module top(Sync,Gate,Done,ena,rst,Tsync,Tgdel,Tgate,Tlen,prev_cnt,prev_cnt_len,prev_state);
	input ena, rst;
	input [7:0]Tsync, Tgdel;
	input [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	input [4:0]prev_state;
	output Sync, Gate, Done;
	wire ena, rst;
	wire [7:0]Tsync, Tgdel;
	wire [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	wire [4:0]prev_state;
	wire Sync, Gate, Done, n_130, n_142, n_164, n_167, n_290, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35;

	nor g63(n_290, Done, n_458);
	not g70(sub_wire0, n_290);
	nor g91(n_130, n_438, prev_cnt_len[5], prev_cnt_len[11], prev_state[1]);
	nor g103(n_142, n_440, prev_cnt_len[15], prev_cnt_len[9], prev_state[3]);
	nor g105(n_167, n_448, prev_cnt[10], prev_cnt[6], prev_cnt[15]);
	nor g111(n_164, n_453, prev_cnt[14], prev_cnt[3], prev_state[3]);
	not g357(n_413, prev_state[1]);
	not g358(n_414, prev_cnt_len[3]);
	not g359(n_415, prev_state[0]);
	not g360(n_416, prev_cnt_len[0]);
	not g361(n_417, prev_cnt_len[7]);
	not g362(n_418, prev_cnt_len[13]);
	not g363(n_419, prev_cnt_len[4]);
	not g364(n_420, prev_cnt_len[10]);
	not g365(n_421, prev_state[2]);
	not g366(n_422, prev_cnt_len[1]);
	not g367(n_423, prev_cnt_len[6]);
	not g368(n_424, prev_cnt_len[12]);
	not g369(n_425, prev_cnt[1]);
	not g370(n_426, prev_state[4]);
	not g371(n_427, rst);
	not g372(n_428, prev_cnt[4]);
	not g373(n_429, prev_cnt[8]);
	not g374(n_430, prev_cnt[12]);
	not g375(n_431, prev_cnt[5]);
	not g376(n_432, prev_cnt[9]);
	not g377(n_433, prev_cnt[13]);
	not g378(n_434, prev_cnt[7]);
	not g379(n_435, prev_cnt[11]);
	not g380(n_436, ena);
	not g381(n_437, prev_cnt[0]);
	nand g382(n_438, n_415, n_414);
	not g383(n_439, n_130);
	nand g384(n_440, n_418, n_417, n_416);
	not g385(n_441, n_142);
	nand g386(n_442, n_421, n_420, n_419);
	nor g387(n_443, n_442, rst, n_426, prev_cnt_len[2]);
	not g388(n_444, n_443);
	nand g389(n_445, n_424, n_423, n_422);
	nor g390(n_446, n_445, n_436, prev_cnt_len[14], prev_cnt_len[8]);
	not g391(n_447, n_446);
	nor g392(Done, n_439, n_441, n_444, n_447);
	nand g393(n_448, n_427, n_426, n_425);
	not g394(n_449, n_167);
	nand g395(n_450, n_430, n_429, n_428);
	nor g396(n_451, n_450, n_436, n_421, prev_cnt[2]);
	not g397(n_452, n_451);
	nand g398(n_453, n_433, n_432, n_431);
	nand g399(n_454, n_413, n_435, n_434);
	not g400(n_455, n_454);
	nand g401(n_456, n_164, n_455, n_415, n_437);
	nor g402(Gate, n_449, n_452, n_456);
	nand g403(n_457, ena, n_427, n_426, n_421);
	nor g404(n_458, n_457, prev_state[3], prev_state[1], n_415);
	and _ECO_0(w_eco0, !prev_state[0], !ena, !prev_cnt_len[14]);
	and _ECO_1(w_eco1, !prev_state[1], !ena, !prev_cnt_len[14]);
	and _ECO_2(w_eco2, !prev_state[0], !prev_cnt_len[6], !prev_cnt_len[12], !prev_cnt_len[14]);
	and _ECO_3(w_eco3, !prev_state[1], prev_cnt_len[8]);
	and _ECO_4(w_eco4, !prev_cnt_len[11], !prev_state[1], prev_state[0], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_5(w_eco5, !prev_state[1], !prev_cnt_len[6], !prev_cnt_len[12], !prev_cnt_len[14]);
	and _ECO_6(w_eco6, !prev_state[0], prev_cnt_len[8]);
	and _ECO_7(w_eco7, prev_state[3], !prev_state[0], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_8(w_eco8, !prev_state[1], prev_state[3], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_9(w_eco9, !prev_state[1], prev_cnt_len[1], !prev_cnt_len[14]);
	and _ECO_10(w_eco10, prev_state[1], !prev_state[0], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_11(w_eco11, !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_12(w_eco12, !prev_cnt_len[11], !prev_state[1], prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_13(w_eco13, prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_14(w_eco14, !prev_state[0], prev_cnt_len[1], !prev_cnt_len[14]);
	and _ECO_15(w_eco15, !prev_state[1], !prev_cnt_len[9], prev_cnt_len[0], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_16(w_eco16, !prev_cnt_len[11], !prev_state[1], prev_state[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_17(w_eco17, prev_state[3], !prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_18(w_eco18, !prev_cnt_len[11], !prev_state[1], prev_cnt_len[3], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_19(w_eco19, !prev_state[1], prev_state[3], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_20(w_eco20, prev_state[3], !prev_state[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_21(w_eco21, prev_state[1], !prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_22(w_eco22, !prev_state[1], prev_state[3], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_23(w_eco23, !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_24(w_eco24, !prev_state[1], !prev_cnt_len[9], !prev_cnt_len[7], !prev_cnt_len[13], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_25(w_eco25, prev_state[1], !prev_state[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_26(w_eco26, prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_27(w_eco27, !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_28(w_eco28, !prev_state[1], !prev_cnt_len[9], prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_29(w_eco29, prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_30(w_eco30, !prev_cnt_len[11], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_31(w_eco31, !prev_state[1], !prev_cnt_len[9], prev_cnt_len[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_32(w_eco32, !prev_cnt_len[11], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_33(w_eco33, !prev_state[1], !prev_cnt_len[9], !prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_34(w_eco34, !prev_state[1], !prev_cnt_len[9], !prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	or _ECO_35(w_eco35, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34);
	xor _ECO_out0(Sync, sub_wire0, w_eco35);

endmodule