module top(Sync,Gate,Done,clk,ena,rst,Tsync,Tgdel,Tgate,Tlen,prev_cnt,prev_cnt_len,prev_state);
	input clk, ena, rst;
	input [7:0]Tsync, Tgdel;
	input [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	input [4:0]prev_state;
	output Sync, Gate, Done;
	wire clk, ena, rst;
	wire [7:0]Tsync, Tgdel;
	wire [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	wire [4:0]prev_state;
	wire Sync, Gate, Done, n_130, n_142, n_164, n_167, n_290, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, sub_wire1, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, sub_wire2, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182;

	nor g63(n_290, Done, n_458);
	not g70(sub_wire1, n_290);
	nor g91(n_130, n_438, prev_cnt_len[5], prev_cnt_len[11], prev_state[1]);
	nor g103(n_142, n_440, prev_cnt_len[15], prev_cnt_len[9], prev_state[3]);
	nor g105(n_167, n_448, prev_cnt[10], prev_cnt[6], prev_cnt[15]);
	nor g111(n_164, n_453, prev_cnt[14], prev_cnt[3], prev_state[3]);
	not g357(n_413, prev_state[1]);
	not g358(n_414, prev_cnt_len[3]);
	not g359(n_415, prev_state[0]);
	not g360(n_416, prev_cnt_len[0]);
	not g361(n_417, prev_cnt_len[7]);
	not g362(n_418, prev_cnt_len[13]);
	not g363(n_419, prev_cnt_len[4]);
	not g364(n_420, prev_cnt_len[10]);
	not g365(n_421, prev_state[2]);
	not g366(n_422, prev_cnt_len[1]);
	not g367(n_423, prev_cnt_len[6]);
	not g368(n_424, prev_cnt_len[12]);
	not g369(n_425, prev_cnt[1]);
	not g370(n_426, prev_state[4]);
	not g371(n_427, rst);
	not g372(n_428, prev_cnt[4]);
	not g373(n_429, prev_cnt[8]);
	not g374(n_430, prev_cnt[12]);
	not g375(n_431, prev_cnt[5]);
	not g376(n_432, prev_cnt[9]);
	not g377(n_433, prev_cnt[13]);
	not g378(n_434, prev_cnt[7]);
	not g379(n_435, prev_cnt[11]);
	not g380(n_436, ena);
	not g381(n_437, prev_cnt[0]);
	nand g382(n_438, n_415, n_414);
	not g383(n_439, n_130);
	nand g384(n_440, n_418, n_417, n_416);
	not g385(n_441, n_142);
	nand g386(n_442, n_421, n_420, n_419);
	nor g387(n_443, n_442, rst, n_426, prev_cnt_len[2]);
	not g388(n_444, n_443);
	nand g389(n_445, n_424, n_423, n_422);
	nor g390(n_446, n_445, n_436, prev_cnt_len[14], prev_cnt_len[8]);
	not g391(n_447, n_446);
	nor g392(sub_wire0, n_439, n_441, n_444, n_447);
	nand g393(n_448, n_427, n_426, n_425);
	not g394(n_449, n_167);
	nand g395(n_450, n_430, n_429, n_428);
	nor g396(n_451, n_450, n_436, n_421, prev_cnt[2]);
	not g397(n_452, n_451);
	nand g398(n_453, n_433, n_432, n_431);
	nand g399(n_454, n_413, n_435, n_434);
	not g400(n_455, n_454);
	nand g401(n_456, n_164, n_455, n_415, n_437);
	nor g402(sub_wire2, n_449, n_452, n_456);
	nand g403(n_457, ena, n_427, n_426, n_421);
	nor g404(n_458, n_457, prev_state[3], prev_state[1], n_415);
	and _ECO_0(w_eco0, prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1(w_eco1, prev_state[4], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_2(w_eco2, !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_3(w_eco3, prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_4(w_eco4, !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_5(w_eco5, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_6(w_eco6, !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_7(w_eco7, !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_8(w_eco8, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_9(w_eco9, !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_10(w_eco10, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_11(w_eco11, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_12(w_eco12, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_13(w_eco13, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_14(w_eco14, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_15(w_eco15, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_16(w_eco16, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_17(w_eco17, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_18(w_eco18, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_19(w_eco19, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_20(w_eco20, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_21(w_eco21, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_22(w_eco22, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_23(w_eco23, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_24(w_eco24, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_25(w_eco25, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_26(w_eco26, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_27(w_eco27, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_28(w_eco28, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_29(w_eco29, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	or _ECO_30(w_eco30, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29);
	xor _ECO_out0(Done, sub_wire0, w_eco30);
	and _ECO_31(w_eco31, prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_32(w_eco32, prev_state[1], prev_state[0]);
	and _ECO_33(w_eco33, !prev_state[3], prev_state[0], !prev_state[2], prev_state[4]);
	and _ECO_34(w_eco34, !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_35(w_eco35, !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_36(w_eco36, !prev_state[3], prev_state[0], !prev_state[2], !rst, ena);
	and _ECO_37(w_eco37, prev_state[4], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_38(w_eco38, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_39(w_eco39, prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_40(w_eco40, !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_41(w_eco41, !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_42(w_eco42, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_43(w_eco43, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_44(w_eco44, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_45(w_eco45, !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_46(w_eco46, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_47(w_eco47, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_48(w_eco48, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_49(w_eco49, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_50(w_eco50, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_51(w_eco51, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_52(w_eco52, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_53(w_eco53, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_54(w_eco54, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_55(w_eco55, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_56(w_eco56, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_57(w_eco57, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_58(w_eco58, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_59(w_eco59, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_60(w_eco60, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_61(w_eco61, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_62(w_eco62, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_63(w_eco63, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	or _ECO_64(w_eco64, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63);
	xor _ECO_out1(Sync, sub_wire1, w_eco64);
	and _ECO_65(w_eco65, !prev_state[3], prev_state[4], prev_cnt[0]);
	and _ECO_66(w_eco66, prev_state[3], prev_state[0], !prev_cnt[0], prev_cnt[2]);
	and _ECO_67(w_eco67, !prev_state[3], !prev_state[0], prev_state[4], prev_cnt[7]);
	and _ECO_68(w_eco68, prev_state[1], !prev_state[3], prev_state[0], ena, prev_cnt[0]);
	and _ECO_69(w_eco69, prev_state[0], !prev_state[4], !ena, !prev_cnt[0], prev_cnt[2]);
	and _ECO_70(w_eco70, prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt[0]);
	and _ECO_71(w_eco71, prev_cnt[15], prev_state[0], !prev_state[4], !ena, !prev_cnt[0]);
	and _ECO_72(w_eco72, !prev_state[3], prev_state[0], !prev_state[2], !rst, ena, prev_cnt[0]);
	and _ECO_73(w_eco73, !prev_state[1], prev_state[0], !prev_state[4], rst, !prev_cnt[0], prev_cnt[2]);
	and _ECO_74(w_eco74, prev_state[3], prev_state[0], prev_state[2], !ena, !prev_cnt[0]);
	and _ECO_75(w_eco75, !prev_state[1], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[0], prev_cnt[2]);
	and _ECO_76(w_eco76, !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_state[2], prev_state[4], !prev_cnt[2]);
	and _ECO_77(w_eco77, prev_state[0], prev_state[2], !prev_state[4], !ena, !prev_cnt[0]);
	and _ECO_78(w_eco78, prev_state[3], !prev_cnt[6], prev_state[0], prev_cnt[1], !prev_cnt[0]);
	and _ECO_79(w_eco79, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_80(w_eco80, !prev_state[1], prev_cnt[15], prev_state[0], !prev_state[4], rst, !prev_cnt[0]);
	and _ECO_81(w_eco81, prev_state[3], prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[0]);
	and _ECO_82(w_eco82, !prev_cnt[6], prev_state[0], prev_cnt[1], !prev_state[4], !ena, !prev_cnt[0]);
	and _ECO_83(w_eco83, prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt[0]);
	and _ECO_84(w_eco84, !prev_state[1], !prev_state[3], !prev_state[0], prev_state[4], !prev_cnt[11]);
	and _ECO_85(w_eco85, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_86(w_eco86, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[4], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_87(w_eco87, !prev_state[1], prev_cnt[15], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[0]);
	and _ECO_88(w_eco88, !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[4], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_89(w_eco89, prev_state[1], !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_90(w_eco90, prev_state[3], prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[0]);
	and _ECO_91(w_eco91, prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_state[4], !ena, !prev_cnt[0]);
	and _ECO_92(w_eco92, !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_state[2], !prev_cnt[1], prev_state[4], !prev_cnt[2]);
	and _ECO_93(w_eco93, !prev_cnt[6], prev_state[0], !prev_state[4], !rst, !ena, !prev_cnt[0]);
	and _ECO_94(w_eco94, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_95(w_eco95, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[4], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_96(w_eco96, !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_state[0], prev_state[4]);
	and _ECO_97(w_eco97, prev_state[1], !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], ena, !prev_cnt[2]);
	and _ECO_98(w_eco98, !prev_state[1], !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[4], !rst, prev_cnt[4], ena, !prev_cnt[0], !prev_cnt[2]);
	and _ECO_99(w_eco99, !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[4], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_100(w_eco100, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_101(w_eco101, !prev_state[3], prev_cnt[3], prev_state[2], !prev_state[4], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_102(w_eco102, !prev_state[3], !prev_cnt[3], !prev_state[0], prev_state[4], prev_cnt[5]);
	and _ECO_103(w_eco103, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_104(w_eco104, !prev_state[1], prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[0]);
	and _ECO_105(w_eco105, !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !rst, ena, !prev_cnt[2]);
	and _ECO_106(w_eco106, !prev_state[1], !prev_cnt[6], prev_state[0], prev_cnt[1], !prev_state[4], rst, !prev_cnt[0]);
	and _ECO_107(w_eco107, prev_state[3], !prev_cnt[6], prev_state[0], !prev_state[4], !rst, !prev_cnt[0]);
	and _ECO_108(w_eco108, !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_109(w_eco109, prev_state[1], !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_110(w_eco110, !prev_state[1], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[0]);
	and _ECO_111(w_eco111, prev_state[1], !prev_state[3], prev_cnt[3], prev_state[2], !prev_state[4], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_112(w_eco112, !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_113(w_eco113, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_114(w_eco114, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_115(w_eco115, !prev_state[3], !prev_cnt[3], !prev_state[0], prev_state[4], !prev_cnt[9], !prev_cnt[13]);
	and _ECO_116(w_eco116, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_117(w_eco117, !prev_state[1], !prev_cnt[6], prev_state[0], prev_state[2], !prev_state[4], !rst, !prev_cnt[0]);
	and _ECO_118(w_eco118, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_state[4], rst, !prev_cnt[0]);
	and _ECO_119(w_eco119, prev_state[1], !prev_state[3], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_120(w_eco120, !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_121(w_eco121, !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_122(w_eco122, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_123(w_eco123, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt[1], !prev_state[4], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_124(w_eco124, !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[4], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_125(w_eco125, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_126(w_eco126, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_127(w_eco127, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_128(w_eco128, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_129(w_eco129, prev_state[1], !prev_state[3], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], rst, ena, !prev_cnt[2]);
	and _ECO_130(w_eco130, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_131(w_eco131, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_132(w_eco132, !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_133(w_eco133, !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_134(w_eco134, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[4], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_135(w_eco135, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_136(w_eco136, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_137(w_eco137, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_138(w_eco138, !prev_state[3], !prev_cnt[14], prev_state[2], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_139(w_eco139, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_140(w_eco140, prev_state[1], !prev_state[3], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_141(w_eco141, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_142(w_eco142, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_143(w_eco143, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_144(w_eco144, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[4], !rst, !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_145(w_eco145, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_146(w_eco146, prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_147(w_eco147, !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_148(w_eco148, !prev_state[3], !prev_cnt[14], prev_state[2], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_149(w_eco149, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_150(w_eco150, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_151(w_eco151, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_152(w_eco152, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_153(w_eco153, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_154(w_eco154, prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_155(w_eco155, !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_156(w_eco156, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_157(w_eco157, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_158(w_eco158, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_159(w_eco159, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_160(w_eco160, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_161(w_eco161, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_162(w_eco162, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_163(w_eco163, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_164(w_eco164, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_165(w_eco165, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_166(w_eco166, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_167(w_eco167, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_168(w_eco168, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_169(w_eco169, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_170(w_eco170, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_171(w_eco171, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_172(w_eco172, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_173(w_eco173, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_174(w_eco174, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_175(w_eco175, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_176(w_eco176, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_177(w_eco177, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_178(w_eco178, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_179(w_eco179, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_state[4], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_180(w_eco180, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_181(w_eco181, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	or _ECO_182(w_eco182, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181);
	xor _ECO_out2(Gate, sub_wire2, w_eco182);

endmodule