module top(next_state,cur_state,at_sendreg,at_senddmaa,at_sendpios,at_senddmas,at_sendbista,at_senddata,lk_txfsmidle,lk_txerror,r2t_waittxid,r2t_rxempty,txtimeout,expire,tptx_reset);
	input [14:0]cur_state;
	input at_sendreg, at_senddmaa, at_sendpios, at_senddmas, at_sendbista, at_senddata, lk_txfsmidle, lk_txerror, r2t_waittxid, r2t_rxempty, txtimeout, expire, tptx_reset;
	output [14:0]next_state;
	wire [14:0]cur_state;
	wire at_sendreg, at_senddmaa, at_sendpios, at_senddmas, at_sendbista, at_senddata, lk_txfsmidle, lk_txerror, r2t_waittxid, r2t_rxempty, txtimeout, expire, tptx_reset;
	wire [14:0]next_state;
	wire n_27, n_62, n_63, n_64, n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_159, n_161, n_162, n_183, n_184, n_185, n_190, n_301, n_302, n_303, n_304, n_305, n_508, n_522, n_530, n_547, n_558, n_566, n_575, n_583, n_594, n_602, n_618, n_625, n_1112, n_1114, n_1115, n_1603, n_1604, n_1628, n_1629, n_1630, n_1631, n_1632, n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640, n_1641, n_1642, n_1643, n_1644, n_1645, n_1646, n_1647, n_1648, n_1649, n_1650, n_1651, n_1652, n_1653, n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661, n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669, n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677, n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685, n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693, n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701, n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1709, n_1710, n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718, n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726, n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734, n_1735, n_1736, n_1737, n_1738, n_1739, n_1740, n_1741, n_1742, n_1743, n_1744, n_1745, n_1746, n_1747, n_1748, n_1749, n_1750, n_1751, n_1752, n_1753, n_1754, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760, n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768, n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776, n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784, n_1785, n_1786, n_1787, n_1788, n_1789, n_1790;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, sub_wire1, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, sub_wire2, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, sub_wire3, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, sub_wire4, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, sub_wire5, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, sub_wire6, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472;

	nor g112(n_76, n_1655, n_184, n_185, n_190);
	nor g110(n_75, n_1657, n_184, n_185, n_190);
	nor g102(n_71, n_183, n_1659, n_185, n_190);
	nor g104(n_72, n_183, n_1661, n_185, n_190);
	nor g106(n_73, n_1663, n_184, n_185, n_190);
	nor g108(n_74, n_1665, n_184, n_185, n_190);
	nor g92(n_66, n_183, n_184, n_1667, n_190);
	nor g94(n_67, n_183, n_184, n_1669, n_190);
	nor g96(n_68, n_183, n_184, n_1671, n_190);
	nor g98(n_69, n_183, n_1673, n_185, n_190);
	nor g83(n_62, n_183, n_184, n_185, n_1675);
	nor g85(n_63, n_183, n_184, n_185, n_1677);
	nor g87(n_64, n_183, n_184, n_185, n_1679);
	nor g90(n_65, n_183, n_184, n_1681, n_190);
	nor g100(n_70, n_183, n_1683, n_185, n_190);
	nand g117(n_305, n_301, n_302, n_303, n_304);
	nor g116(n_304, n_74, n_75, n_76);
	nor g115(n_303, n_70, n_71, n_72, n_73);
	nor g114(n_302, n_66, n_67, n_68, n_69);
	nor g113(n_301, n_62, n_63, n_64, n_65);
	nor g76(n_1112, at_senddmas, at_senddmaa, at_sendbista, at_senddata);
	nor g719(n_27, lk_txfsmidle, txtimeout);
	nand g739(n_159, lk_txfsmidle, r2t_rxempty);
	nor g772(n_625, n_305, tptx_reset);
	nor g801(n_1115, n_27, lk_txfsmidle);
	nor g802(n_1114, n_27, lk_txerror);
	not g1440(n_1628, at_senddata);
	not g1441(n_1629, at_sendbista);
	not g1442(n_1630, at_senddmaa);
	not g1443(n_1631, at_senddmas);
	not g1444(n_1632, lk_txfsmidle);
	not g1445(n_1633, r2t_rxempty);
	not g1446(n_1634, tptx_reset);
	not g1447(n_1635, lk_txerror);
	not g1448(n_1636, expire);
	not g1449(n_1637, cur_state[11]);
	not g1450(n_1638, cur_state[12]);
	not g1451(n_1639, cur_state[13]);
	not g1452(n_1640, cur_state[14]);
	not g1453(n_1641, cur_state[7]);
	not g1454(n_1642, cur_state[8]);
	not g1455(n_1643, cur_state[9]);
	not g1456(n_1644, cur_state[10]);
	not g1457(n_1645, cur_state[3]);
	not g1458(n_1646, cur_state[4]);
	not g1459(n_1647, cur_state[5]);
	not g1460(n_1648, cur_state[6]);
	not g1461(n_1649, cur_state[0]);
	not g1462(n_1650, cur_state[1]);
	not g1463(n_1651, cur_state[2]);
	not g1464(n_1652, at_sendpios);
	not g1465(n_1653, at_sendreg);
	not g1466(n_1654, r2t_waittxid);
	nand g1467(n_1655, cur_state[14], n_1639, n_1638, n_1637);
	nand g1468(n_184, n_1644, n_1643, n_1642, n_1641);
	nand g1469(n_185, n_1648, n_1647, n_1646, n_1645);
	nand g1470(n_190, n_1651, n_1650, n_1649);
	not g1471(n_1656, n_76);
	nand g1472(n_1657, n_1640, cur_state[13], n_1638, n_1637);
	not g1473(n_1658, n_75);
	nand g1474(n_183, n_1640, n_1639, n_1638, n_1637);
	nand g1475(n_1659, n_1644, cur_state[9], n_1642, n_1641);
	not g1476(n_1660, n_71);
	nand g1477(n_1661, cur_state[10], n_1643, n_1642, n_1641);
	not g1478(n_1662, n_72);
	nand g1479(n_1663, n_1640, n_1639, n_1638, cur_state[11]);
	not g1480(n_1664, n_73);
	nand g1481(n_1665, n_1640, n_1639, cur_state[12], n_1637);
	not g1482(n_1666, n_74);
	nand g1483(n_1667, n_1648, n_1647, cur_state[4], n_1645);
	not g1484(n_1668, n_66);
	nand g1485(n_1669, n_1648, cur_state[5], n_1646, n_1645);
	not g1486(n_1670, n_67);
	nand g1487(n_1671, cur_state[6], n_1647, n_1646, n_1645);
	not g1488(n_1672, n_68);
	nand g1489(n_1673, n_1644, n_1643, n_1642, cur_state[7]);
	not g1490(n_1674, n_69);
	nand g1491(n_1675, n_1651, n_1650, cur_state[0]);
	not g1492(n_1676, n_62);
	nand g1493(n_1677, n_1651, cur_state[1], n_1649);
	not g1494(n_1678, n_63);
	nand g1495(n_1679, cur_state[2], n_1650, n_1649);
	not g1496(n_1680, n_64);
	nand g1497(n_1681, n_1648, n_1647, n_1646, cur_state[3]);
	not g1498(n_1682, n_65);
	nand g1499(n_1683, n_1644, n_1643, cur_state[8], n_1641);
	not g1500(n_1684, n_70);
	nor g1501(n_1603, n_1676, tptx_reset);
	not g1502(n_1685, n_1603);
	not g1503(n_1686, n_159);
	nand g1504(n_161, n_1686, n_1653, n_1652);
	not g1505(n_1687, n_161);
	nand g1506(n_162, n_1687, n_1630, n_1631);
	nor g1507(n_1688, n_162, at_sendbista, n_1628);
	not g1508(n_1689, n_1688);
	nor g1509(next_state[7], n_1685, n_1689);
	not g1510(n_1690, n_1112);
	not g1511(n_1691, n_27);
	not g1512(n_1692, n_625);
	not g1513(n_1693, n_1115);
	not g1514(n_1694, n_1114);
	nor g1515(n_1695, n_1685, r2t_rxempty);
	not g1516(n_1696, n_1695);
	nor g1517(n_1604, n_1678, tptx_reset);
	not g1518(n_1697, n_1604);
	nor g1519(n_1698, n_1697, r2t_waittxid);
	not g1520(n_1699, n_1698);
	nand g1521(next_state[1], n_1696, n_1699);
	nor g1522(n_530, n_1656, tptx_reset);
	not g1523(n_1700, n_530);
	nor g1524(n_547, n_1658, tptx_reset);
	not g1525(n_1701, n_547);
	nor g1526(n_566, n_1666, tptx_reset);
	not g1527(n_1702, n_566);
	nor g1528(n_583, n_1664, tptx_reset);
	not g1529(n_1703, n_583);
	nor g1530(n_602, n_1662, tptx_reset);
	not g1531(n_1704, n_602);
	nand g1532(n_1705, n_1701, n_1702, n_1703, n_1704);
	not g1533(n_1706, n_1705);
	nand g1534(n_1707, n_1700, n_1706);
	not g1535(n_1708, n_1707);
	nand g1536(n_1709, n_1693, n_1694);
	not g1537(n_1710, n_1709);
	nor g1538(n_1711, n_1708, n_1710);
	not g1539(n_1712, n_1711);
	nor g1540(n_522, n_1672, tptx_reset);
	not g1541(n_1713, n_522);
	nor g1542(n_1714, n_1713, n_1636);
	not g1543(n_1715, n_1714);
	nor g1544(n_1716, n_1700, n_1691);
	not g1545(n_1717, n_1716);
	nor g1546(n_1718, n_1701, n_1691);
	not g1547(n_1719, n_1718);
	nor g1548(n_558, n_1668, tptx_reset);
	not g1549(n_1720, n_558);
	nor g1550(n_1721, n_1720, n_1636);
	not g1551(n_1722, n_1721);
	nor g1552(n_1723, n_1702, n_1691);
	not g1553(n_1724, n_1723);
	nor g1554(n_575, n_1682, tptx_reset);
	not g1555(n_1725, n_575);
	nor g1556(n_1726, n_1725, n_1636);
	not g1557(n_1727, n_1726);
	nor g1558(n_1728, n_1703, n_1691);
	not g1559(n_1729, n_1728);
	nor g1560(n_594, n_1680, tptx_reset);
	not g1561(n_1730, n_594);
	nor g1562(n_1731, n_1730, n_1636);
	not g1563(n_1732, n_1731);
	nor g1564(n_1733, n_1704, n_1691);
	not g1565(n_1734, n_1733);
	nor g1566(n_618, n_1684, tptx_reset);
	not g1567(n_1735, n_618);
	nor g1568(n_1736, n_1735, n_1636);
	not g1569(n_1737, n_1736);
	nor g1570(n_508, n_27, n_1632, n_1635);
	not g1571(n_1738, n_508);
	nor g1572(n_1739, n_1701, n_1738);
	not g1573(n_1740, n_1739);
	nor g1574(n_1741, n_1702, n_1738);
	not g1575(n_1742, n_1741);
	nor g1576(n_1743, n_1703, n_1738);
	not g1577(n_1744, n_1743);
	nor g1578(n_1745, n_1704, n_1738);
	not g1579(n_1746, n_1745);
	nor g1580(n_1747, n_1700, n_1738);
	not g1581(n_1748, n_1747);
	nand g1582(next_state[14], n_1715, n_1717);
	nor g1583(n_1749, n_1670, tptx_reset);
	not g1584(n_1750, n_1749);
	nand g1585(next_state[13], n_1750, n_1719);
	nand g1586(next_state[12], n_1722, n_1724);
	nand g1587(next_state[11], n_1727, n_1729);
	nand g1588(next_state[10], n_1732, n_1734);
	nor g1589(n_1751, n_1674, tptx_reset);
	not g1590(n_1752, n_1751);
	nor g1591(n_1753, n_1735, expire);
	not g1592(n_1754, n_1753);
	nand g1593(next_state[8], n_1752, n_1754);
	nand g1594(sub_wire0, n_1737, n_1692);
	nor g1595(n_1755, n_161, n_1630, at_senddmas);
	not g1596(n_1756, n_1755);
	nor g1597(n_1757, n_1756, n_1685);
	not g1598(n_1758, n_1757);
	nand g1599(sub_wire1, n_1758, n_1740);
	nor g1600(n_1759, n_161, n_1685, n_1631);
	not g1601(n_1760, n_1759);
	nor g1602(n_1761, n_1720, expire);
	not g1603(n_1762, n_1761);
	nand g1604(sub_wire2, n_1760, n_1762, n_1742);
	nor g1605(n_1763, n_159, at_sendreg, n_1652);
	not g1606(n_1764, n_1763);
	nor g1607(n_1765, n_1764, n_1685);
	not g1608(n_1766, n_1765);
	nor g1609(n_1767, n_1725, expire);
	not g1610(n_1768, n_1767);
	nand g1611(sub_wire3, n_1766, n_1768, n_1744);
	nor g1612(n_1769, n_159, n_1685, n_1653);
	not g1613(n_1770, n_1769);
	nor g1614(n_1771, n_1730, expire);
	not g1615(n_1772, n_1771);
	nand g1616(sub_wire4, n_1770, n_1772, n_1746);
	nor g1617(n_1773, n_1685, n_162, n_1629);
	not g1618(n_1774, n_1773);
	nor g1619(n_1775, n_1713, expire);
	not g1620(n_1776, n_1775);
	nand g1621(sub_wire5, n_1774, n_1776, n_1748);
	nor g1622(n_1777, n_1660, tptx_reset);
	not g1623(n_1778, n_1777);
	nor g1624(n_1779, n_1685, lk_txfsmidle, n_1633);
	not g1625(n_1780, n_1779);
	nor g1626(n_1781, at_sendreg, at_sendpios, n_1632, n_1633);
	not g1627(n_1782, n_1781);
	nor g1628(n_1783, n_1690, n_1782, n_1685);
	not g1629(n_1784, n_1783);
	nor g1630(n_1785, n_1697, n_1654);
	not g1631(n_1786, n_1785);
	nand g1632(n_1787, n_1778, n_1780, n_1784, n_1786);
	not g1633(n_1788, n_1787);
	nand g1634(n_1789, n_1788, n_1634);
	not g1635(n_1790, n_1789);
	nand g1636(sub_wire6, n_1790, n_1712);
	and _ECO_0(w_eco0, !tptx_reset, !lk_txerror, expire, cur_state[3], !cur_state[0], cur_state[1]);
	and _ECO_1(w_eco1, !at_senddmas, !at_senddmaa, !tptx_reset, cur_state[3], cur_state[0], cur_state[1]);
	and _ECO_2(w_eco2, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[3], !cur_state[0], cur_state[1]);
	and _ECO_3(w_eco3, lk_txfsmidle, !tptx_reset, expire, cur_state[3], !cur_state[0], cur_state[1]);
	and _ECO_4(w_eco4, !tptx_reset, !lk_txerror, expire, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_5(w_eco5, !tptx_reset, !lk_txerror, expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_6(w_eco6, !at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_7(w_eco7, !at_senddmas, !at_senddmaa, !tptx_reset, cur_state[3], cur_state[0], cur_state[2]);
	and _ECO_8(w_eco8, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_9(w_eco9, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1]);
	and _ECO_10(w_eco10, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_11(w_eco11, lk_txfsmidle, !tptx_reset, expire, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_12(w_eco12, lk_txfsmidle, !tptx_reset, expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_13(w_eco13, !tptx_reset, !lk_txerror, expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_14(w_eco14, !tptx_reset, !lk_txerror, expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_15(w_eco15, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_16(w_eco16, !at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_17(w_eco17, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_18(w_eco18, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2]);
	and _ECO_19(w_eco19, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1]);
	and _ECO_20(w_eco20, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_21(w_eco21, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_22(w_eco22, lk_txfsmidle, !tptx_reset, expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_23(w_eco23, lk_txfsmidle, !tptx_reset, expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_24(w_eco24, !tptx_reset, !lk_txerror, expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_25(w_eco25, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_26(w_eco26, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_27(w_eco27, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_28(w_eco28, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_29(w_eco29, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_30(w_eco30, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_31(w_eco31, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2]);
	and _ECO_32(w_eco32, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_33(w_eco33, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_34(w_eco34, lk_txfsmidle, !tptx_reset, expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_35(w_eco35, !tptx_reset, !lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_36(w_eco36, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_37(w_eco37, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_38(w_eco38, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_39(w_eco39, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_40(w_eco40, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_41(w_eco41, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_42(w_eco42, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_43(w_eco43, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_44(w_eco44, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_45(w_eco45, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_46(w_eco46, lk_txfsmidle, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_47(w_eco47, !tptx_reset, !lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_48(w_eco48, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_49(w_eco49, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_50(w_eco50, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_51(w_eco51, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_52(w_eco52, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_53(w_eco53, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_54(w_eco54, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_55(w_eco55, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_56(w_eco56, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_57(w_eco57, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_58(w_eco58, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_59(w_eco59, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_60(w_eco60, lk_txfsmidle, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_61(w_eco61, !tptx_reset, !lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_62(w_eco62, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_63(w_eco63, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_64(w_eco64, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_65(w_eco65, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_66(w_eco66, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_67(w_eco67, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_68(w_eco68, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_69(w_eco69, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_70(w_eco70, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_71(w_eco71, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_72(w_eco72, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_73(w_eco73, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_74(w_eco74, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_75(w_eco75, !tptx_reset, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_76(w_eco76, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_77(w_eco77, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_78(w_eco78, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_79(w_eco79, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_80(w_eco80, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_81(w_eco81, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_82(w_eco82, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_83(w_eco83, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_84(w_eco84, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_85(w_eco85, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_86(w_eco86, !tptx_reset, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_87(w_eco87, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_88(w_eco88, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_89(w_eco89, !at_senddmas, !at_senddmaa, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_90(w_eco90, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_91(w_eco91, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_92(w_eco92, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_93(w_eco93, !tptx_reset, expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_94(w_eco94, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_95(w_eco95, !tptx_reset, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_96(w_eco96, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_97(w_eco97, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_98(w_eco98, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_99(w_eco99, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_100(w_eco100, !tptx_reset, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_101(w_eco101, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_102(w_eco102, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_103(w_eco103, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_104(w_eco104, !at_senddmas, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendreg);
	or _ECO_105(w_eco105, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104);
	xor _ECO_out0(next_state[9], sub_wire0, w_eco105);
	and _ECO_106(w_eco106, !at_senddmas, !lk_txerror, expire, !cur_state[0]);
	and _ECO_107(w_eco107, !at_senddmas, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_108(w_eco108, !at_senddmas, tptx_reset);
	and _ECO_109(w_eco109, !at_senddmas, cur_state[11], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_110(w_eco110, !at_senddmas, lk_txfsmidle, expire, !cur_state[0]);
	and _ECO_111(w_eco111, at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_112(w_eco112, !at_senddmas, at_senddmaa, cur_state[0], !at_sendpios, at_sendreg);
	and _ECO_113(w_eco113, !at_senddmas, !cur_state[1], !cur_state[2]);
	and _ECO_114(w_eco114, at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_115(w_eco115, at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_116(w_eco116, !at_senddmas, expire, cur_state[11], !cur_state[3], cur_state[4]);
	and _ECO_117(w_eco117, at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_118(w_eco118, !at_senddmas, !lk_txerror, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_119(w_eco119, !at_senddmas, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_120(w_eco120, at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_121(w_eco121, at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_122(w_eco122, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_123(w_eco123, !at_senddmas, cur_state[7], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_124(w_eco124, at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_125(w_eco125, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_126(w_eco126, at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_127(w_eco127, !at_senddmas, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_128(w_eco128, !at_senddmas, lk_txfsmidle, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_129(w_eco129, !at_senddmas, !lk_txerror, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_130(w_eco130, at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_131(w_eco131, at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_132(w_eco132, at_senddmaa, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_133(w_eco133, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_134(w_eco134, !at_senddmas, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_135(w_eco135, !at_senddmas, expire, cur_state[7], !cur_state[3], cur_state[4]);
	and _ECO_136(w_eco136, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_137(w_eco137, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_138(w_eco138, at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_139(w_eco139, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_140(w_eco140, !at_senddmas, at_senddmaa, !r2t_rxempty, cur_state[0], !at_sendpios);
	and _ECO_141(w_eco141, !at_senddmas, !lk_txerror, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_142(w_eco142, !at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_143(w_eco143, !at_senddmas, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_144(w_eco144, at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_145(w_eco145, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_146(w_eco146, at_senddmaa, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_147(w_eco147, !at_senddmas, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_148(w_eco148, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_149(w_eco149, !at_senddmas, !lk_txfsmidle, lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4]);
	and _ECO_150(w_eco150, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_151(w_eco151, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_152(w_eco152, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_153(w_eco153, !at_senddmas, at_senddmaa, !lk_txfsmidle, cur_state[0], !at_sendpios);
	and _ECO_154(w_eco154, !at_senddmas, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_155(w_eco155, !at_senddmas, expire, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_156(w_eco156, !at_senddmas, lk_txfsmidle, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_157(w_eco157, !at_senddmas, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_158(w_eco158, at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_159(w_eco159, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_160(w_eco160, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_161(w_eco161, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_162(w_eco162, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_163(w_eco163, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_164(w_eco164, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_165(w_eco165, !at_senddmas, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_166(w_eco166, !at_senddmas, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_167(w_eco167, !at_senddmas, expire, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_168(w_eco168, at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_169(w_eco169, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_170(w_eco170, !at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_171(w_eco171, !at_senddmas, !lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_172(w_eco172, !at_senddmas, !lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_173(w_eco173, at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_174(w_eco174, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_175(w_eco175, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_176(w_eco176, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_177(w_eco177, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_178(w_eco178, !at_senddmas, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_179(w_eco179, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_180(w_eco180, at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_181(w_eco181, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_182(w_eco182, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_183(w_eco183, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_184(w_eco184, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_185(w_eco185, !at_senddmas, !lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_186(w_eco186, !at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_187(w_eco187, !at_senddmas, !lk_txfsmidle, lk_txerror, !expire, cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_188(w_eco188, !at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0]);
	and _ECO_189(w_eco189, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_190(w_eco190, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_191(w_eco191, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_192(w_eco192, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_193(w_eco193, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_194(w_eco194, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_195(w_eco195, at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_196(w_eco196, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_197(w_eco197, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_198(w_eco198, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_199(w_eco199, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_200(w_eco200, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_201(w_eco201, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_202(w_eco202, !at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_203(w_eco203, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_204(w_eco204, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_205(w_eco205, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_206(w_eco206, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_207(w_eco207, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_208(w_eco208, at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_209(w_eco209, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_210(w_eco210, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_211(w_eco211, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_212(w_eco212, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_213(w_eco213, !at_senddmas, !lk_txfsmidle, lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_214(w_eco214, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_215(w_eco215, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_216(w_eco216, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_217(w_eco217, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_218(w_eco218, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios);
	and _ECO_219(w_eco219, at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_220(w_eco220, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_221(w_eco221, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_222(w_eco222, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_223(w_eco223, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_224(w_eco224, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_225(w_eco225, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_226(w_eco226, at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios);
	and _ECO_227(w_eco227, at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	or _ECO_228(w_eco228, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227);
	xor _ECO_out1(next_state[5], sub_wire1, w_eco228);
	and _ECO_229(w_eco229, at_senddmas, !lk_txerror, expire, !cur_state[0]);
	and _ECO_230(w_eco230, at_senddmas, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_231(w_eco231, at_senddmas, tptx_reset);
	and _ECO_232(w_eco232, at_senddmas, cur_state[11], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_233(w_eco233, at_senddmas, lk_txfsmidle, expire, !cur_state[0]);
	and _ECO_234(w_eco234, at_senddmas, !lk_txerror, cur_state[11], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_235(w_eco235, at_senddmas, !cur_state[1], !cur_state[2]);
	and _ECO_236(w_eco236, !at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_237(w_eco237, at_senddmas, lk_txfsmidle, r2t_rxempty, cur_state[0], !at_sendreg);
	and _ECO_238(w_eco238, !at_senddmas, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_239(w_eco239, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_240(w_eco240, at_senddmas, expire, cur_state[11], !cur_state[3], cur_state[4]);
	and _ECO_241(w_eco241, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_242(w_eco242, at_senddmas, lk_txfsmidle, cur_state[11], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_243(w_eco243, !tptx_reset, !lk_txerror, !expire, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_244(w_eco244, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_245(w_eco245, at_senddmas, !lk_txerror, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_246(w_eco246, !at_senddmas, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_247(w_eco247, at_senddmas, cur_state[7], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_248(w_eco248, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_249(w_eco249, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_250(w_eco250, at_senddmas, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_251(w_eco251, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_252(w_eco252, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_253(w_eco253, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_254(w_eco254, at_senddmas, expire, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_255(w_eco255, at_senddmas, !lk_txerror, cur_state[7], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_256(w_eco256, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_257(w_eco257, !tptx_reset, !lk_txerror, !expire, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_258(w_eco258, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_259(w_eco259, at_senddmas, !lk_txerror, cur_state[11], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_260(w_eco260, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_261(w_eco261, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_262(w_eco262, at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_263(w_eco263, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_264(w_eco264, !at_senddmas, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_265(w_eco265, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_266(w_eco266, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_267(w_eco267, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_268(w_eco268, at_senddmas, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_269(w_eco269, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_270(w_eco270, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_271(w_eco271, at_senddmas, expire, cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_272(w_eco272, at_senddmas, expire, cur_state[7], !cur_state[3], cur_state[4]);
	and _ECO_273(w_eco273, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_274(w_eco274, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_275(w_eco275, !at_senddmas, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_276(w_eco276, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_277(w_eco277, at_senddmas, expire, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_278(w_eco278, at_senddmas, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_279(w_eco279, at_senddmas, lk_txfsmidle, cur_state[7], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_280(w_eco280, at_senddmas, !lk_txerror, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_281(w_eco281, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4]);
	and _ECO_282(w_eco282, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_283(w_eco283, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_284(w_eco284, !tptx_reset, !lk_txerror, !expire, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_285(w_eco285, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_286(w_eco286, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_287(w_eco287, at_senddmas, lk_txfsmidle, cur_state[11], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_288(w_eco288, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_289(w_eco289, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_290(w_eco290, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_291(w_eco291, at_senddmas, !lk_txerror, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_292(w_eco292, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_293(w_eco293, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_294(w_eco294, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_295(w_eco295, at_senddmas, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_296(w_eco296, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_297(w_eco297, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_298(w_eco298, at_senddmas, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_299(w_eco299, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_300(w_eco300, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_301(w_eco301, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_302(w_eco302, at_senddmas, expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_303(w_eco303, at_senddmas, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_304(w_eco304, at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_305(w_eco305, at_senddmas, !lk_txerror, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_306(w_eco306, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_307(w_eco307, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_308(w_eco308, !tptx_reset, !lk_txerror, !expire, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_309(w_eco309, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_310(w_eco310, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_311(w_eco311, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_312(w_eco312, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_313(w_eco313, at_senddmas, !lk_txerror, cur_state[7], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_314(w_eco314, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_315(w_eco315, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_316(w_eco316, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_317(w_eco317, !at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_318(w_eco318, at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_319(w_eco319, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_320(w_eco320, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_321(w_eco321, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_322(w_eco322, at_senddmas, !lk_txerror, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_323(w_eco323, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_324(w_eco324, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_325(w_eco325, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_326(w_eco326, at_senddmas, expire, cur_state[12], cur_state[13], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_327(w_eco327, at_senddmas, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_328(w_eco328, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_329(w_eco329, at_senddmas, expire, cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_330(w_eco330, at_senddmas, expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_331(w_eco331, at_senddmas, expire, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_332(w_eco332, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_333(w_eco333, at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_334(w_eco334, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4]);
	and _ECO_335(w_eco335, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_336(w_eco336, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_337(w_eco337, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_338(w_eco338, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_339(w_eco339, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_340(w_eco340, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_341(w_eco341, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_342(w_eco342, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_343(w_eco343, !at_senddmas, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_344(w_eco344, !at_senddmas, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_345(w_eco345, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_346(w_eco346, at_senddmas, lk_txfsmidle, cur_state[7], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_347(w_eco347, at_senddmas, !lk_txerror, !cur_state[12], cur_state[14], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_348(w_eco348, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_349(w_eco349, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_350(w_eco350, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_351(w_eco351, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_352(w_eco352, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_353(w_eco353, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_354(w_eco354, !at_senddmas, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_355(w_eco355, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_356(w_eco356, at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_357(w_eco357, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_358(w_eco358, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_359(w_eco359, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_360(w_eco360, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_361(w_eco361, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_362(w_eco362, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_363(w_eco363, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_364(w_eco364, at_senddmas, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_365(w_eco365, at_senddmas, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_366(w_eco366, !at_senddmas, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_367(w_eco367, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_368(w_eco368, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_369(w_eco369, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_370(w_eco370, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_371(w_eco371, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_372(w_eco372, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_373(w_eco373, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_374(w_eco374, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_375(w_eco375, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_376(w_eco376, !at_senddmas, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_377(w_eco377, !at_senddmas, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_378(w_eco378, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_379(w_eco379, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_380(w_eco380, at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[14], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_381(w_eco381, at_senddmas, !lk_txerror, !cur_state[12], cur_state[13], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_382(w_eco382, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_383(w_eco383, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_384(w_eco384, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_385(w_eco385, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_386(w_eco386, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_387(w_eco387, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_388(w_eco388, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_389(w_eco389, at_senddmas, !lk_txerror, !cur_state[8], cur_state[10], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_390(w_eco390, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_391(w_eco391, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_392(w_eco392, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_393(w_eco393, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_394(w_eco394, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_395(w_eco395, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_396(w_eco396, at_senddmas, expire, cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_397(w_eco397, at_senddmas, expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_398(w_eco398, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_399(w_eco399, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_400(w_eco400, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_401(w_eco401, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_402(w_eco402, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_403(w_eco403, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_404(w_eco404, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_405(w_eco405, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_406(w_eco406, !at_senddmas, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_407(w_eco407, !at_senddmas, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_408(w_eco408, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_409(w_eco409, at_senddmas, lk_txfsmidle, !cur_state[12], cur_state[13], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_410(w_eco410, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_411(w_eco411, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_412(w_eco412, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_413(w_eco413, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_414(w_eco414, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_415(w_eco415, !at_senddmas, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_416(w_eco416, !at_senddmas, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_417(w_eco417, at_senddmas, lk_txfsmidle, !cur_state[8], cur_state[10], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_418(w_eco418, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_419(w_eco419, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_420(w_eco420, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_421(w_eco421, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_422(w_eco422, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_423(w_eco423, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_424(w_eco424, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_425(w_eco425, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_426(w_eco426, !at_senddmas, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_427(w_eco427, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_428(w_eco428, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_429(w_eco429, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_430(w_eco430, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_431(w_eco431, !at_senddmas, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_432(w_eco432, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_433(w_eco433, !at_senddmas, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_434(w_eco434, !at_senddmas, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_435(w_eco435, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_436(w_eco436, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_437(w_eco437, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_438(w_eco438, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_439(w_eco439, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_440(w_eco440, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_441(w_eco441, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_442(w_eco442, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_443(w_eco443, at_senddmas, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_444(w_eco444, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_445(w_eco445, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_446(w_eco446, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_447(w_eco447, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	or _ECO_448(w_eco448, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447);
	xor _ECO_out2(next_state[4], sub_wire2, w_eco448);
	and _ECO_449(w_eco449, !lk_txerror, expire, !cur_state[0], at_sendreg);
	and _ECO_450(w_eco450, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_451(w_eco451, !r2t_rxempty, cur_state[0], !at_sendpios, at_sendreg);
	and _ECO_452(w_eco452, lk_txfsmidle, expire, !cur_state[0], at_sendreg);
	and _ECO_453(w_eco453, tptx_reset, at_sendreg);
	and _ECO_454(w_eco454, !lk_txerror, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_455(w_eco455, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_456(w_eco456, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_457(w_eco457, lk_txfsmidle, r2t_rxempty, cur_state[0], at_sendpios, at_sendreg);
	and _ECO_458(w_eco458, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_459(w_eco459, !lk_txfsmidle, cur_state[0], !at_sendpios, at_sendreg);
	and _ECO_460(w_eco460, cur_state[11], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_461(w_eco461, expire, cur_state[11], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_462(w_eco462, lk_txfsmidle, cur_state[11], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_463(w_eco463, !tptx_reset, !lk_txerror, !expire, cur_state[11], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_464(w_eco464, !cur_state[1], !cur_state[2], at_sendreg);
	and _ECO_465(w_eco465, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_466(w_eco466, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_467(w_eco467, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_468(w_eco468, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_469(w_eco469, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_470(w_eco470, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_471(w_eco471, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_472(w_eco472, !tptx_reset, !expire, cur_state[3], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_473(w_eco473, !tptx_reset, !lk_txerror, !expire, !cur_state[3], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_474(w_eco474, !lk_txerror, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_475(w_eco475, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_476(w_eco476, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_477(w_eco477, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_478(w_eco478, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_479(w_eco479, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_480(w_eco480, expire, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_481(w_eco481, !lk_txerror, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_482(w_eco482, !tptx_reset, !lk_txerror, !expire, cur_state[7], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_483(w_eco483, !lk_txfsmidle, lk_txerror, !expire, cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_484(w_eco484, lk_txfsmidle, !tptx_reset, !expire, !cur_state[3], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_485(w_eco485, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_486(w_eco486, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_487(w_eco487, !tptx_reset, !expire, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_488(w_eco488, !lk_txerror, cur_state[11], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_489(w_eco489, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_490(w_eco490, lk_txfsmidle, !cur_state[8], cur_state[9], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_491(w_eco491, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_492(w_eco492, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_493(w_eco493, cur_state[7], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_494(w_eco494, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_495(w_eco495, expire, cur_state[7], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_496(w_eco496, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_497(w_eco497, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_498(w_eco498, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_499(w_eco499, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_500(w_eco500, expire, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_501(w_eco501, lk_txfsmidle, cur_state[7], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_502(w_eco502, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_503(w_eco503, !lk_txerror, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_504(w_eco504, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_505(w_eco505, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_506(w_eco506, !tptx_reset, !expire, cur_state[7], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_507(w_eco507, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_508(w_eco508, lk_txfsmidle, cur_state[11], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_509(w_eco509, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_510(w_eco510, !lk_txerror, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_511(w_eco511, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_512(w_eco512, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_513(w_eco513, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_514(w_eco514, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_515(w_eco515, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_516(w_eco516, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_517(w_eco517, expire, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_518(w_eco518, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_519(w_eco519, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_520(w_eco520, expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_521(w_eco521, lk_txfsmidle, !cur_state[12], cur_state[14], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_522(w_eco522, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_523(w_eco523, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_524(w_eco524, !lk_txerror, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_525(w_eco525, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_526(w_eco526, !lk_txfsmidle, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_527(w_eco527, !tptx_reset, !expire, cur_state[7], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_528(w_eco528, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_529(w_eco529, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_530(w_eco530, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_531(w_eco531, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_532(w_eco532, !lk_txerror, cur_state[7], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_533(w_eco533, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_534(w_eco534, !lk_txfsmidle, lk_txerror, !expire, cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_535(w_eco535, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_536(w_eco536, lk_txfsmidle, !cur_state[8], cur_state[9], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_537(w_eco537, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_538(w_eco538, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_539(w_eco539, !lk_txerror, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_540(w_eco540, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_541(w_eco541, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_542(w_eco542, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_543(w_eco543, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_544(w_eco544, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_545(w_eco545, expire, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_546(w_eco546, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_547(w_eco547, expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_548(w_eco548, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[0], at_sendreg);
	and _ECO_549(w_eco549, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_550(w_eco550, expire, !cur_state[8], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_551(w_eco551, lk_txfsmidle, !cur_state[12], cur_state[13], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_552(w_eco552, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_553(w_eco553, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_554(w_eco554, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_555(w_eco555, lk_txfsmidle, cur_state[7], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_556(w_eco556, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_557(w_eco557, !lk_txerror, !cur_state[12], cur_state[14], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_558(w_eco558, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_559(w_eco559, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_560(w_eco560, lk_txfsmidle, !cur_state[8], cur_state[10], cur_state[3], cur_state[4], !cur_state[0], at_sendreg);
	and _ECO_561(w_eco561, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_562(w_eco562, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_563(w_eco563, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_564(w_eco564, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_565(w_eco565, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_566(w_eco566, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_567(w_eco567, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_568(w_eco568, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_569(w_eco569, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_570(w_eco570, expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_571(w_eco571, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_572(w_eco572, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_573(w_eco573, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_574(w_eco574, lk_txfsmidle, !cur_state[12], cur_state[14], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_575(w_eco575, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_576(w_eco576, !lk_txerror, !cur_state[12], cur_state[13], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_577(w_eco577, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_578(w_eco578, !lk_txfsmidle, lk_txerror, !expire, !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_579(w_eco579, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_580(w_eco580, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_581(w_eco581, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_582(w_eco582, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_583(w_eco583, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_584(w_eco584, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_585(w_eco585, !lk_txerror, !cur_state[8], cur_state[10], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_586(w_eco586, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_587(w_eco587, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_588(w_eco588, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_589(w_eco589, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_590(w_eco590, expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_591(w_eco591, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_592(w_eco592, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_593(w_eco593, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_594(w_eco594, expire, !cur_state[8], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_595(w_eco595, lk_txfsmidle, !cur_state[12], cur_state[13], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_596(w_eco596, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_597(w_eco597, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_598(w_eco598, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_599(w_eco599, lk_txfsmidle, !cur_state[8], cur_state[10], cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_600(w_eco600, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_601(w_eco601, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_602(w_eco602, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_603(w_eco603, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_604(w_eco604, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_605(w_eco605, !lk_txfsmidle, lk_txerror, cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_606(w_eco606, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_607(w_eco607, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, !at_sendreg);
	and _ECO_608(w_eco608, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_609(w_eco609, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_610(w_eco610, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_611(w_eco611, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_612(w_eco612, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, !at_sendreg);
	and _ECO_613(w_eco613, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_614(w_eco614, !lk_txfsmidle, lk_txerror, cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_615(w_eco615, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_616(w_eco616, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	or _ECO_617(w_eco617, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616);
	xor _ECO_out3(next_state[3], sub_wire3, w_eco617);
	and _ECO_618(w_eco618, at_senddmas, at_sendbista, cur_state[0], !at_sendreg);
	and _ECO_619(w_eco619, !at_sendbista, !r2t_rxempty, cur_state[0], at_sendreg);
	and _ECO_620(w_eco620, !at_sendbista, !lk_txfsmidle, cur_state[0], at_sendreg);
	and _ECO_621(w_eco621, at_sendbista, !lk_txerror, expire, !cur_state[0], !at_sendreg);
	and _ECO_622(w_eco622, !at_sendbista, !lk_txerror, expire, !cur_state[0], at_sendreg);
	and _ECO_623(w_eco623, at_sendbista, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_624(w_eco624, !at_sendbista, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_625(w_eco625, at_sendbista, tptx_reset, !at_sendreg);
	and _ECO_626(w_eco626, !at_sendbista, tptx_reset, at_sendreg);
	and _ECO_627(w_eco627, at_sendbista, cur_state[11], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_628(w_eco628, !at_sendbista, cur_state[11], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_629(w_eco629, at_sendbista, lk_txfsmidle, expire, !cur_state[0], !at_sendreg);
	and _ECO_630(w_eco630, !at_sendbista, lk_txfsmidle, expire, !cur_state[0], at_sendreg);
	and _ECO_631(w_eco631, !at_sendbista, !tptx_reset, !lk_txerror, !expire, cur_state[3], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_632(w_eco632, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1]);
	and _ECO_633(w_eco633, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_634(w_eco634, at_sendbista, cur_state[0], !cur_state[1], !cur_state[2], !at_sendreg);
	and _ECO_635(w_eco635, !at_sendbista, !cur_state[1], !cur_state[2], at_sendreg);
	and _ECO_636(w_eco636, !tptx_reset, !lk_txerror, !expire, cur_state[3], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_637(w_eco637, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, cur_state[3], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_638(w_eco638, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_639(w_eco639, at_sendbista, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_640(w_eco640, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2]);
	and _ECO_641(w_eco641, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_642(w_eco642, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_643(w_eco643, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_644(w_eco644, !at_senddmaa, at_sendbista, !r2t_rxempty, cur_state[0], !at_sendpios, !at_sendreg);
	and _ECO_645(w_eco645, at_sendbista, expire, !cur_state[1], !cur_state[2], !at_sendreg);
	and _ECO_646(w_eco646, lk_txfsmidle, !tptx_reset, !expire, cur_state[3], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_647(w_eco647, at_sendbista, cur_state[7], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_648(w_eco648, !at_sendbista, !tptx_reset, !expire, cur_state[3], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_649(w_eco649, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1]);
	and _ECO_650(w_eco650, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_651(w_eco651, at_sendbista, !lk_txerror, !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_652(w_eco652, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_653(w_eco653, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_654(w_eco654, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_655(w_eco655, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_656(w_eco656, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_657(w_eco657, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_658(w_eco658, !at_senddmaa, at_sendbista, !lk_txfsmidle, cur_state[0], !at_sendpios, !at_sendreg);
	and _ECO_659(w_eco659, !at_sendbista, cur_state[7], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_660(w_eco660, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_661(w_eco661, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2]);
	and _ECO_662(w_eco662, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1]);
	and _ECO_663(w_eco663, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_664(w_eco664, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_665(w_eco665, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_666(w_eco666, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_667(w_eco667, at_sendbista, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_668(w_eco668, !at_sendbista, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_669(w_eco669, at_sendbista, lk_txfsmidle, !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_670(w_eco670, !at_sendbista, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_671(w_eco671, !at_sendbista, !lk_txerror, cur_state[11], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_672(w_eco672, !at_sendbista, !tptx_reset, !lk_txerror, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_673(w_eco673, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_674(w_eco674, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_675(w_eco675, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_676(w_eco676, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_677(w_eco677, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_678(w_eco678, at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], cur_state[0], !at_sendreg);
	and _ECO_679(w_eco679, !at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_680(w_eco680, at_sendbista, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_681(w_eco681, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_682(w_eco682, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2]);
	and _ECO_683(w_eco683, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_684(w_eco684, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_685(w_eco685, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_686(w_eco686, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_687(w_eco687, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_688(w_eco688, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_689(w_eco689, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_690(w_eco690, !at_sendbista, lk_txfsmidle, cur_state[11], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_691(w_eco691, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_692(w_eco692, !at_sendbista, !tptx_reset, !expire, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_693(w_eco693, !at_sendbista, expire, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_694(w_eco694, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_695(w_eco695, !tptx_reset, !lk_txerror, !expire, !cur_state[4], !cur_state[6], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_696(w_eco696, !at_sendbista, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_697(w_eco697, !at_sendbista, !lk_txerror, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_698(w_eco698, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_699(w_eco699, at_sendbista, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_700(w_eco700, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_701(w_eco701, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_702(w_eco702, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_703(w_eco703, at_sendbista, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_704(w_eco704, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_705(w_eco705, !at_sendbista, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_706(w_eco706, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_707(w_eco707, !at_sendbista, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_708(w_eco708, !at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_709(w_eco709, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_710(w_eco710, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_711(w_eco711, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_712(w_eco712, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_713(w_eco713, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_714(w_eco714, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_715(w_eco715, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_716(w_eco716, at_sendbista, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_717(w_eco717, !at_sendbista, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_718(w_eco718, !at_sendbista, !lk_txerror, cur_state[7], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_719(w_eco719, !at_sendbista, !tptx_reset, !lk_txerror, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_720(w_eco720, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], !cur_state[6], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_721(w_eco721, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_722(w_eco722, !at_sendbista, lk_txfsmidle, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_723(w_eco723, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_724(w_eco724, !at_sendbista, expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_725(w_eco725, !at_sendbista, lk_txfsmidle, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_726(w_eco726, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_727(w_eco727, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_728(w_eco728, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_729(w_eco729, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_730(w_eco730, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_731(w_eco731, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_732(w_eco732, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_733(w_eco733, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_734(w_eco734, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_735(w_eco735, at_sendbista, expire, !cur_state[12], !cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], !at_sendreg);
	and _ECO_736(w_eco736, at_sendbista, lk_txfsmidle, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !at_sendreg);
	and _ECO_737(w_eco737, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_738(w_eco738, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_739(w_eco739, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_740(w_eco740, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_741(w_eco741, at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], !at_sendreg);
	and _ECO_742(w_eco742, !at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_743(w_eco743, at_sendbista, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_744(w_eco744, !at_sendbista, lk_txfsmidle, cur_state[7], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_745(w_eco745, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_746(w_eco746, !at_sendbista, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_747(w_eco747, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_748(w_eco748, !at_sendbista, expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_749(w_eco749, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_750(w_eco750, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_751(w_eco751, !at_sendbista, !lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_752(w_eco752, at_sendbista, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_753(w_eco753, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_754(w_eco754, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_755(w_eco755, at_sendbista, !lk_txfsmidle, lk_txerror, !expire, cur_state[12], !cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_756(w_eco756, !at_sendbista, !lk_txfsmidle, lk_txerror, cur_state[12], !cur_state[8], !cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_757(w_eco757, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_758(w_eco758, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_759(w_eco759, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_760(w_eco760, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_761(w_eco761, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_762(w_eco762, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_763(w_eco763, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_764(w_eco764, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_765(w_eco765, at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !cur_state[1], !cur_state[2], !at_sendreg);
	and _ECO_766(w_eco766, at_sendbista, !cur_state[12], !cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_767(w_eco767, at_sendbista, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_768(w_eco768, !at_sendbista, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_769(w_eco769, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_770(w_eco770, !at_sendbista, lk_txfsmidle, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_771(w_eco771, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_772(w_eco772, !at_sendbista, !lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_773(w_eco773, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_774(w_eco774, !at_sendbista, expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_775(w_eco775, !at_sendbista, !lk_txfsmidle, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_776(w_eco776, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_777(w_eco777, !at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_778(w_eco778, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_779(w_eco779, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_780(w_eco780, !at_sendbista, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0], at_sendreg);
	and _ECO_781(w_eco781, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_782(w_eco782, !at_sendbista, !lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_783(w_eco783, !at_sendbista, !tptx_reset, !lk_txerror, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_784(w_eco784, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_785(w_eco785, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_786(w_eco786, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_787(w_eco787, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_788(w_eco788, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_789(w_eco789, !at_sendbista, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_790(w_eco790, !at_sendbista, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_791(w_eco791, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_792(w_eco792, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_793(w_eco793, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_794(w_eco794, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_795(w_eco795, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_796(w_eco796, at_sendbista, expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !at_sendreg);
	and _ECO_797(w_eco797, at_sendbista, lk_txfsmidle, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !at_sendreg);
	and _ECO_798(w_eco798, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_799(w_eco799, !at_sendbista, lk_txfsmidle, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_800(w_eco800, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_801(w_eco801, !at_sendbista, expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_802(w_eco802, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_803(w_eco803, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_804(w_eco804, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_805(w_eco805, !at_sendbista, lk_txfsmidle, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], cur_state[6], !cur_state[0], at_sendreg);
	and _ECO_806(w_eco806, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_807(w_eco807, !at_sendbista, !lk_txfsmidle, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_808(w_eco808, !lk_txfsmidle, !tptx_reset, lk_txerror, !expire, cur_state[12], !cur_state[8], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_809(w_eco809, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_810(w_eco810, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_811(w_eco811, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_812(w_eco812, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_813(w_eco813, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_814(w_eco814, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_815(w_eco815, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_816(w_eco816, !at_sendbista, !lk_txfsmidle, expire, !cur_state[8], !cur_state[10], !cur_state[3], cur_state[4], at_sendreg);
	and _ECO_817(w_eco817, !at_sendbista, !lk_txfsmidle, expire, !cur_state[8], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_818(w_eco818, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_819(w_eco819, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_820(w_eco820, at_sendbista, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[1], !cur_state[2], !at_sendreg);
	and _ECO_821(w_eco821, at_sendbista, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_822(w_eco822, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_823(w_eco823, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !at_sendreg);
	and _ECO_824(w_eco824, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_825(w_eco825, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendreg);
	and _ECO_826(w_eco826, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_827(w_eco827, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_828(w_eco828, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_829(w_eco829, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_830(w_eco830, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], at_sendreg);
	and _ECO_831(w_eco831, at_sendbista, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_832(w_eco832, !at_sendbista, !lk_txfsmidle, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], at_sendreg);
	and _ECO_833(w_eco833, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !at_sendreg);
	and _ECO_834(w_eco834, !at_senddmas, at_senddmaa, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendreg);
	and _ECO_835(w_eco835, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios, at_sendreg);
	and _ECO_836(w_eco836, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_837(w_eco837, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], !at_sendpios, at_sendreg);
	and _ECO_838(w_eco838, !lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], at_sendreg);
	and _ECO_839(w_eco839, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	and _ECO_840(w_eco840, !at_sendbista, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !cur_state[1], !at_sendreg);
	and _ECO_841(w_eco841, !at_senddmas, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios, at_sendreg);
	and _ECO_842(w_eco842, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], !at_sendpios, at_sendreg);
	and _ECO_843(w_eco843, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], cur_state[2], !at_sendreg);
	or _ECO_844(w_eco844, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843);
	xor _ECO_out4(next_state[2], sub_wire4, w_eco844);
	and _ECO_845(w_eco845, !at_sendbista, !r2t_rxempty, !tptx_reset, cur_state[0]);
	and _ECO_846(w_eco846, at_senddmas, at_sendbista, lk_txfsmidle, r2t_rxempty, cur_state[0]);
	and _ECO_847(w_eco847, at_sendbista, tptx_reset);
	and _ECO_848(w_eco848, !at_sendbista, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1]);
	and _ECO_849(w_eco849, at_sendbista, r2t_rxempty, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_850(w_eco850, at_sendbista, r2t_rxempty, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_851(w_eco851, at_sendbista, r2t_rxempty, cur_state[11], !cur_state[3], cur_state[4]);
	and _ECO_852(w_eco852, !at_senddmas, at_senddmaa, at_sendbista, !lk_txfsmidle, r2t_rxempty, cur_state[0]);
	and _ECO_853(w_eco853, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1]);
	and _ECO_854(w_eco854, !at_sendbista, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2]);
	and _ECO_855(w_eco855, at_sendbista, r2t_rxempty, !lk_txerror, !cur_state[0], !r2t_waittxid);
	and _ECO_856(w_eco856, at_sendbista, txtimeout, !lk_txerror, cur_state[3], !cur_state[0], cur_state[1]);
	and _ECO_857(w_eco857, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, cur_state[3]);
	and _ECO_858(w_eco858, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1]);
	and _ECO_859(w_eco859, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[8], cur_state[9], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_860(w_eco860, at_sendbista, r2t_rxempty, cur_state[0], !cur_state[1], !cur_state[2]);
	and _ECO_861(w_eco861, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2]);
	and _ECO_862(w_eco862, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_863(w_eco863, at_sendbista, lk_txfsmidle, r2t_rxempty, !cur_state[0], !r2t_waittxid);
	and _ECO_864(w_eco864, at_sendbista, txtimeout, !lk_txerror, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_865(w_eco865, at_sendbista, lk_txfsmidle, !lk_txerror, cur_state[3], !cur_state[0], cur_state[1]);
	and _ECO_866(w_eco866, !at_sendbista, !r2t_rxempty, !tptx_reset, cur_state[11], !cur_state[3], cur_state[4]);
	and _ECO_867(w_eco867, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, cur_state[3], !cur_state[0], r2t_waittxid);
	and _ECO_868(w_eco868, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, cur_state[3]);
	and _ECO_869(w_eco869, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1]);
	and _ECO_870(w_eco870, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2]);
	and _ECO_871(w_eco871, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1]);
	and _ECO_872(w_eco872, at_sendbista, txtimeout, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_873(w_eco873, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5]);
	and _ECO_874(w_eco874, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_875(w_eco875, !at_senddmas, !r2t_rxempty, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_876(w_eco876, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_877(w_eco877, at_sendbista, lk_txfsmidle, cur_state[3], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_878(w_eco878, !lk_txfsmidle, !txtimeout, !tptx_reset, lk_txerror, cur_state[3], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_879(w_eco879, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !expire, cur_state[3], !r2t_waittxid);
	and _ECO_880(w_eco880, at_sendbista, lk_txfsmidle, r2t_rxempty, !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_881(w_eco881, at_sendbista, r2t_rxempty, !cur_state[1], !cur_state[2], !r2t_waittxid);
	and _ECO_882(w_eco882, at_sendbista, lk_txfsmidle, cur_state[3], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_883(w_eco883, at_sendbista, lk_txfsmidle, cur_state[3], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_884(w_eco884, at_sendbista, !lk_txerror, cur_state[3], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_885(w_eco885, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_886(w_eco886, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, cur_state[3], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_887(w_eco887, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[1], !cur_state[2]);
	and _ECO_888(w_eco888, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, cur_state[3], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_889(w_eco889, lk_txfsmidle, !tptx_reset, !expire, cur_state[3], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_890(w_eco890, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2]);
	and _ECO_891(w_eco891, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_892(w_eco892, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1]);
	and _ECO_893(w_eco893, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2]);
	and _ECO_894(w_eco894, at_sendbista, txtimeout, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_895(w_eco895, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1]);
	and _ECO_896(w_eco896, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], r2t_waittxid);
	and _ECO_897(w_eco897, at_sendbista, r2t_rxempty, cur_state[7], !cur_state[3], cur_state[4]);
	and _ECO_898(w_eco898, !at_senddmas, !lk_txfsmidle, !tptx_reset, cur_state[3], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_899(w_eco899, !at_senddmaa, at_sendbista, lk_txfsmidle, r2t_rxempty, cur_state[0], !at_sendpios, at_sendreg);
	and _ECO_900(w_eco900, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_901(w_eco901, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_902(w_eco902, at_sendbista, lk_txfsmidle, r2t_rxempty, !lk_txerror, !cur_state[0], cur_state[2]);
	and _ECO_903(w_eco903, at_sendbista, r2t_rxempty, !lk_txerror, !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_904(w_eco904, at_sendbista, lk_txfsmidle, !lk_txerror, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_905(w_eco905, at_sendbista, !lk_txerror, cur_state[3], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_906(w_eco906, at_sendbista, !lk_txerror, cur_state[3], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_907(w_eco907, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_908(w_eco908, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_909(w_eco909, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, cur_state[3], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_910(w_eco910, !at_sendbista, !tptx_reset, cur_state[3], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_911(w_eco911, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, cur_state[3], cur_state[2], r2t_waittxid);
	and _ECO_912(w_eco912, !at_sendbista, !r2t_rxempty, !tptx_reset, cur_state[7], !cur_state[3], cur_state[4]);
	and _ECO_913(w_eco913, lk_txfsmidle, !tptx_reset, !expire, cur_state[3], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_914(w_eco914, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, cur_state[3], cur_state[1], !r2t_waittxid);
	and _ECO_915(w_eco915, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, cur_state[3], !cur_state[0], cur_state[2]);
	and _ECO_916(w_eco916, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, cur_state[3], cur_state[1], !cur_state[2]);
	and _ECO_917(w_eco917, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, cur_state[3], cur_state[2], !r2t_waittxid);
	and _ECO_918(w_eco918, at_sendbista, r2t_rxempty, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_919(w_eco919, !at_senddmas, at_sendbista, !lk_txfsmidle, r2t_rxempty, cur_state[0], at_sendpios);
	and _ECO_920(w_eco920, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[5], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_921(w_eco921, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2]);
	and _ECO_922(w_eco922, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_923(w_eco923, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_924(w_eco924, !lk_txfsmidle, !txtimeout, !tptx_reset, lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_925(w_eco925, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_926(w_eco926, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_927(w_eco927, at_sendbista, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_928(w_eco928, at_sendbista, txtimeout, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_929(w_eco929, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_930(w_eco930, !at_sendbista, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_931(w_eco931, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_932(w_eco932, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, !cur_state[8], cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_933(w_eco933, r2t_rxempty, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_934(w_eco934, at_sendbista, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_935(w_eco935, r2t_rxempty, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_936(w_eco936, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_937(w_eco937, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_938(w_eco938, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_939(w_eco939, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_940(w_eco940, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_941(w_eco941, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], r2t_waittxid);
	and _ECO_942(w_eco942, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[4], cur_state[6], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_943(w_eco943, at_sendbista, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_944(w_eco944, at_sendbista, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_945(w_eco945, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_946(w_eco946, !lk_txfsmidle, !txtimeout, !tptx_reset, lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_947(w_eco947, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_948(w_eco948, at_sendbista, lk_txfsmidle, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_949(w_eco949, at_sendbista, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_950(w_eco950, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_951(w_eco951, !at_sendbista, !tptx_reset, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_952(w_eco952, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[4], cur_state[5], cur_state[2], r2t_waittxid);
	and _ECO_953(w_eco953, lk_txfsmidle, !tptx_reset, !expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_954(w_eco954, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_955(w_eco955, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], cur_state[1], !r2t_waittxid);
	and _ECO_956(w_eco956, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], cur_state[1], !cur_state[2]);
	and _ECO_957(w_eco957, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[4], cur_state[5], cur_state[2], !r2t_waittxid);
	and _ECO_958(w_eco958, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_959(w_eco959, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_960(w_eco960, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_961(w_eco961, r2t_rxempty, !tptx_reset, !expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_962(w_eco962, at_sendbista, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_963(w_eco963, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[14], !cur_state[8], cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_964(w_eco964, r2t_rxempty, !tptx_reset, !expire, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_965(w_eco965, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_966(w_eco966, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_967(w_eco967, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_968(w_eco968, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4]);
	and _ECO_969(w_eco969, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_970(w_eco970, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_971(w_eco971, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_972(w_eco972, at_sendbista, lk_txfsmidle, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_973(w_eco973, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_974(w_eco974, at_sendbista, !lk_txfsmidle, !txtimeout, r2t_rxempty, lk_txerror, cur_state[12], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_975(w_eco975, !lk_txfsmidle, !txtimeout, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_976(w_eco976, at_sendbista, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_977(w_eco977, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, !expire, cur_state[8], cur_state[4], !r2t_waittxid);
	and _ECO_978(w_eco978, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_979(w_eco979, !at_sendbista, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], r2t_waittxid);
	and _ECO_980(w_eco980, at_sendbista, r2t_rxempty, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_981(w_eco981, at_sendbista, txtimeout, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_982(w_eco982, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_983(w_eco983, at_sendbista, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_984(w_eco984, at_sendbista, !lk_txerror, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_985(w_eco985, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_986(w_eco986, !at_sendbista, !tptx_reset, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_987(w_eco987, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[4], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_988(w_eco988, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_989(w_eco989, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_990(w_eco990, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_991(w_eco991, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_992(w_eco992, txtimeout, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_993(w_eco993, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_994(w_eco994, at_sendbista, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_995(w_eco995, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[13], !cur_state[8], cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_996(w_eco996, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_997(w_eco997, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_998(w_eco998, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_999(w_eco999, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_1000(w_eco1000, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1001(w_eco1001, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1002(w_eco1002, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1003(w_eco1003, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_1004(w_eco1004, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_1005(w_eco1005, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_1006(w_eco1006, at_sendbista, lk_txfsmidle, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1007(w_eco1007, at_sendbista, lk_txfsmidle, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1008(w_eco1008, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1009(w_eco1009, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1010(w_eco1010, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1011(w_eco1011, at_sendbista, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1012(w_eco1012, at_sendbista, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1013(w_eco1013, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1014(w_eco1014, !at_sendbista, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1015(w_eco1015, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[2], r2t_waittxid);
	and _ECO_1016(w_eco1016, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1017(w_eco1017, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[12], cur_state[8], !cur_state[3], cur_state[4], !r2t_waittxid);
	and _ECO_1018(w_eco1018, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], r2t_waittxid);
	and _ECO_1019(w_eco1019, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1020(w_eco1020, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1021(w_eco1021, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_1022(w_eco1022, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1023(w_eco1023, r2t_rxempty, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1024(w_eco1024, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1025(w_eco1025, txtimeout, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[4], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1026(w_eco1026, at_sendbista, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1027(w_eco1027, at_sendbista, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1028(w_eco1028, !at_sendbista, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1029(w_eco1029, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1030(w_eco1030, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1031(w_eco1031, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1032(w_eco1032, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[14], !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_1033(w_eco1033, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1034(w_eco1034, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_1035(w_eco1035, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_1036(w_eco1036, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1037(w_eco1037, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1038(w_eco1038, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_1039(w_eco1039, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, expire, !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_1040(w_eco1040, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], r2t_waittxid);
	and _ECO_1041(w_eco1041, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_1042(w_eco1042, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1043(w_eco1043, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1044(w_eco1044, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1045(w_eco1045, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1046(w_eco1046, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4]);
	and _ECO_1047(w_eco1047, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1048(w_eco1048, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1049(w_eco1049, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1050(w_eco1050, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1051(w_eco1051, !at_sendbista, !lk_txfsmidle, txtimeout, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1052(w_eco1052, !at_sendbista, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_1053(w_eco1053, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1054(w_eco1054, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1055(w_eco1055, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[1], !cur_state[2]);
	and _ECO_1056(w_eco1056, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1057(w_eco1057, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[4], cur_state[5], !cur_state[0], cur_state[2]);
	and _ECO_1058(w_eco1058, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1059(w_eco1059, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_1060(w_eco1060, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1061(w_eco1061, r2t_rxempty, !tptx_reset, !expire, cur_state[11], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1062(w_eco1062, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[4], !cur_state[6]);
	and _ECO_1063(w_eco1063, at_sendbista, r2t_rxempty, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1064(w_eco1064, at_sendbista, r2t_rxempty, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1065(w_eco1065, at_sendbista, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1066(w_eco1066, at_sendbista, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1067(w_eco1067, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1068(w_eco1068, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1069(w_eco1069, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1070(w_eco1070, !at_sendbista, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[13], !cur_state[8], cur_state[10], !cur_state[3], cur_state[4]);
	and _ECO_1071(w_eco1071, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_1072(w_eco1072, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_1073(w_eco1073, !at_sendbista, !lk_txfsmidle, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1074(w_eco1074, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1075(w_eco1075, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1076(w_eco1076, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1077(w_eco1077, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, cur_state[12], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4]);
	and _ECO_1078(w_eco1078, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1079(w_eco1079, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10]);
	and _ECO_1080(w_eco1080, !at_sendbista, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], r2t_waittxid);
	and _ECO_1081(w_eco1081, at_sendbista, lk_txfsmidle, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1082(w_eco1082, at_sendbista, lk_txfsmidle, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1083(w_eco1083, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1084(w_eco1084, at_sendbista, r2t_rxempty, !cur_state[12], !cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], !r2t_waittxid);
	and _ECO_1085(w_eco1085, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1086(w_eco1086, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1087(w_eco1087, at_sendbista, r2t_rxempty, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1088(w_eco1088, at_sendbista, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1089(w_eco1089, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1090(w_eco1090, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4]);
	and _ECO_1091(w_eco1091, !at_sendbista, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1092(w_eco1092, r2t_rxempty, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1093(w_eco1093, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1094(w_eco1094, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[2], r2t_waittxid);
	and _ECO_1095(w_eco1095, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4]);
	and _ECO_1096(w_eco1096, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_1097(w_eco1097, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1098(w_eco1098, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1099(w_eco1099, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1100(w_eco1100, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1101(w_eco1101, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_1102(w_eco1102, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1103(w_eco1103, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1104(w_eco1104, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1105(w_eco1105, r2t_rxempty, !tptx_reset, !expire, cur_state[7], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1106(w_eco1106, !lk_txfsmidle, txtimeout, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1107(w_eco1107, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1108(w_eco1108, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1109(w_eco1109, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1110(w_eco1110, at_sendbista, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1111(w_eco1111, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1112(w_eco1112, !at_sendbista, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], cur_state[9], !cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1113(w_eco1113, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1114(w_eco1114, at_sendbista, txtimeout, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1115(w_eco1115, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1116(w_eco1116, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1117(w_eco1117, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1118(w_eco1118, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[4], !cur_state[6]);
	and _ECO_1119(w_eco1119, !at_senddmas, at_senddmaa, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1120(w_eco1120, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1], at_sendpios);
	and _ECO_1121(w_eco1121, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1122(w_eco1122, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1123(w_eco1123, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1124(w_eco1124, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1125(w_eco1125, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1126(w_eco1126, !at_sendbista, !tptx_reset, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1127(w_eco1127, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[2], r2t_waittxid);
	and _ECO_1128(w_eco1128, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1129(w_eco1129, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[2], r2t_waittxid);
	and _ECO_1130(w_eco1130, !at_sendbista, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], r2t_waittxid);
	and _ECO_1131(w_eco1131, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1132(w_eco1132, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1133(w_eco1133, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10]);
	and _ECO_1134(w_eco1134, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4], !cur_state[1], !cur_state[2]);
	and _ECO_1135(w_eco1135, at_sendbista, lk_txfsmidle, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1136(w_eco1136, at_sendbista, lk_txfsmidle, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1137(w_eco1137, at_sendbista, r2t_rxempty, !cur_state[12], !cur_state[14], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1138(w_eco1138, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[13], cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1139(w_eco1139, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1140(w_eco1140, at_sendbista, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1141(w_eco1141, at_sendbista, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1142(w_eco1142, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1143(w_eco1143, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1144(w_eco1144, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1145(w_eco1145, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1146(w_eco1146, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[4], !cur_state[6]);
	and _ECO_1147(w_eco1147, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1148(w_eco1148, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_1149(w_eco1149, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1150(w_eco1150, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1151(w_eco1151, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1152(w_eco1152, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1153(w_eco1153, !lk_txfsmidle, txtimeout, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1154(w_eco1154, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1155(w_eco1155, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !r2t_waittxid);
	and _ECO_1156(w_eco1156, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_1157(w_eco1157, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], cur_state[6], cur_state[2], r2t_waittxid);
	and _ECO_1158(w_eco1158, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[14], !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1159(w_eco1159, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1160(w_eco1160, at_sendbista, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1161(w_eco1161, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1162(w_eco1162, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1163(w_eco1163, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[14], !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1164(w_eco1164, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, expire, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1165(w_eco1165, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1166(w_eco1166, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[4], !cur_state[6]);
	and _ECO_1167(w_eco1167, !at_senddmas, !r2t_rxempty, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2], at_sendpios);
	and _ECO_1168(w_eco1168, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1169(w_eco1169, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1170(w_eco1170, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1171(w_eco1171, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1172(w_eco1172, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1173(w_eco1173, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1174(w_eco1174, !at_sendbista, !lk_txfsmidle, txtimeout, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1175(w_eco1175, !at_sendbista, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_1176(w_eco1176, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1177(w_eco1177, txtimeout, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1178(w_eco1178, !at_sendbista, !lk_txfsmidle, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[1], !cur_state[2]);
	and _ECO_1179(w_eco1179, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10]);
	and _ECO_1180(w_eco1180, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1181(w_eco1181, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], !r2t_waittxid);
	and _ECO_1182(w_eco1182, !at_sendbista, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1183(w_eco1183, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], !cur_state[6]);
	and _ECO_1184(w_eco1184, at_sendbista, lk_txfsmidle, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1185(w_eco1185, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1186(w_eco1186, at_sendbista, r2t_rxempty, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], !r2t_waittxid);
	and _ECO_1187(w_eco1187, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1188(w_eco1188, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1189(w_eco1189, at_sendbista, r2t_rxempty, !lk_txerror, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1190(w_eco1190, at_sendbista, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[1], !cur_state[2]);
	and _ECO_1191(w_eco1191, at_sendbista, r2t_rxempty, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1192(w_eco1192, at_sendbista, !lk_txerror, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1193(w_eco1193, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[1], !cur_state[2]);
	and _ECO_1194(w_eco1194, r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1195(w_eco1195, lk_txfsmidle, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1196(w_eco1196, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1197(w_eco1197, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1198(w_eco1198, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[7], cur_state[8], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[2]);
	and _ECO_1199(w_eco1199, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[13], !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1200(w_eco1200, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1201(w_eco1201, !at_sendbista, !r2t_rxempty, !tptx_reset, expire, !cur_state[12], cur_state[13], !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1202(w_eco1202, !at_sendbista, txtimeout, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[4], !cur_state[6]);
	and _ECO_1203(w_eco1203, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1204(w_eco1204, !at_sendbista, !txtimeout, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1205(w_eco1205, !at_sendbista, !tptx_reset, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1206(w_eco1206, !at_sendbista, !lk_txfsmidle, !txtimeout, !tptx_reset, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[2], r2t_waittxid);
	and _ECO_1207(w_eco1207, r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1208(w_eco1208, !at_sendbista, !lk_txfsmidle, txtimeout, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[1]);
	and _ECO_1209(w_eco1209, lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1210(w_eco1210, at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1211(w_eco1211, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], !cur_state[2]);
	and _ECO_1212(w_eco1212, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1213(w_eco1213, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[1], !r2t_waittxid);
	and _ECO_1214(w_eco1214, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, lk_txerror, expire, !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1215(w_eco1215, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, expire, !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1216(w_eco1216, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1217(w_eco1217, !at_sendbista, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1218(w_eco1218, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], !cur_state[6]);
	and _ECO_1219(w_eco1219, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1220(w_eco1220, r2t_rxempty, !tptx_reset, !expire, !cur_state[12], !cur_state[14], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1221(w_eco1221, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1222(w_eco1222, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1223(w_eco1223, at_sendbista, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1224(w_eco1224, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1225(w_eco1225, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1226(w_eco1226, !at_sendbista, lk_txfsmidle, !r2t_rxempty, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[4], !cur_state[6]);
	and _ECO_1227(w_eco1227, !at_sendbista, lk_txfsmidle, !tptx_reset, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1228(w_eco1228, !at_sendbista, !lk_txfsmidle, txtimeout, !tptx_reset, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[2]);
	and _ECO_1229(w_eco1229, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !tptx_reset, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1230(w_eco1230, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1231(w_eco1231, lk_txfsmidle, !tptx_reset, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1232(w_eco1232, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[1], !cur_state[2]);
	and _ECO_1233(w_eco1233, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[2], !r2t_waittxid);
	and _ECO_1234(w_eco1234, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[1], !r2t_waittxid);
	and _ECO_1235(w_eco1235, !at_sendbista, !lk_txfsmidle, txtimeout, !r2t_rxempty, !tptx_reset, !expire, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[4], !cur_state[5], !cur_state[6]);
	and _ECO_1236(w_eco1236, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[1], !cur_state[2]);
	and _ECO_1237(w_eco1237, !at_sendbista, !lk_txfsmidle, !tptx_reset, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[4], cur_state[6], cur_state[2], !r2t_waittxid);
	or _ECO_1238(w_eco1238, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237);
	xor _ECO_out5(next_state[6], sub_wire5, w_eco1238);
	and _ECO_1239(w_eco1239, r2t_rxempty, !expire, cur_state[3], !cur_state[0]);
	and _ECO_1240(w_eco1240, at_senddata, r2t_rxempty, cur_state[0]);
	assign w_eco1241 = tptx_reset;
	and _ECO_1242(w_eco1242, !expire, cur_state[3], !cur_state[0], r2t_waittxid);
	and _ECO_1243(w_eco1243, r2t_rxempty, !expire, !cur_state[4], cur_state[5], !cur_state[0]);
	and _ECO_1244(w_eco1244, r2t_rxempty, !expire, cur_state[10], !cur_state[0]);
	and _ECO_1245(w_eco1245, r2t_rxempty, !expire, cur_state[9], !cur_state[0]);
	and _ECO_1246(w_eco1246, !r2t_rxempty, cur_state[3], cur_state[0], cur_state[1]);
	and _ECO_1247(w_eco1247, lk_txfsmidle, r2t_rxempty, cur_state[0]);
	and _ECO_1248(w_eco1248, r2t_rxempty, !cur_state[1], !cur_state[2]);
	and _ECO_1249(w_eco1249, !r2t_rxempty, cur_state[3], cur_state[0], cur_state[2]);
	and _ECO_1250(w_eco1250, !r2t_rxempty, !expire, cur_state[3], cur_state[1]);
	and _ECO_1251(w_eco1251, !r2t_rxempty, !cur_state[4], cur_state[5], cur_state[0], cur_state[1]);
	and _ECO_1252(w_eco1252, !expire, !cur_state[4], cur_state[5], !cur_state[0], r2t_waittxid);
	and _ECO_1253(w_eco1253, cur_state[3], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1254(w_eco1254, r2t_rxempty, cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_1255(w_eco1255, !r2t_rxempty, !expire, cur_state[3], cur_state[2]);
	and _ECO_1256(w_eco1256, !r2t_rxempty, !cur_state[4], cur_state[5], cur_state[0], cur_state[2]);
	and _ECO_1257(w_eco1257, !r2t_rxempty, !cur_state[4], cur_state[6], cur_state[0], cur_state[1]);
	and _ECO_1258(w_eco1258, !r2t_rxempty, !expire, !cur_state[4], cur_state[5], cur_state[1]);
	and _ECO_1259(w_eco1259, !expire, !cur_state[4], cur_state[6], !cur_state[0], r2t_waittxid);
	and _ECO_1260(w_eco1260, r2t_rxempty, cur_state[11], !cur_state[3], cur_state[4]);
	and _ECO_1261(w_eco1261, at_senddmas, !at_sendbista, r2t_rxempty, cur_state[0]);
	and _ECO_1262(w_eco1262, !r2t_rxempty, !cur_state[4], cur_state[6], cur_state[0], cur_state[2]);
	and _ECO_1263(w_eco1263, !cur_state[4], cur_state[5], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1264(w_eco1264, !r2t_rxempty, !expire, !cur_state[4], cur_state[5], cur_state[2]);
	and _ECO_1265(w_eco1265, !r2t_rxempty, !expire, !cur_state[4], cur_state[6], cur_state[1]);
	and _ECO_1266(w_eco1266, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_1267(w_eco1267, at_senddmaa, !at_sendbista, r2t_rxempty, cur_state[0]);
	and _ECO_1268(w_eco1268, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1269(w_eco1269, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1270(w_eco1270, !cur_state[4], cur_state[6], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1271(w_eco1271, !r2t_rxempty, !expire, !cur_state[4], cur_state[6], cur_state[2]);
	and _ECO_1272(w_eco1272, r2t_rxempty, cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_1273(w_eco1273, r2t_rxempty, cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0]);
	and _ECO_1274(w_eco1274, r2t_rxempty, !expire, cur_state[8], !cur_state[0]);
	and _ECO_1275(w_eco1275, r2t_rxempty, !cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_1276(w_eco1276, r2t_rxempty, cur_state[7], !cur_state[3], cur_state[4]);
	and _ECO_1277(w_eco1277, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1278(w_eco1278, r2t_rxempty, cur_state[11], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1279(w_eco1279, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1280(w_eco1280, !expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1281(w_eco1281, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1282(w_eco1282, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1283(w_eco1283, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], cur_state[4]);
	and _ECO_1284(w_eco1284, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1285(w_eco1285, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1286(w_eco1286, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_1287(w_eco1287, !expire, !cur_state[4], cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1288(w_eco1288, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_1289(w_eco1289, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1290(w_eco1290, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[1]);
	and _ECO_1291(w_eco1291, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1292(w_eco1292, r2t_rxempty, cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0]);
	and _ECO_1293(w_eco1293, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], !cur_state[0], r2t_waittxid);
	and _ECO_1294(w_eco1294, txtimeout, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_1295(w_eco1295, r2t_rxempty, !cur_state[12], cur_state[13], !cur_state[3], cur_state[4]);
	and _ECO_1296(w_eco1296, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1297(w_eco1297, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[1]);
	and _ECO_1298(w_eco1298, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[1]);
	and _ECO_1299(w_eco1299, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[0], cur_state[2]);
	and _ECO_1300(w_eco1300, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1301(w_eco1301, r2t_rxempty, !cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_1302(w_eco1302, r2t_rxempty, cur_state[7], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1303(w_eco1303, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1304(w_eco1304, r2t_rxempty, !cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[0]);
	and _ECO_1305(w_eco1305, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], !cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1306(w_eco1306, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1307(w_eco1307, txtimeout, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1308(w_eco1308, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], cur_state[0], cur_state[2]);
	and _ECO_1309(w_eco1309, r2t_rxempty, !expire, cur_state[12], !cur_state[0]);
	and _ECO_1310(w_eco1310, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1311(w_eco1311, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[1]);
	and _ECO_1312(w_eco1312, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1313(w_eco1313, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1314(w_eco1314, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1315(w_eco1315, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[2]);
	and _ECO_1316(w_eco1316, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1317(w_eco1317, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_1318(w_eco1318, !r2t_rxempty, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[1]);
	and _ECO_1319(w_eco1319, txtimeout, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_1320(w_eco1320, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1321(w_eco1321, r2t_rxempty, !cur_state[12], cur_state[14], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1322(w_eco1322, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1323(w_eco1323, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], !cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1324(w_eco1324, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1325(w_eco1325, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1326(w_eco1326, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1327(w_eco1327, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1328(w_eco1328, txtimeout, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1329(w_eco1329, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[1]);
	and _ECO_1330(w_eco1330, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_1331(w_eco1331, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1332(w_eco1332, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], r2t_waittxid);
	and _ECO_1333(w_eco1333, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1334(w_eco1334, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], r2t_waittxid);
	and _ECO_1335(w_eco1335, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[2]);
	and _ECO_1336(w_eco1336, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1337(w_eco1337, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], r2t_waittxid);
	and _ECO_1338(w_eco1338, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1339(w_eco1339, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[1]);
	and _ECO_1340(w_eco1340, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1341(w_eco1341, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], r2t_waittxid);
	and _ECO_1342(w_eco1342, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1343(w_eco1343, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1344(w_eco1344, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1345(w_eco1345, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_1346(w_eco1346, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], !cur_state[0], r2t_waittxid);
	and _ECO_1347(w_eco1347, !r2t_rxempty, !expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[2]);
	and _ECO_1348(w_eco1348, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[1]);
	and _ECO_1349(w_eco1349, r2t_rxempty, !cur_state[12], cur_state[13], !cur_state[3], !cur_state[5], !cur_state[6]);
	and _ECO_1350(w_eco1350, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1351(w_eco1351, r2t_rxempty, !cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[0]);
	and _ECO_1352(w_eco1352, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1353(w_eco1353, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1354(w_eco1354, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1355(w_eco1355, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1356(w_eco1356, txtimeout, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1357(w_eco1357, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[9], !cur_state[0], cur_state[2]);
	and _ECO_1358(w_eco1358, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1359(w_eco1359, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1360(w_eco1360, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1361(w_eco1361, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1362(w_eco1362, !expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[2], r2t_waittxid);
	and _ECO_1363(w_eco1363, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[1]);
	and _ECO_1364(w_eco1364, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1365(w_eco1365, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1366(w_eco1366, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[1]);
	and _ECO_1367(w_eco1367, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1368(w_eco1368, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], cur_state[4], cur_state[2]);
	and _ECO_1369(w_eco1369, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1370(w_eco1370, txtimeout, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1371(w_eco1371, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1372(w_eco1372, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1373(w_eco1373, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1374(w_eco1374, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1375(w_eco1375, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1376(w_eco1376, !txtimeout, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1377(w_eco1377, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], !cur_state[7], cur_state[8], !cur_state[0], cur_state[2]);
	and _ECO_1378(w_eco1378, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[9], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1379(w_eco1379, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1380(w_eco1380, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1381(w_eco1381, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1382(w_eco1382, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1383(w_eco1383, txtimeout, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1384(w_eco1384, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[1]);
	and _ECO_1385(w_eco1385, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1386(w_eco1386, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1387(w_eco1387, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1388(w_eco1388, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1389(w_eco1389, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1390(w_eco1390, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_1391(w_eco1391, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1392(w_eco1392, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1393(w_eco1393, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1394(w_eco1394, lk_txfsmidle, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], !cur_state[2], r2t_waittxid);
	and _ECO_1395(w_eco1395, lk_txfsmidle, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[1], !r2t_waittxid);
	and _ECO_1396(w_eco1396, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1397(w_eco1397, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1398(w_eco1398, !txtimeout, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[2], !r2t_waittxid);
	and _ECO_1399(w_eco1399, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1400(w_eco1400, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[0], !cur_state[1], !cur_state[2], r2t_waittxid);
	and _ECO_1401(w_eco1401, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1402(w_eco1402, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[1]);
	and _ECO_1403(w_eco1403, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1404(w_eco1404, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1405(w_eco1405, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1406(w_eco1406, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[1], !r2t_waittxid);
	and _ECO_1407(w_eco1407, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1408(w_eco1408, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], cur_state[4], cur_state[2]);
	and _ECO_1409(w_eco1409, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1410(w_eco1410, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], r2t_waittxid);
	and _ECO_1411(w_eco1411, !r2t_rxempty, !cur_state[11], cur_state[12], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[2]);
	and _ECO_1412(w_eco1412, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1413(w_eco1413, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1414(w_eco1414, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], r2t_waittxid);
	and _ECO_1415(w_eco1415, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1416(w_eco1416, lk_txfsmidle, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1417(w_eco1417, !txtimeout, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1418(w_eco1418, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1419(w_eco1419, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1420(w_eco1420, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1421(w_eco1421, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1422(w_eco1422, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1423(w_eco1423, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1424(w_eco1424, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], cur_state[4], !cur_state[0], cur_state[2]);
	and _ECO_1425(w_eco1425, !lk_txfsmidle, txtimeout, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1426(w_eco1426, lk_txfsmidle, !lk_txerror, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[9], cur_state[10], !cur_state[0], cur_state[2]);
	and _ECO_1427(w_eco1427, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1428(w_eco1428, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1429(w_eco1429, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1430(w_eco1430, lk_txfsmidle, !r2t_rxempty, lk_txerror, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[2], !r2t_waittxid);
	and _ECO_1431(w_eco1431, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[1], !cur_state[2]);
	and _ECO_1432(w_eco1432, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[10], !cur_state[3], cur_state[4], cur_state[2], !r2t_waittxid);
	and _ECO_1433(w_eco1433, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1434(w_eco1434, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1435(w_eco1435, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1436(w_eco1436, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1437(w_eco1437, !r2t_rxempty, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[1]);
	and _ECO_1438(w_eco1438, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[1]);
	and _ECO_1439(w_eco1439, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1440(w_eco1440, lk_txfsmidle, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1441(w_eco1441, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1442(w_eco1442, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1443(w_eco1443, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1444(w_eco1444, txtimeout, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1445(w_eco1445, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[14], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1446(w_eco1446, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1447(w_eco1447, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1448(w_eco1448, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1449(w_eco1449, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1]);
	and _ECO_1450(w_eco1450, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1451(w_eco1451, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1452(w_eco1452, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1453(w_eco1453, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1454(w_eco1454, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], cur_state[12], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1455(w_eco1455, !r2t_rxempty, !expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[2]);
	and _ECO_1456(w_eco1456, !r2t_rxempty, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[8], cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], cur_state[2]);
	and _ECO_1457(w_eco1457, !lk_txfsmidle, txtimeout, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1458(w_eco1458, lk_txfsmidle, !lk_txerror, !cur_state[11], !cur_state[12], cur_state[13], !cur_state[7], !cur_state[9], !cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1459(w_eco1459, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1460(w_eco1460, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], cur_state[10], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2]);
	and _ECO_1461(w_eco1461, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1462(w_eco1462, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1463(w_eco1463, !txtimeout, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1464(w_eco1464, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !r2t_waittxid);
	and _ECO_1465(w_eco1465, !txtimeout, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1466(w_eco1466, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1467(w_eco1467, lk_txfsmidle, !r2t_rxempty, lk_txerror, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1468(w_eco1468, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1469(w_eco1469, !lk_txfsmidle, !txtimeout, !r2t_rxempty, expire, !cur_state[11], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[8], !cur_state[9], !cur_state[3], !cur_state[5], !cur_state[6], !cur_state[0], cur_state[2], !r2t_waittxid);
	and _ECO_1470(w_eco1470, lk_txfsmidle, !r2t_rxempty, lk_txerror, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !cur_state[2]);
	and _ECO_1471(w_eco1471, !lk_txfsmidle, !txtimeout, !r2t_rxempty, !expire, !cur_state[11], !cur_state[12], !cur_state[13], !cur_state[14], !cur_state[7], !cur_state[10], !cur_state[0], cur_state[1], !cur_state[2]);
	or _ECO_1472(w_eco1472, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471);
	xor _ECO_out6(next_state[0], sub_wire6, w_eco1472);

endmodule