//
// Conformal-LEC: Version 11.10-d208 (10-Mar-2012) (64 bit executable)
//
module top(clk, rst, enb, out, reg_0, reg_1, fib, reg_0_p, reg_1_p, fib_p, State
    , State_p);
input  clk, rst, enb;
input   [16:0] reg_0_p;
input   [16:0] reg_1_p;
input   [16:0] fib_p;
input   [2:0] State_p;
output  [16:0] out;
output  [16:0] reg_0;
output  [16:0] reg_1;
output  [16:0] fib;
output  [2:0] State;
wire  \g318/inv_sel0 , \g318/w_0 , \g318/w_1 , \g312/inv_sel0 , \g312/w_0 , 
    \g312/w_1 , \g306/inv_sel0 , \g306/w_0 , \g306/w_1 , \g300/inv_sel0 , 
    \g300/w_0 , \g300/w_1 , \g294/inv_sel0 , \g294/w_0 , \g294/w_1 , 
    \g288/inv_sel0 , \g288/w_0 , \g288/w_1 , \g282/inv_sel0 , \g282/w_0 , 
    \g282/w_1 , \g276/inv_sel0 , \g276/w_0 , \g276/w_1 , \g270/inv_sel0 , 
    \g270/w_0 , \g270/w_1 , \g264/inv_sel0 , \g264/w_0 , \g264/w_1 , 
    \g258/inv_sel0 , \g258/w_0 , \g258/w_1 , \g252/inv_sel0 , \g252/w_0 , 
    \g252/w_1 , \g246/inv_sel0 , \g246/w_0 , \g246/w_1 , \g240/inv_sel0 , 
    \g240/w_0 , \g240/w_1 , \g234/inv_sel0 , \g234/w_0 , \g234/w_1 , 
    \g228/inv_sel0 , \g228/w_0 , \g228/w_1 , \g222/inv_sel0 , \g222/w_0 , 
    \g222/w_1 , \g216/inv_sel0 , \g216/w_0 , \g216/w_1 , \g215/inv_sel0 , 
    \g215/w_0 , \g215/w_1 , \g214/inv_sel0 , \g214/w_0 , \g214/w_1 , 
    \g209/inv_sel0 , \g209/w_0 , \g209/w_1 , \g208/inv_sel0 , \g208/w_0 , 
    \g208/w_1 , \g207/inv_sel0 , \g207/w_0 , \g207/w_1 , \g202/inv_sel0 , 
    \g202/w_0 , \g202/w_1 , \g201/inv_sel0 , \g201/w_0 , \g201/w_1 , 
    \g200/inv_sel0 , \g200/w_0 , \g200/w_1 , \g195/inv_sel0 , \g195/w_0 , 
    \g195/w_1 , \g194/inv_sel0 , \g194/w_0 , \g194/w_1 , \g193/inv_sel0 , 
    \g193/w_0 , \g193/w_1 , \g188/inv_sel0 , \g188/w_0 , \g188/w_1 , 
    \g187/inv_sel0 , \g187/w_0 , \g187/w_1 , \g186/inv_sel0 , \g186/w_0 , 
    \g186/w_1 , \g181/inv_sel0 , \g181/w_0 , \g181/w_1 , \g180/inv_sel0 , 
    \g180/w_0 , \g180/w_1 , \g179/inv_sel0 , \g179/w_0 , \g179/w_1 , 
    \g174/inv_sel0 , \g174/w_0 , \g174/w_1 , \g173/inv_sel0 , \g173/w_0 , 
    \g173/w_1 , \g172/inv_sel0 , \g172/w_0 , \g172/w_1 , \g167/inv_sel0 , 
    \g167/w_0 , \g167/w_1 , \g166/inv_sel0 , \g166/w_0 , \g166/w_1 , 
    \g165/inv_sel0 , \g165/w_0 , \g165/w_1 , \g160/inv_sel0 , \g160/w_0 , 
    \g160/w_1 , \g159/inv_sel0 , \g159/w_0 , \g159/w_1 , \g158/inv_sel0 , 
    \g158/w_0 , \g158/w_1 , \g153/inv_sel0 , \g153/w_0 , \g153/w_1 , 
    \g152/inv_sel0 , \g152/w_0 , \g152/w_1 , \g151/inv_sel0 , \g151/w_0 , 
    \g151/w_1 , \g146/inv_sel0 , \g146/w_0 , \g146/w_1 , \g145/inv_sel0 , 
    \g145/w_0 , \g145/w_1 , \g144/inv_sel0 , \g144/w_0 , \g144/w_1 , 
    \g139/inv_sel0 , \g139/w_0 , \g139/w_1 , \g138/inv_sel0 , \g138/w_0 , 
    \g138/w_1 , \g137/inv_sel0 , \g137/w_0 , \g137/w_1 , \g132/inv_sel0 , 
    \g132/w_0 , \g132/w_1 , \g131/inv_sel0 , \g131/w_0 , \g131/w_1 , 
    \g130/inv_sel0 , \g130/w_0 , \g130/w_1 , \g125/inv_sel0 , \g125/w_0 , 
    \g125/w_1 , \g124/inv_sel0 , \g124/w_0 , \g124/w_1 , \g123/inv_sel0 , 
    \g123/w_0 , \g123/w_1 , \g118/inv_sel0 , \g118/w_0 , \g118/w_1 , 
    \g117/inv_sel0 , \g117/w_0 , \g117/w_1 , \g116/inv_sel0 , \g116/w_0 , 
    \g116/w_1 , \g111/inv_sel0 , \g111/w_0 , \g111/w_1 , \g110/inv_sel0 , 
    \g110/w_0 , \g110/w_1 , \g109/inv_sel0 , \g109/w_0 , \g109/w_1 , 
    \g104/inv_sel0 , \g104/w_0 , \g104/w_1 , \g103/inv_sel0 , \g103/w_0 , 
    \g103/w_1 , \g102/inv_sel0 , \g102/w_0 , \g102/w_1 , \g97/inv_sel0 , 
    \g97/w_0 , \g97/w_1 , \g91/inv_sel0 , \g91/w_0 , \g91/w_1 , \g85/inv_sel0 , 
    \g85/w_0 , \g85/w_1 , \g79/inv_sel0 , \g79/w_0 , \g79/w_1 , \g73/inv_sel0 , 
    \g73/w_0 , \g73/w_1 , \g67/inv_sel0 , \g67/w_0 , \g67/w_1 , \g61/inv_sel0 , 
    \g61/w_0 , \g61/w_1 , \g55/inv_sel0 , \g55/w_0 , \g55/w_1 , \g49/inv_sel0 , 
    \g49/w_0 , \g49/w_1 , \g43/inv_sel0 , \g43/w_0 , \g43/w_1 , \g37/inv_sel0 , 
    \g37/w_0 , \g37/w_1 , \g31/inv_sel0 , \g31/w_0 , \g31/w_1 , \g25/inv_sel0 , 
    \g25/w_0 , \g25/w_1 , \g1008/inv_sel0 , \g1008/w_0 , \g1008/w_1 , 
    \g13/inv_sel0 , \g13/w_0 , \g13/w_1 , \g9/inv_sel0 , \g9/w_0 , \g9/w_1 , 
    \g3/inv_sel0 , \g3/w_0 , \g3/w_1 , n_1708, n_1707, n_1706, n_1705, n_1704, 
    n_1703, n_1702, n_1701, n_1700, n_1699, n_1698, n_1697, n_1422, n_1421, 
    n_1420, n_1419, n_1418, n_1417, n_1416, n_1415, n_1414, n_1413, n_1412, 
    n_1411, n_1410, n_1409, n_1408, n_1407, n_1406, n_1405, n_1404, n_1403, 
    n_1402, n_1401, n_1400, n_1399, n_1398, n_1397, n_1396, n_1395, n_1394, 
    n_1393, n_1392, n_1391, n_1390, n_1389, n_1388, n_1387, n_1220, n_1219, 
    n_1218, n_1217, n_1216, n_1215, n_1214, n_1213, n_1212, n_1211, n_1210, 
    n_1209, n_1208, n_1207, n_1206, n_1205, n_1203, n_1202, n_1201, n_1200, 
    n_1199, n_1198, n_1197, n_1196, n_1195, n_1194, n_1193, n_1192, n_1191, 
    n_1190, n_1189, n_1188, n_1187, n_1186, n_1185, n_1184, n_1183, n_1182, 
    n_1181, n_1180, n_1179, n_1178, n_1177, n_1176, n_1175, n_1174, n_1173, 
    n_1172, n_1171, n_1170, n_1169, n_1168, n_1167, n_1166, n_1165, n_1164, 
    n_1163, n_1162, n_1161, n_1160, n_1159, n_1158, n_1157, n_1156, n_1155, 
    n_1154, n_1153, n_1152, n_1151, n_1150, n_1149, n_1148, n_1147, n_1146, 
    n_1145, n_1144, n_1143, n_1142, n_1141, n_1140, n_1139, n_1138, n_1137, 
    n_1136, n_1135, n_1134, n_1133, n_1132, n_1131, n_1130, n_1129, n_1128, 
    n_1127, n_1126, n_1125, n_1124, n_1123, n_1122, n_1121, n_1120, n_1119, 
    n_1116, n_1115, n_881, n_598, n_595, n_594, n_395, n_393, n_392, n_391, 
    n_390, n_387, n_386, n_385, n_384, n_381, n_380, n_379, n_378, n_375, 
    n_374, n_373, n_372, n_369, n_368, n_367, n_366, n_363, n_362, n_361, 
    n_360, n_357, n_356, n_355, n_354, n_351, n_350, n_349, n_348, n_345, 
    n_344, n_343, n_342, n_339, n_338, n_337, n_336, n_333, n_332, n_331, 
    n_330, n_327, n_326, n_325, n_324, n_321, n_320, n_319, n_318, n_315, 
    n_314, n_313, n_312, n_309, n_308, n_307, n_306, n_303, n_302, n_301, 
    n_300, n_297, n_296, n_295, n_294, n_291, n_290, n_289, n_288, n_287, 
    n_286, n_282, n_281, n_280, n_279, n_278, n_277, n_273, n_272, n_271, 
    n_270, n_269, n_268, n_264, n_263, n_262, n_261, n_260, n_259, n_255, 
    n_254, n_253, n_252, n_251, n_250, n_246, n_245, n_244, n_243, n_242, 
    n_241, n_237, n_236, n_235, n_234, n_233, n_232, n_228, n_227, n_226, 
    n_208, n_207, n_206, n_205, n_201, n_200, n_199, n_198, n_197, n_196, 
    n_192, n_191, n_190, n_189, n_188, n_187, n_183, n_182, n_181, n_180, 
    n_179, n_178, n_174, n_173, n_172, n_171, n_170, n_169, n_165, n_164, 
    n_163, n_162, n_161, n_160, n_156, n_155, n_154, n_153, n_152, n_151, 
    n_147, n_146, n_145, n_144, n_143, n_142, n_138, n_137, n_136, n_135, 
    n_130, n_129, n_128, n_127, n_122, n_121, n_120, n_119, n_114, n_113, 
    n_112, n_111, n_106, n_105, n_104, n_103, n_98, n_97, n_96, n_95, n_90, 
    n_89, n_88, n_87, n_81, n_77, n_73, n_69, n_65, n_61, n_57, n_53, n_49, 
    n_45, n_41, n_37, n_33, n_29, n_25, n_21, n_17, n_14, n_12, n_10, n_8, 
    add_107_31_n_225, add_107_31_n_222, add_107_31_n_220, add_107_31_n_217, 
    add_107_31_n_214, add_107_31_n_211, add_107_31_n_209, add_107_31_n_205, 
    add_107_31_n_202, add_107_31_n_200, add_107_31_n_196, add_107_31_n_191, 
    add_107_31_n_189, add_107_31_n_188, add_107_31_n_187, add_107_31_n_185, 
    add_107_31_n_184, add_107_31_n_182, add_107_31_n_181, add_107_31_n_178, 
    add_107_31_n_176, add_107_31_n_169, add_107_31_n_166, add_107_31_n_164, 
    add_107_31_n_162, add_107_31_n_160, add_107_31_n_158, add_107_31_n_154, 
    add_107_31_n_152, add_107_31_n_151, add_107_31_n_147, add_107_31_n_142, 
    add_107_31_n_139, add_107_31_n_134, add_107_31_n_132, add_107_31_n_130, 
    add_107_31_n_129, add_107_31_n_124, add_107_31_n_122, add_107_31_n_120, 
    add_107_31_n_119, add_107_31_n_114, add_107_31_n_112, add_107_31_n_110, 
    add_107_31_n_109, add_107_31_n_108, add_107_31_n_106, add_107_31_n_103, 
    add_107_31_n_102, add_107_31_n_100, add_107_31_n_99, add_107_31_n_98, 
    add_107_31_n_97, add_107_31_n_96, add_107_31_n_94, add_107_31_n_93, 
    add_107_31_n_92, add_107_31_n_91, add_107_31_n_90, add_107_31_n_88, 
    add_107_31_n_87, add_107_31_n_86, add_107_31_n_85, add_107_31_n_84, 
    add_107_31_n_82, add_107_31_n_81, add_107_31_n_80, add_107_31_n_79, 
    add_107_31_n_78, add_107_31_n_76, add_107_31_n_75, add_107_31_n_74, 
    add_107_31_n_73, add_107_31_n_72, add_107_31_n_70, add_107_31_n_69, 
    add_107_31_n_68, add_107_31_n_67, add_107_31_n_66, add_107_31_n_64, 
    add_107_31_n_63, add_107_31_n_62, add_107_31_n_61, add_107_31_n_59, 
    add_107_31_n_56, add_107_31_n_53, enb, rst, clk;
wire   [2:0] State;
wire   [16:0] fib;
wire   [16:0] reg_1;
wire   [16:0] reg_0;
wire   [16:0] out;
wire   [2:0] State_p;
wire   [16:0] fib_p;
wire   [16:0] reg_1_p;
wire   [16:0] reg_0_p;
  assign State[2] = 1'b0;
  or \g318/org (n_390, \g318/w_0 , \g318/w_1 );
  and \g318/a_1 (\g318/w_1 , n_1387, reg_0_p[9]);
  and \g318/a_0 (\g318/w_0 , \g318/inv_sel0 , reg_1_p[9]);
  not \g318/i_0 (\g318/inv_sel0 , n_1387);
  or \g312/org (n_384, \g312/w_0 , \g312/w_1 );
  and \g312/a_1 (\g312/w_1 , n_1387, reg_0_p[10]);
  and \g312/a_0 (\g312/w_0 , \g312/inv_sel0 , reg_1_p[10]);
  not \g312/i_0 (\g312/inv_sel0 , n_1387);
  or \g306/org (n_378, \g306/w_0 , \g306/w_1 );
  and \g306/a_1 (\g306/w_1 , n_1387, reg_0_p[11]);
  and \g306/a_0 (\g306/w_0 , \g306/inv_sel0 , reg_1_p[11]);
  not \g306/i_0 (\g306/inv_sel0 , n_1387);
  or \g300/org (n_372, \g300/w_0 , \g300/w_1 );
  and \g300/a_1 (\g300/w_1 , n_1387, reg_0_p[12]);
  and \g300/a_0 (\g300/w_0 , \g300/inv_sel0 , reg_1_p[12]);
  not \g300/i_0 (\g300/inv_sel0 , n_1387);
  or \g294/org (n_366, \g294/w_0 , \g294/w_1 );
  and \g294/a_1 (\g294/w_1 , n_1387, reg_0_p[13]);
  and \g294/a_0 (\g294/w_0 , \g294/inv_sel0 , reg_1_p[13]);
  not \g294/i_0 (\g294/inv_sel0 , n_1387);
  or \g288/org (n_360, \g288/w_0 , \g288/w_1 );
  and \g288/a_1 (\g288/w_1 , n_1387, reg_0_p[14]);
  and \g288/a_0 (\g288/w_0 , \g288/inv_sel0 , reg_1_p[14]);
  not \g288/i_0 (\g288/inv_sel0 , n_1387);
  or \g282/org (n_354, \g282/w_0 , \g282/w_1 );
  and \g282/a_1 (\g282/w_1 , n_1387, reg_0_p[15]);
  and \g282/a_0 (\g282/w_0 , \g282/inv_sel0 , reg_1_p[15]);
  not \g282/i_0 (\g282/inv_sel0 , n_1387);
  or \g276/org (n_348, \g276/w_0 , \g276/w_1 );
  and \g276/a_1 (\g276/w_1 , n_1387, reg_0_p[16]);
  and \g276/a_0 (\g276/w_0 , \g276/inv_sel0 , reg_1_p[16]);
  not \g276/i_0 (\g276/inv_sel0 , n_1387);
  or \g270/org (n_342, \g270/w_0 , \g270/w_1 );
  and \g270/a_1 (\g270/w_1 , n_1387, reg_0_p[8]);
  and \g270/a_0 (\g270/w_0 , \g270/inv_sel0 , reg_1_p[8]);
  not \g270/i_0 (\g270/inv_sel0 , n_1387);
  or \g264/org (n_336, \g264/w_0 , \g264/w_1 );
  and \g264/a_1 (\g264/w_1 , n_1387, reg_0_p[5]);
  and \g264/a_0 (\g264/w_0 , \g264/inv_sel0 , reg_1_p[5]);
  not \g264/i_0 (\g264/inv_sel0 , n_1387);
  or \g258/org (n_330, \g258/w_0 , \g258/w_1 );
  and \g258/a_1 (\g258/w_1 , n_1387, reg_0_p[6]);
  and \g258/a_0 (\g258/w_0 , \g258/inv_sel0 , reg_1_p[6]);
  not \g258/i_0 (\g258/inv_sel0 , n_1387);
  or \g252/org (n_324, \g252/w_0 , \g252/w_1 );
  and \g252/a_1 (\g252/w_1 , n_1387, reg_0_p[7]);
  and \g252/a_0 (\g252/w_0 , \g252/inv_sel0 , reg_1_p[7]);
  not \g252/i_0 (\g252/inv_sel0 , n_1387);
  or \g246/org (n_318, \g246/w_0 , \g246/w_1 );
  and \g246/a_1 (\g246/w_1 , n_1387, reg_0_p[3]);
  and \g246/a_0 (\g246/w_0 , \g246/inv_sel0 , reg_1_p[3]);
  not \g246/i_0 (\g246/inv_sel0 , n_1387);
  or \g240/org (n_312, \g240/w_0 , \g240/w_1 );
  and \g240/a_1 (\g240/w_1 , n_1387, reg_0_p[4]);
  and \g240/a_0 (\g240/w_0 , \g240/inv_sel0 , reg_1_p[4]);
  not \g240/i_0 (\g240/inv_sel0 , n_1387);
  or \g234/org (n_306, \g234/w_0 , \g234/w_1 );
  and \g234/a_1 (\g234/w_1 , n_1387, reg_0_p[0]);
  and \g234/a_0 (\g234/w_0 , \g234/inv_sel0 , reg_1_p[0]);
  not \g234/i_0 (\g234/inv_sel0 , n_1387);
  or \g228/org (n_300, \g228/w_0 , \g228/w_1 );
  and \g228/a_1 (\g228/w_1 , n_1387, reg_0_p[1]);
  and \g228/a_0 (\g228/w_0 , \g228/inv_sel0 , reg_1_p[1]);
  not \g228/i_0 (\g228/inv_sel0 , n_1387);
  or \g222/org (n_294, \g222/w_0 , \g222/w_1 );
  and \g222/a_1 (\g222/w_1 , n_1387, reg_0_p[2]);
  and \g222/a_0 (\g222/w_0 , \g222/inv_sel0 , reg_1_p[2]);
  not \g222/i_0 (\g222/inv_sel0 , n_1387);
  or \g216/org (n_288, \g216/w_0 , \g216/w_1 );
  and \g216/a_1 (\g216/w_1 , State_p[0], n_286);
  and \g216/a_0 (\g216/w_0 , \g216/inv_sel0 , n_287);
  not \g216/i_0 (\g216/inv_sel0 , State_p[0]);
  or \g215/org (n_286, \g215/w_0 , \g215/w_1 );
  and \g215/a_1 (\g215/w_1 , State_p[1], fib_p[9]);
  and \g215/a_0 (\g215/w_0 , \g215/inv_sel0 , reg_1_p[9]);
  not \g215/i_0 (\g215/inv_sel0 , State_p[1]);
  or \g214/org (n_287, \g214/w_0 , \g214/w_1 );
  and \g214/a_1 (\g214/w_1 , State_p[1], n_53);
  and \g214/a_0 (\g214/w_0 , \g214/inv_sel0 , reg_0_p[9]);
  not \g214/i_0 (\g214/inv_sel0 , State_p[1]);
  or \g209/org (n_279, \g209/w_0 , \g209/w_1 );
  and \g209/a_1 (\g209/w_1 , State_p[0], n_277);
  and \g209/a_0 (\g209/w_0 , \g209/inv_sel0 , n_278);
  not \g209/i_0 (\g209/inv_sel0 , State_p[0]);
  or \g208/org (n_277, \g208/w_0 , \g208/w_1 );
  and \g208/a_1 (\g208/w_1 , State_p[1], fib_p[10]);
  and \g208/a_0 (\g208/w_0 , \g208/inv_sel0 , reg_1_p[10]);
  not \g208/i_0 (\g208/inv_sel0 , State_p[1]);
  or \g207/org (n_278, \g207/w_0 , \g207/w_1 );
  and \g207/a_1 (\g207/w_1 , State_p[1], n_57);
  and \g207/a_0 (\g207/w_0 , \g207/inv_sel0 , reg_0_p[10]);
  not \g207/i_0 (\g207/inv_sel0 , State_p[1]);
  or \g202/org (n_270, \g202/w_0 , \g202/w_1 );
  and \g202/a_1 (\g202/w_1 , State_p[0], n_268);
  and \g202/a_0 (\g202/w_0 , \g202/inv_sel0 , n_269);
  not \g202/i_0 (\g202/inv_sel0 , State_p[0]);
  or \g201/org (n_268, \g201/w_0 , \g201/w_1 );
  and \g201/a_1 (\g201/w_1 , State_p[1], fib_p[11]);
  and \g201/a_0 (\g201/w_0 , \g201/inv_sel0 , reg_1_p[11]);
  not \g201/i_0 (\g201/inv_sel0 , State_p[1]);
  or \g200/org (n_269, \g200/w_0 , \g200/w_1 );
  and \g200/a_1 (\g200/w_1 , State_p[1], n_61);
  and \g200/a_0 (\g200/w_0 , \g200/inv_sel0 , reg_0_p[11]);
  not \g200/i_0 (\g200/inv_sel0 , State_p[1]);
  or \g195/org (n_261, \g195/w_0 , \g195/w_1 );
  and \g195/a_1 (\g195/w_1 , State_p[0], n_259);
  and \g195/a_0 (\g195/w_0 , \g195/inv_sel0 , n_260);
  not \g195/i_0 (\g195/inv_sel0 , State_p[0]);
  or \g194/org (n_259, \g194/w_0 , \g194/w_1 );
  and \g194/a_1 (\g194/w_1 , State_p[1], fib_p[12]);
  and \g194/a_0 (\g194/w_0 , \g194/inv_sel0 , reg_1_p[12]);
  not \g194/i_0 (\g194/inv_sel0 , State_p[1]);
  or \g193/org (n_260, \g193/w_0 , \g193/w_1 );
  and \g193/a_1 (\g193/w_1 , State_p[1], n_65);
  and \g193/a_0 (\g193/w_0 , \g193/inv_sel0 , reg_0_p[12]);
  not \g193/i_0 (\g193/inv_sel0 , State_p[1]);
  or \g188/org (n_252, \g188/w_0 , \g188/w_1 );
  and \g188/a_1 (\g188/w_1 , State_p[0], n_250);
  and \g188/a_0 (\g188/w_0 , \g188/inv_sel0 , n_251);
  not \g188/i_0 (\g188/inv_sel0 , State_p[0]);
  or \g187/org (n_250, \g187/w_0 , \g187/w_1 );
  and \g187/a_1 (\g187/w_1 , State_p[1], fib_p[13]);
  and \g187/a_0 (\g187/w_0 , \g187/inv_sel0 , reg_1_p[13]);
  not \g187/i_0 (\g187/inv_sel0 , State_p[1]);
  or \g186/org (n_251, \g186/w_0 , \g186/w_1 );
  and \g186/a_1 (\g186/w_1 , State_p[1], n_69);
  and \g186/a_0 (\g186/w_0 , \g186/inv_sel0 , reg_0_p[13]);
  not \g186/i_0 (\g186/inv_sel0 , State_p[1]);
  or \g181/org (n_243, \g181/w_0 , \g181/w_1 );
  and \g181/a_1 (\g181/w_1 , State_p[0], n_241);
  and \g181/a_0 (\g181/w_0 , \g181/inv_sel0 , n_242);
  not \g181/i_0 (\g181/inv_sel0 , State_p[0]);
  or \g180/org (n_241, \g180/w_0 , \g180/w_1 );
  and \g180/a_1 (\g180/w_1 , State_p[1], fib_p[14]);
  and \g180/a_0 (\g180/w_0 , \g180/inv_sel0 , reg_1_p[14]);
  not \g180/i_0 (\g180/inv_sel0 , State_p[1]);
  or \g179/org (n_242, \g179/w_0 , \g179/w_1 );
  and \g179/a_1 (\g179/w_1 , State_p[1], n_73);
  and \g179/a_0 (\g179/w_0 , \g179/inv_sel0 , reg_0_p[14]);
  not \g179/i_0 (\g179/inv_sel0 , State_p[1]);
  or \g174/org (n_234, \g174/w_0 , \g174/w_1 );
  and \g174/a_1 (\g174/w_1 , State_p[0], n_232);
  and \g174/a_0 (\g174/w_0 , \g174/inv_sel0 , n_233);
  not \g174/i_0 (\g174/inv_sel0 , State_p[0]);
  or \g173/org (n_232, \g173/w_0 , \g173/w_1 );
  and \g173/a_1 (\g173/w_1 , State_p[1], fib_p[15]);
  and \g173/a_0 (\g173/w_0 , \g173/inv_sel0 , reg_1_p[15]);
  not \g173/i_0 (\g173/inv_sel0 , State_p[1]);
  or \g172/org (n_233, \g172/w_0 , \g172/w_1 );
  and \g172/a_1 (\g172/w_1 , State_p[1], n_77);
  and \g172/a_0 (\g172/w_0 , \g172/inv_sel0 , reg_0_p[15]);
  not \g172/i_0 (\g172/inv_sel0 , State_p[1]);
  or \g167/org (n_1708, \g167/w_0 , \g167/w_1 );
  and \g167/a_1 (\g167/w_1 , State_p[0], n_1706);
  and \g167/a_0 (\g167/w_0 , \g167/inv_sel0 , n_1707);
  not \g167/i_0 (\g167/inv_sel0 , State_p[0]);
  or \g166/org (n_1706, \g166/w_0 , \g166/w_1 );
  and \g166/a_1 (\g166/w_1 , State_p[1], fib_p[16]);
  and \g166/a_0 (\g166/w_0 , \g166/inv_sel0 , reg_1_p[16]);
  not \g166/i_0 (\g166/inv_sel0 , State_p[1]);
  or \g165/org (n_1707, \g165/w_0 , \g165/w_1 );
  and \g165/a_1 (\g165/w_1 , State_p[1], n_81);
  and \g165/a_0 (\g165/w_0 , \g165/inv_sel0 , reg_0_p[16]);
  not \g165/i_0 (\g165/inv_sel0 , State_p[1]);
  or \g160/org (n_1702, \g160/w_0 , \g160/w_1 );
  and \g160/a_1 (\g160/w_1 , State_p[0], n_1700);
  and \g160/a_0 (\g160/w_0 , \g160/inv_sel0 , n_1701);
  not \g160/i_0 (\g160/inv_sel0 , State_p[0]);
  or \g159/org (n_1700, \g159/w_0 , \g159/w_1 );
  and \g159/a_1 (\g159/w_1 , State_p[1], fib_p[8]);
  and \g159/a_0 (\g159/w_0 , \g159/inv_sel0 , reg_1_p[8]);
  not \g159/i_0 (\g159/inv_sel0 , State_p[1]);
  or \g158/org (n_1701, \g158/w_0 , \g158/w_1 );
  and \g158/a_1 (\g158/w_1 , State_p[1], n_49);
  and \g158/a_0 (\g158/w_0 , \g158/inv_sel0 , reg_0_p[8]);
  not \g158/i_0 (\g158/inv_sel0 , State_p[1]);
  or \g153/org (n_207, \g153/w_0 , \g153/w_1 );
  and \g153/a_1 (\g153/w_1 , State_p[0], n_205);
  and \g153/a_0 (\g153/w_0 , \g153/inv_sel0 , n_206);
  not \g153/i_0 (\g153/inv_sel0 , State_p[0]);
  or \g152/org (n_205, \g152/w_0 , \g152/w_1 );
  and \g152/a_1 (\g152/w_1 , State_p[1], fib_p[5]);
  and \g152/a_0 (\g152/w_0 , \g152/inv_sel0 , reg_1_p[5]);
  not \g152/i_0 (\g152/inv_sel0 , State_p[1]);
  or \g151/org (n_206, \g151/w_0 , \g151/w_1 );
  and \g151/a_1 (\g151/w_1 , State_p[1], n_37);
  and \g151/a_0 (\g151/w_0 , \g151/inv_sel0 , reg_0_p[5]);
  not \g151/i_0 (\g151/inv_sel0 , State_p[1]);
  or \g146/org (n_198, \g146/w_0 , \g146/w_1 );
  and \g146/a_1 (\g146/w_1 , State_p[0], n_196);
  and \g146/a_0 (\g146/w_0 , \g146/inv_sel0 , n_197);
  not \g146/i_0 (\g146/inv_sel0 , State_p[0]);
  or \g145/org (n_196, \g145/w_0 , \g145/w_1 );
  and \g145/a_1 (\g145/w_1 , State_p[1], fib_p[6]);
  and \g145/a_0 (\g145/w_0 , \g145/inv_sel0 , reg_1_p[6]);
  not \g145/i_0 (\g145/inv_sel0 , State_p[1]);
  or \g144/org (n_197, \g144/w_0 , \g144/w_1 );
  and \g144/a_1 (\g144/w_1 , State_p[1], n_41);
  and \g144/a_0 (\g144/w_0 , \g144/inv_sel0 , reg_0_p[6]);
  not \g144/i_0 (\g144/inv_sel0 , State_p[1]);
  or \g139/org (n_189, \g139/w_0 , \g139/w_1 );
  and \g139/a_1 (\g139/w_1 , State_p[0], n_187);
  and \g139/a_0 (\g139/w_0 , \g139/inv_sel0 , n_188);
  not \g139/i_0 (\g139/inv_sel0 , State_p[0]);
  or \g138/org (n_187, \g138/w_0 , \g138/w_1 );
  and \g138/a_1 (\g138/w_1 , State_p[1], fib_p[7]);
  and \g138/a_0 (\g138/w_0 , \g138/inv_sel0 , reg_1_p[7]);
  not \g138/i_0 (\g138/inv_sel0 , State_p[1]);
  or \g137/org (n_188, \g137/w_0 , \g137/w_1 );
  and \g137/a_1 (\g137/w_1 , State_p[1], n_45);
  and \g137/a_0 (\g137/w_0 , \g137/inv_sel0 , reg_0_p[7]);
  not \g137/i_0 (\g137/inv_sel0 , State_p[1]);
  or \g132/org (n_180, \g132/w_0 , \g132/w_1 );
  and \g132/a_1 (\g132/w_1 , State_p[0], n_178);
  and \g132/a_0 (\g132/w_0 , \g132/inv_sel0 , n_179);
  not \g132/i_0 (\g132/inv_sel0 , State_p[0]);
  or \g131/org (n_178, \g131/w_0 , \g131/w_1 );
  and \g131/a_1 (\g131/w_1 , State_p[1], fib_p[3]);
  and \g131/a_0 (\g131/w_0 , \g131/inv_sel0 , reg_1_p[3]);
  not \g131/i_0 (\g131/inv_sel0 , State_p[1]);
  or \g130/org (n_179, \g130/w_0 , \g130/w_1 );
  and \g130/a_1 (\g130/w_1 , State_p[1], n_29);
  and \g130/a_0 (\g130/w_0 , \g130/inv_sel0 , reg_0_p[3]);
  not \g130/i_0 (\g130/inv_sel0 , State_p[1]);
  or \g125/org (n_171, \g125/w_0 , \g125/w_1 );
  and \g125/a_1 (\g125/w_1 , State_p[0], n_169);
  and \g125/a_0 (\g125/w_0 , \g125/inv_sel0 , n_170);
  not \g125/i_0 (\g125/inv_sel0 , State_p[0]);
  or \g124/org (n_169, \g124/w_0 , \g124/w_1 );
  and \g124/a_1 (\g124/w_1 , State_p[1], fib_p[4]);
  and \g124/a_0 (\g124/w_0 , \g124/inv_sel0 , reg_1_p[4]);
  not \g124/i_0 (\g124/inv_sel0 , State_p[1]);
  or \g123/org (n_170, \g123/w_0 , \g123/w_1 );
  and \g123/a_1 (\g123/w_1 , State_p[1], n_33);
  and \g123/a_0 (\g123/w_0 , \g123/inv_sel0 , reg_0_p[4]);
  not \g123/i_0 (\g123/inv_sel0 , State_p[1]);
  or \g118/org (n_162, \g118/w_0 , \g118/w_1 );
  and \g118/a_1 (\g118/w_1 , State_p[0], n_160);
  and \g118/a_0 (\g118/w_0 , \g118/inv_sel0 , n_161);
  not \g118/i_0 (\g118/inv_sel0 , State_p[0]);
  or \g117/org (n_160, \g117/w_0 , \g117/w_1 );
  and \g117/a_1 (\g117/w_1 , State_p[1], fib_p[0]);
  and \g117/a_0 (\g117/w_0 , \g117/inv_sel0 , reg_1_p[0]);
  not \g117/i_0 (\g117/inv_sel0 , State_p[1]);
  or \g116/org (n_161, \g116/w_0 , \g116/w_1 );
  and \g116/a_1 (\g116/w_1 , State_p[1], n_17);
  and \g116/a_0 (\g116/w_0 , \g116/inv_sel0 , reg_0_p[0]);
  not \g116/i_0 (\g116/inv_sel0 , State_p[1]);
  or \g111/org (n_153, \g111/w_0 , \g111/w_1 );
  and \g111/a_1 (\g111/w_1 , State_p[0], n_151);
  and \g111/a_0 (\g111/w_0 , \g111/inv_sel0 , n_152);
  not \g111/i_0 (\g111/inv_sel0 , State_p[0]);
  or \g110/org (n_151, \g110/w_0 , \g110/w_1 );
  and \g110/a_1 (\g110/w_1 , State_p[1], fib_p[1]);
  and \g110/a_0 (\g110/w_0 , \g110/inv_sel0 , reg_1_p[1]);
  not \g110/i_0 (\g110/inv_sel0 , State_p[1]);
  or \g109/org (n_152, \g109/w_0 , \g109/w_1 );
  and \g109/a_1 (\g109/w_1 , State_p[1], n_21);
  and \g109/a_0 (\g109/w_0 , \g109/inv_sel0 , reg_0_p[1]);
  not \g109/i_0 (\g109/inv_sel0 , State_p[1]);
  or \g104/org (n_144, \g104/w_0 , \g104/w_1 );
  and \g104/a_1 (\g104/w_1 , State_p[0], n_142);
  and \g104/a_0 (\g104/w_0 , \g104/inv_sel0 , n_143);
  not \g104/i_0 (\g104/inv_sel0 , State_p[0]);
  or \g103/org (n_142, \g103/w_0 , \g103/w_1 );
  and \g103/a_1 (\g103/w_1 , State_p[1], fib_p[2]);
  and \g103/a_0 (\g103/w_0 , \g103/inv_sel0 , reg_1_p[2]);
  not \g103/i_0 (\g103/inv_sel0 , State_p[1]);
  or \g102/org (n_143, \g102/w_0 , \g102/w_1 );
  and \g102/a_1 (\g102/w_1 , State_p[1], n_25);
  and \g102/a_0 (\g102/w_0 , \g102/inv_sel0 , reg_0_p[2]);
  not \g102/i_0 (\g102/inv_sel0 , State_p[1]);
  or \g97/org (n_135, \g97/w_0 , \g97/w_1 );
  and \g97/a_1 (\g97/w_1 , n_1387, reg_1_p[9]);
  and \g97/a_0 (\g97/w_0 , \g97/inv_sel0 , n_53);
  not \g97/i_0 (\g97/inv_sel0 , n_1387);
  or \g91/org (n_127, \g91/w_0 , \g91/w_1 );
  and \g91/a_1 (\g91/w_1 , n_1387, reg_1_p[10]);
  and \g91/a_0 (\g91/w_0 , \g91/inv_sel0 , n_57);
  not \g91/i_0 (\g91/inv_sel0 , n_1387);
  or \g85/org (n_119, \g85/w_0 , \g85/w_1 );
  and \g85/a_1 (\g85/w_1 , n_1387, reg_1_p[11]);
  and \g85/a_0 (\g85/w_0 , \g85/inv_sel0 , n_61);
  not \g85/i_0 (\g85/inv_sel0 , n_1387);
  or \g79/org (n_111, \g79/w_0 , \g79/w_1 );
  and \g79/a_1 (\g79/w_1 , n_1387, reg_1_p[12]);
  and \g79/a_0 (\g79/w_0 , \g79/inv_sel0 , n_65);
  not \g79/i_0 (\g79/inv_sel0 , n_1387);
  or \g73/org (n_103, \g73/w_0 , \g73/w_1 );
  and \g73/a_1 (\g73/w_1 , n_1387, reg_1_p[13]);
  and \g73/a_0 (\g73/w_0 , \g73/inv_sel0 , n_69);
  not \g73/i_0 (\g73/inv_sel0 , n_1387);
  or \g67/org (n_95, \g67/w_0 , \g67/w_1 );
  and \g67/a_1 (\g67/w_1 , n_1387, reg_1_p[14]);
  and \g67/a_0 (\g67/w_0 , \g67/inv_sel0 , n_73);
  not \g67/i_0 (\g67/inv_sel0 , n_1387);
  or \g61/org (n_87, \g61/w_0 , \g61/w_1 );
  and \g61/a_1 (\g61/w_1 , n_1387, reg_1_p[15]);
  and \g61/a_0 (\g61/w_0 , \g61/inv_sel0 , n_77);
  not \g61/i_0 (\g61/inv_sel0 , n_1387);
  or \g55/org (n_1419, \g55/w_0 , \g55/w_1 );
  and \g55/a_1 (\g55/w_1 , n_1387, reg_1_p[16]);
  and \g55/a_0 (\g55/w_0 , \g55/inv_sel0 , n_81);
  not \g55/i_0 (\g55/inv_sel0 , n_1387);
  or \g49/org (n_1415, \g49/w_0 , \g49/w_1 );
  and \g49/a_1 (\g49/w_1 , n_1387, reg_1_p[8]);
  and \g49/a_0 (\g49/w_0 , \g49/inv_sel0 , n_49);
  not \g49/i_0 (\g49/inv_sel0 , n_1387);
  or \g43/org (n_1411, \g43/w_0 , \g43/w_1 );
  and \g43/a_1 (\g43/w_1 , n_1387, reg_1_p[5]);
  and \g43/a_0 (\g43/w_0 , \g43/inv_sel0 , n_37);
  not \g43/i_0 (\g43/inv_sel0 , n_1387);
  or \g37/org (n_1407, \g37/w_0 , \g37/w_1 );
  and \g37/a_1 (\g37/w_1 , n_1387, reg_1_p[6]);
  and \g37/a_0 (\g37/w_0 , \g37/inv_sel0 , n_41);
  not \g37/i_0 (\g37/inv_sel0 , n_1387);
  or \g31/org (n_1403, \g31/w_0 , \g31/w_1 );
  and \g31/a_1 (\g31/w_1 , n_1387, reg_1_p[7]);
  and \g31/a_0 (\g31/w_0 , \g31/inv_sel0 , n_45);
  not \g31/i_0 (\g31/inv_sel0 , n_1387);
  or \g25/org (n_1399, \g25/w_0 , \g25/w_1 );
  and \g25/a_1 (\g25/w_1 , n_1387, reg_1_p[3]);
  and \g25/a_0 (\g25/w_0 , \g25/inv_sel0 , n_29);
  not \g25/i_0 (\g25/inv_sel0 , n_1387);
  or \g1008/org (n_1395, \g1008/w_0 , \g1008/w_1 );
  and \g1008/a_1 (\g1008/w_1 , n_1387, reg_1_p[4]);
  and \g1008/a_0 (\g1008/w_0 , \g1008/inv_sel0 , n_33);
  not \g1008/i_0 (\g1008/inv_sel0 , n_1387);
  or \g13/org (n_1391, \g13/w_0 , \g13/w_1 );
  and \g13/a_1 (\g13/w_1 , n_1387, reg_1_p[2]);
  and \g13/a_0 (\g13/w_0 , \g13/inv_sel0 , n_25);
  not \g13/i_0 (\g13/inv_sel0 , n_1387);
  or \g9/org (n_1389, \g9/w_0 , \g9/w_1 );
  and \g9/a_1 (\g9/w_1 , n_1387, reg_1_p[0]);
  and \g9/a_0 (\g9/w_0 , \g9/inv_sel0 , n_17);
  not \g9/i_0 (\g9/inv_sel0 , n_1387);
  or \g3/org (n_1388, \g3/w_0 , \g3/w_1 );
  and \g3/a_1 (\g3/w_1 , n_1387, reg_1_p[1]);
  and \g3/a_0 (\g3/w_0 , \g3/inv_sel0 , n_21);
  not \g3/i_0 (\g3/inv_sel0 , n_1387);
  assign fib[16] = out[16];
  assign fib[15] = out[15];
  assign fib[14] = out[14];
  assign fib[13] = out[13];
  assign fib[12] = out[12];
  assign fib[11] = out[11];
  assign fib[10] = out[10];
  assign fib[9] = out[9];
  assign fib[8] = out[8];
  assign fib[7] = out[7];
  assign fib[6] = out[6];
  assign fib[5] = out[5];
  assign fib[4] = out[4];
  assign fib[3] = out[3];
  assign fib[2] = out[2];
  assign fib[1] = out[1];
  assign fib[0] = out[0];
  xor add_107_31_g1(n_17, reg_0_p[0], reg_1_p[0]);
  nor add_107_31_g10(add_107_31_n_62, reg_0_p[3], reg_1_p[3]);
  nand add_107_31_g103(add_107_31_n_162, add_107_31_n_132, add_107_31_n_134);
  nand add_107_31_g106(add_107_31_n_200, add_107_31_n_67, n_1134);
  nand add_107_31_g107(add_107_31_n_142, add_107_31_n_112, add_107_31_n_139);
  nand add_107_31_g108(add_107_31_n_202, add_107_31_n_109, add_107_31_n_142);
  nand add_107_31_g11(add_107_31_n_63, reg_0_p[3], reg_1_p[3]);
  nand add_107_31_g111(add_107_31_n_205, n_1139, n_1142);
  nand add_107_31_g114(add_107_31_n_166, n_1149, n_1151);
  nor add_107_31_g115(add_107_31_n_152, add_107_31_n_96, add_107_31_n_151);
  nor add_107_31_g118(add_107_31_n_176, add_107_31_n_96, add_107_31_n_154);
  nor add_107_31_g12(add_107_31_n_72, reg_0_p[4], reg_1_p[4]);
  nor add_107_31_g124(add_107_31_n_160, add_107_31_n_158, add_107_31_n_151);
  nor add_107_31_g127(add_107_31_n_182, add_107_31_n_154, add_107_31_n_158);
  nor add_107_31_g128(add_107_31_n_164, add_107_31_n_162, add_107_31_n_151);
  nand add_107_31_g13(add_107_31_n_67, reg_0_p[4], reg_1_p[4]);
  nor add_107_31_g131(add_107_31_n_185, add_107_31_n_154, add_107_31_n_162);
  nand add_107_31_g134(add_107_31_n_209, add_107_31_n_79, n_1164);
  nand add_107_31_g135(add_107_31_n_169, add_107_31_n_122, add_107_31_n_166);
  nand add_107_31_g136(add_107_31_n_211, add_107_31_n_119, add_107_31_n_169);
  nand add_107_31_g139(add_107_31_n_214, n_1165, n_1168);
  nor add_107_31_g14(add_107_31_n_68, reg_0_p[5], reg_1_p[5]);
  nand add_107_31_g142(add_107_31_n_217, add_107_31_n_151, n_1169);
  nand add_107_31_g143(add_107_31_n_178, add_107_31_n_176, add_107_31_n_166);
  nand add_107_31_g144(add_107_31_n_220, n_1171, add_107_31_n_178);
  nand add_107_31_g145(add_107_31_n_181, n_1172, add_107_31_n_166);
  nand add_107_31_g146(add_107_31_n_222, n_1176, add_107_31_n_181);
  nand add_107_31_g147(add_107_31_n_184, add_107_31_n_182, add_107_31_n_166);
  nand add_107_31_g148(add_107_31_n_225, n_1180, add_107_31_n_184);
  nand add_107_31_g149(add_107_31_n_187, add_107_31_n_185, add_107_31_n_166);
  nand add_107_31_g15(add_107_31_n_69, reg_0_p[5], reg_1_p[5]);
  nand add_107_31_g150(add_107_31_n_189, n_1187, add_107_31_n_187);
  xnor add_107_31_g157(n_25, add_107_31_n_103, n_1205);
  nor add_107_31_g16(add_107_31_n_78, reg_0_p[6], reg_1_p[6]);
  xnor add_107_31_g160(n_29, add_107_31_n_196, n_1206);
  xnor add_107_31_g162(n_33, add_107_31_n_139, n_1207);
  xnor add_107_31_g165(n_37, add_107_31_n_200, n_1208);
  xnor add_107_31_g167(n_41, add_107_31_n_202, n_1209);
  nand add_107_31_g17(add_107_31_n_73, reg_0_p[6], reg_1_p[6]);
  xnor add_107_31_g170(n_45, add_107_31_n_205, n_1210);
  xnor add_107_31_g172(n_49, add_107_31_n_166, n_1211);
  xnor add_107_31_g175(n_53, add_107_31_n_209, n_1212);
  xnor add_107_31_g177(n_57, add_107_31_n_211, n_1213);
  nor add_107_31_g18(add_107_31_n_74, reg_0_p[7], reg_1_p[7]);
  xnor add_107_31_g180(n_61, add_107_31_n_214, n_1214);
  xnor add_107_31_g183(n_65, add_107_31_n_217, n_1215);
  xnor add_107_31_g186(n_69, add_107_31_n_220, n_1216);
  xnor add_107_31_g188(n_73, add_107_31_n_222, n_1217);
  nand add_107_31_g19(add_107_31_n_75, reg_0_p[7], reg_1_p[7]);
  xnor add_107_31_g191(n_77, add_107_31_n_225, n_1218);
  xnor add_107_31_g193(n_81, add_107_31_n_189, n_1219);
  nand add_107_31_g2(add_107_31_n_53, reg_0_p[0], reg_1_p[0]);
  nor add_107_31_g20(add_107_31_n_84, reg_0_p[8], reg_1_p[8]);
  nand add_107_31_g21(add_107_31_n_79, reg_0_p[8], reg_1_p[8]);
  nor add_107_31_g22(add_107_31_n_80, reg_0_p[9], reg_1_p[9]);
  nand add_107_31_g23(add_107_31_n_81, reg_0_p[9], reg_1_p[9]);
  nor add_107_31_g24(add_107_31_n_90, reg_0_p[10], reg_1_p[10]);
  nand add_107_31_g25(add_107_31_n_85, reg_0_p[10], reg_1_p[10]);
  nor add_107_31_g26(add_107_31_n_86, reg_0_p[11], reg_1_p[11]);
  nand add_107_31_g27(add_107_31_n_87, reg_0_p[11], reg_1_p[11]);
  nor add_107_31_g28(add_107_31_n_96, reg_0_p[12], reg_1_p[12]);
  nand add_107_31_g29(add_107_31_n_91, reg_0_p[12], reg_1_p[12]);
  nor add_107_31_g30(add_107_31_n_92, reg_0_p[13], reg_1_p[13]);
  nand add_107_31_g31(add_107_31_n_93, reg_0_p[13], reg_1_p[13]);
  nor add_107_31_g32(add_107_31_n_102, reg_0_p[14], reg_1_p[14]);
  nand add_107_31_g33(add_107_31_n_97, reg_0_p[14], reg_1_p[14]);
  nor add_107_31_g34(add_107_31_n_98, reg_0_p[15], reg_1_p[15]);
  nand add_107_31_g35(add_107_31_n_99, reg_0_p[15], reg_1_p[15]);
  nor add_107_31_g36(add_107_31_n_188, reg_0_p[16], reg_1_p[16]);
  nand add_107_31_g37(add_107_31_n_191, reg_0_p[16], reg_1_p[16]);
  nand add_107_31_g40(add_107_31_n_103, add_107_31_n_59, n_1133);
  nor add_107_31_g41(add_107_31_n_64, add_107_31_n_61, add_107_31_n_62);
  nor add_107_31_g44(add_107_31_n_106, add_107_31_n_66, add_107_31_n_62);
  nor add_107_31_g45(add_107_31_n_70, add_107_31_n_67, add_107_31_n_68);
  nor add_107_31_g48(add_107_31_n_112, add_107_31_n_72, add_107_31_n_68);
  nor add_107_31_g49(add_107_31_n_76, add_107_31_n_73, add_107_31_n_74);
  nor add_107_31_g52(add_107_31_n_114, add_107_31_n_78, add_107_31_n_74);
  nor add_107_31_g53(add_107_31_n_82, add_107_31_n_79, add_107_31_n_80);
  nor add_107_31_g56(add_107_31_n_122, add_107_31_n_84, add_107_31_n_80);
  nor add_107_31_g57(add_107_31_n_88, add_107_31_n_85, add_107_31_n_86);
  nor add_107_31_g6(add_107_31_n_56, reg_0_p[1], reg_1_p[1]);
  nor add_107_31_g60(add_107_31_n_124, add_107_31_n_90, add_107_31_n_86);
  nor add_107_31_g61(add_107_31_n_94, add_107_31_n_91, add_107_31_n_92);
  nor add_107_31_g64(add_107_31_n_132, add_107_31_n_96, add_107_31_n_92);
  nor add_107_31_g65(add_107_31_n_100, add_107_31_n_97, add_107_31_n_98);
  nor add_107_31_g68(add_107_31_n_134, add_107_31_n_102, add_107_31_n_98);
  nand add_107_31_g7(add_107_31_n_59, reg_0_p[1], reg_1_p[1]);
  nand add_107_31_g71(add_107_31_n_196, add_107_31_n_61, n_1189);
  nand add_107_31_g72(add_107_31_n_108, add_107_31_n_106, add_107_31_n_103);
  nand add_107_31_g73(add_107_31_n_139, n_1129, add_107_31_n_108);
  nor add_107_31_g74(add_107_31_n_110, add_107_31_n_78, add_107_31_n_109);
  nor add_107_31_g8(add_107_31_n_66, reg_0_p[2], reg_1_p[2]);
  nand add_107_31_g83(add_107_31_n_147, add_107_31_n_112, add_107_31_n_114);
  nor add_107_31_g84(add_107_31_n_120, add_107_31_n_90, add_107_31_n_119);
  nand add_107_31_g9(add_107_31_n_61, reg_0_p[2], reg_1_p[2]);
  nand add_107_31_g93(add_107_31_n_154, add_107_31_n_122, add_107_31_n_124);
  nor add_107_31_g94(add_107_31_n_130, add_107_31_n_102, add_107_31_n_129);
  not g7(reg_1[1], n_1697);
  not g19(State[1], n_595);
  not g29(State[0], n_598);
  xor g54(n_881, enb, State_p[0]);
  xor g681(n_21, add_107_31_n_53, n_1220);
  not g889(n_1115, State_p[1]);
  not g893(n_1119, n_881);
  not g894(n_1120, add_107_31_n_62);
  not g895(n_1121, add_107_31_n_96);
  not g896(n_1122, add_107_31_n_92);
  not g897(n_1123, add_107_31_n_132);
  not g898(n_1124, add_107_31_n_102);
  not g899(n_1125, add_107_31_n_98);
  not g900(n_1126, add_107_31_n_134);
  not g901(n_1127, add_107_31_n_72);
  not g902(n_1128, add_107_31_n_63);
  nor g903(n_1129, n_1128, add_107_31_n_64);
  not g904(n_1130, add_107_31_n_66);
  not g905(n_1131, add_107_31_n_53);
  not g906(n_1132, add_107_31_n_56);
  nand g907(n_1133, n_1131, n_1132);
  nand g908(n_1134, n_1127, add_107_31_n_139);
  not g909(n_1135, add_107_31_n_68);
  not g910(n_1136, add_107_31_n_69);
  nor g911(add_107_31_n_109, n_1136, add_107_31_n_70);
  not g912(n_1137, add_107_31_n_73);
  not g913(n_1138, add_107_31_n_78);
  nor g914(n_1139, n_1137, add_107_31_n_110);
  nand g915(n_1140, n_1138, add_107_31_n_112);
  not g916(n_1141, n_1140);
  nand g917(n_1142, add_107_31_n_139, n_1141);
  not g918(n_1143, add_107_31_n_75);
  not g919(n_1144, add_107_31_n_74);
  nor g920(n_1145, n_1143, add_107_31_n_76);
  not g921(n_1146, n_1145);
  not g922(n_1147, add_107_31_n_114);
  nor g923(n_1148, n_1147, add_107_31_n_109);
  nor g924(n_1149, n_1146, n_1148);
  not g925(n_1150, add_107_31_n_147);
  nand g926(n_1151, add_107_31_n_139, n_1150);
  not g927(n_1152, add_107_31_n_87);
  not g928(n_1153, add_107_31_n_85);
  not g929(n_1154, add_107_31_n_86);
  nor g930(n_1155, n_1152, add_107_31_n_88);
  not g931(n_1156, n_1155);
  not g932(n_1157, add_107_31_n_90);
  not g933(n_1158, add_107_31_n_124);
  not g934(n_1159, add_107_31_n_81);
  not g935(n_1160, add_107_31_n_80);
  nor g936(add_107_31_n_119, n_1159, add_107_31_n_82);
  nor g937(n_1161, n_1158, add_107_31_n_119);
  nor g938(add_107_31_n_151, n_1156, n_1161);
  not g939(n_1162, add_107_31_n_84);
  not g940(n_1163, add_107_31_n_154);
  nand g941(add_107_31_n_158, n_1124, add_107_31_n_132);
  nand g942(n_1164, add_107_31_n_166, n_1162);
  nor g943(n_1165, n_1153, add_107_31_n_120);
  nand g944(n_1166, n_1157, add_107_31_n_122);
  not g945(n_1167, n_1166);
  nand g946(n_1168, add_107_31_n_166, n_1167);
  nand g947(n_1169, add_107_31_n_166, n_1163);
  not g948(n_1170, add_107_31_n_91);
  nor g949(n_1171, add_107_31_n_152, n_1170);
  nor g950(n_1172, n_1123, add_107_31_n_154);
  not g951(n_1173, add_107_31_n_93);
  nor g952(add_107_31_n_129, n_1173, add_107_31_n_94);
  not g953(n_1174, add_107_31_n_129);
  nor g954(n_1175, n_1123, add_107_31_n_151);
  nor g955(n_1176, n_1174, n_1175);
  not g956(n_1177, add_107_31_n_97);
  nor g957(n_1178, n_1177, add_107_31_n_130);
  not g958(n_1179, n_1178);
  nor g959(n_1180, add_107_31_n_160, n_1179);
  not g960(n_1181, add_107_31_n_99);
  nor g961(n_1182, n_1181, add_107_31_n_100);
  not g962(n_1183, n_1182);
  nor g963(n_1184, n_1126, add_107_31_n_129);
  nor g964(n_1185, n_1183, n_1184);
  not g965(n_1186, n_1185);
  nor g966(n_1187, add_107_31_n_164, n_1186);
  not g967(n_1188, add_107_31_n_188);
  nand g968(n_1189, add_107_31_n_103, n_1130);
  not g971(n_1190, n_14);
  nor g972(n_1191, rst, n_1115);
  not g973(n_1192, n_1191);
  nand g974(n_1193, n_12, n_1192);
  nor g975(n_1194, n_1190, enb);
  not g976(n_1195, n_1194);
  nor g977(n_1196, n_1190, n_1116);
  not g978(n_1197, n_1196);
  nand g979(n_595, n_1193, n_1195, n_1197);
  not g981(n_1198, n_594);
  nor g982(n_1199, enb, n_1115);
  not g983(n_1200, n_1199);
  nor g984(n_1201, n_1119, State_p[1]);
  not g985(n_1202, n_1201);
  nand g986(n_1203, n_1200, n_1202);
  nand g987(n_598, n_1198, n_1203);
  nand g989(n_1205, n_1130, add_107_31_n_61);
  nand g990(n_1206, n_1120, add_107_31_n_63);
  nand g991(n_1207, n_1127, add_107_31_n_67);
  nand g992(n_1208, n_1135, add_107_31_n_69);
  nand g993(n_1209, n_1138, add_107_31_n_73);
  nand g994(n_1210, n_1144, add_107_31_n_75);
  nand g995(n_1211, n_1162, add_107_31_n_79);
  nand g996(n_1212, n_1160, add_107_31_n_81);
  nand g997(n_1213, n_1157, add_107_31_n_85);
  nand g998(n_1214, n_1154, add_107_31_n_87);
  nand g999(n_1215, n_1121, add_107_31_n_91);
  nand g1000(n_1216, n_1122, add_107_31_n_93);
  nand g1001(n_1217, n_1124, add_107_31_n_97);
  nand g1002(n_1218, n_1125, add_107_31_n_99);
  nand g1003(n_1219, n_1188, add_107_31_n_191);
  nand g1004(n_1220, n_1132, add_107_31_n_59);
  or g2(n_1387, n_1115, State_p[0]);
  not g4(n_8, n_1388);
  or g5(n_10, n_8, rst);
  or g6(n_1697, n_10, State_p[2]);
  or g10(n_1390, n_1389, rst);
  or g11(reg_1[0], n_1390, State_p[2]);
  not g14(n_1392, n_1391);
  or g15(n_1393, n_1392, rst);
  or g16(n_1394, n_1393, State_p[2]);
  not g17(reg_1[2], n_1394);
  not g20(n_1396, n_1395);
  or g21(n_1397, n_1396, rst);
  or g22(n_1398, n_1397, State_p[2]);
  not g23(reg_1[4], n_1398);
  not g26(n_1400, n_1399);
  or g27(n_1401, n_1400, rst);
  or g28(n_1402, n_1401, State_p[2]);
  not g1009(reg_1[3], n_1402);
  not g32(n_1404, n_1403);
  or g33(n_1405, n_1404, rst);
  or g34(n_1406, n_1405, State_p[2]);
  not g35(reg_1[7], n_1406);
  not g38(n_1408, n_1407);
  or g39(n_1409, n_1408, rst);
  or g40(n_1410, n_1409, State_p[2]);
  not g41(reg_1[6], n_1410);
  not g44(n_1412, n_1411);
  or g45(n_1413, n_1412, rst);
  or g46(n_1414, n_1413, State_p[2]);
  not g47(reg_1[5], n_1414);
  not g50(n_1416, n_1415);
  or g51(n_1417, n_1416, rst);
  or g52(n_1418, n_1417, State_p[2]);
  not g53(reg_1[8], n_1418);
  not g56(n_1420, n_1419);
  or g57(n_1421, n_1420, rst);
  or g58(n_1422, n_1421, State_p[2]);
  not g59(reg_1[16], n_1422);
  not g62(n_88, n_87);
  or g63(n_89, n_88, rst);
  or g64(n_90, n_89, State_p[2]);
  not g65(reg_1[15], n_90);
  not g68(n_96, n_95);
  or g69(n_97, n_96, rst);
  or g70(n_98, n_97, State_p[2]);
  not g71(reg_1[14], n_98);
  not g74(n_104, n_103);
  or g75(n_105, n_104, rst);
  or g76(n_106, n_105, State_p[2]);
  not g77(reg_1[13], n_106);
  not g80(n_112, n_111);
  or g81(n_113, n_112, rst);
  or g82(n_114, n_113, State_p[2]);
  not g83(reg_1[12], n_114);
  not g86(n_120, n_119);
  or g87(n_121, n_120, rst);
  or g88(n_122, n_121, State_p[2]);
  not g89(reg_1[11], n_122);
  not g92(n_128, n_127);
  or g93(n_129, n_128, rst);
  or g94(n_130, n_129, State_p[2]);
  not g95(reg_1[10], n_130);
  not g98(n_136, n_135);
  or g99(n_137, n_136, rst);
  or g100(n_138, n_137, State_p[2]);
  not g101(reg_1[9], n_138);
  not g105(n_145, n_144);
  or g106(n_146, n_145, rst);
  or g107(n_147, n_146, State_p[2]);
  not g108(out[2], n_147);
  not g112(n_154, n_153);
  or g113(n_155, n_154, rst);
  or g114(n_156, n_155, State_p[2]);
  not g115(out[1], n_156);
  not g119(n_163, n_162);
  or g120(n_164, n_163, rst);
  or g121(n_165, n_164, State_p[2]);
  not g122(out[0], n_165);
  not g126(n_172, n_171);
  or g127(n_173, n_172, rst);
  or g128(n_174, n_173, State_p[2]);
  not g129(out[4], n_174);
  not g133(n_181, n_180);
  or g134(n_182, n_181, rst);
  or g135(n_183, n_182, State_p[2]);
  not g136(out[3], n_183);
  not g140(n_190, n_189);
  or g141(n_191, n_190, rst);
  or g142(n_192, n_191, State_p[2]);
  not g143(out[7], n_192);
  not g147(n_199, n_198);
  or g148(n_200, n_199, rst);
  or g149(n_201, n_200, State_p[2]);
  not g150(out[6], n_201);
  not g154(n_208, n_207);
  or g155(n_1698, n_208, rst);
  or g156(n_1699, n_1698, State_p[2]);
  not g157(out[5], n_1699);
  not g161(n_1703, n_1702);
  or g162(n_1704, n_1703, rst);
  or g163(n_1705, n_1704, State_p[2]);
  not g164(out[8], n_1705);
  not g168(n_226, n_1708);
  or g169(n_227, n_226, rst);
  or g170(n_228, n_227, State_p[2]);
  not g171(out[16], n_228);
  not g175(n_235, n_234);
  or g176(n_236, n_235, rst);
  or g177(n_237, n_236, State_p[2]);
  not g178(out[15], n_237);
  not g182(n_244, n_243);
  or g183(n_245, n_244, rst);
  or g184(n_246, n_245, State_p[2]);
  not g185(out[14], n_246);
  not g189(n_253, n_252);
  or g190(n_254, n_253, rst);
  or g191(n_255, n_254, State_p[2]);
  not g192(out[13], n_255);
  not g196(n_262, n_261);
  or g197(n_263, n_262, rst);
  or g198(n_264, n_263, State_p[2]);
  not g199(out[12], n_264);
  not g203(n_271, n_270);
  or g204(n_272, n_271, rst);
  or g205(n_273, n_272, State_p[2]);
  not g206(out[11], n_273);
  not g210(n_280, n_279);
  or g211(n_281, n_280, rst);
  or g212(n_282, n_281, State_p[2]);
  not g213(out[10], n_282);
  not g217(n_289, n_288);
  or g218(n_290, n_289, rst);
  or g219(n_291, n_290, State_p[2]);
  not g220(out[9], n_291);
  not g223(n_295, n_294);
  or g224(n_296, n_295, rst);
  or g225(n_297, n_296, State_p[2]);
  not g226(reg_0[2], n_297);
  not g229(n_301, n_300);
  or g230(n_302, n_301, rst);
  or g231(n_303, n_302, State_p[2]);
  not g232(reg_0[1], n_303);
  not g235(n_307, n_306);
  or g236(n_308, n_307, rst);
  or g237(n_309, n_308, State_p[2]);
  not g238(reg_0[0], n_309);
  not g241(n_313, n_312);
  or g242(n_314, n_313, rst);
  or g243(n_315, n_314, State_p[2]);
  not g244(reg_0[4], n_315);
  not g247(n_319, n_318);
  or g248(n_320, n_319, rst);
  or g249(n_321, n_320, State_p[2]);
  not g250(reg_0[3], n_321);
  not g253(n_325, n_324);
  or g254(n_326, n_325, rst);
  or g255(n_327, n_326, State_p[2]);
  not g256(reg_0[7], n_327);
  not g259(n_331, n_330);
  or g260(n_332, n_331, rst);
  or g261(n_333, n_332, State_p[2]);
  not g262(reg_0[6], n_333);
  not g265(n_337, n_336);
  or g266(n_338, n_337, rst);
  or g267(n_339, n_338, State_p[2]);
  not g268(reg_0[5], n_339);
  not g271(n_343, n_342);
  or g272(n_344, n_343, rst);
  or g273(n_345, n_344, State_p[2]);
  not g274(reg_0[8], n_345);
  not g277(n_349, n_348);
  or g278(n_350, n_349, rst);
  or g279(n_351, n_350, State_p[2]);
  not g280(reg_0[16], n_351);
  not g283(n_355, n_354);
  or g284(n_356, n_355, rst);
  or g285(n_357, n_356, State_p[2]);
  not g286(reg_0[15], n_357);
  not g289(n_361, n_360);
  or g290(n_362, n_361, rst);
  or g291(n_363, n_362, State_p[2]);
  not g292(reg_0[14], n_363);
  not g295(n_367, n_366);
  or g296(n_368, n_367, rst);
  or g297(n_369, n_368, State_p[2]);
  not g298(reg_0[13], n_369);
  not g301(n_373, n_372);
  or g302(n_374, n_373, rst);
  or g303(n_375, n_374, State_p[2]);
  not g304(reg_0[12], n_375);
  not g307(n_379, n_378);
  or g308(n_380, n_379, rst);
  or g309(n_381, n_380, State_p[2]);
  not g310(reg_0[11], n_381);
  not g313(n_385, n_384);
  or g314(n_386, n_385, rst);
  or g315(n_387, n_386, State_p[2]);
  not g316(reg_0[10], n_387);
  not g319(n_391, n_390);
  or g320(n_392, n_391, rst);
  or g321(n_393, n_392, State_p[2]);
  not g322(reg_0[9], n_393);
  not g323(n_395, State_p[0]);
  or g324(n_12, n_395, rst);
  or g326(n_14, n_1115, State_p[2]);
  or g327(n_594, rst, State_p[2]);
  not g328(n_1116, State_p[2]);
endmodule

