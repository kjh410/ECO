module top(z,a,shiftCnt);
	input [31:0]a;
	input [4:0]shiftCnt;
	output [31:0]z;
	wire \m21_4_mux_24_18_g32/inv_sel0, \m21_4_mux_24_18_g32/w_0, \m21_4_mux_24_18_g32/w_1, \m21_4_mux_24_18_g31/inv_sel0, \m21_4_mux_24_18_g31/w_0, \m21_4_mux_24_18_g31/w_1, \m21_4_mux_24_18_g30/inv_sel0, \m21_4_mux_24_18_g30/w_0, \m21_4_mux_24_18_g30/w_1, \m21_4_mux_24_18_g29/inv_sel0, \m21_4_mux_24_18_g29/w_0, \m21_4_mux_24_18_g29/w_1, \m21_4_mux_24_18_g28/inv_sel0, \m21_4_mux_24_18_g28/w_0, \m21_4_mux_24_18_g28/w_1, \m21_4_mux_24_18_g27/inv_sel0, \m21_4_mux_24_18_g27/w_0, \m21_4_mux_24_18_g27/w_1, \m21_4_mux_24_18_g26/inv_sel0, \m21_4_mux_24_18_g26/w_0, \m21_4_mux_24_18_g26/w_1, \m21_4_mux_24_18_g25/inv_sel0, \m21_4_mux_24_18_g25/w_0, \m21_4_mux_24_18_g25/w_1, \m21_4_mux_24_18_g24/inv_sel0, \m21_4_mux_24_18_g24/w_0, \m21_4_mux_24_18_g24/w_1, \m21_4_mux_24_18_g23/inv_sel0, \m21_4_mux_24_18_g23/w_0, \m21_4_mux_24_18_g23/w_1, \m21_4_mux_24_18_g22/inv_sel0, \m21_4_mux_24_18_g22/w_0, \m21_4_mux_24_18_g22/w_1, \m21_4_mux_24_18_g21/inv_sel0, \m21_4_mux_24_18_g21/w_0, \m21_4_mux_24_18_g21/w_1, \m21_4_mux_24_18_g20/inv_sel0, \m21_4_mux_24_18_g20/w_0, \m21_4_mux_24_18_g20/w_1, \m21_4_mux_24_18_g19/inv_sel0, \m21_4_mux_24_18_g19/w_0, \m21_4_mux_24_18_g19/w_1, \m21_4_mux_24_18_g18/inv_sel0, \m21_4_mux_24_18_g18/w_0, \m21_4_mux_24_18_g18/w_1, \m21_4_mux_24_18_g17/inv_sel0, \m21_4_mux_24_18_g17/w_0, \m21_4_mux_24_18_g17/w_1, \m21_3_mux_24_18_g9/inv_sel0, \m21_3_mux_24_18_g9/w_0, \m21_3_mux_24_18_g9/w_1, \m21_3_mux_24_18_g32/inv_sel0, \m21_3_mux_24_18_g32/w_0, \m21_3_mux_24_18_g32/w_1, \m21_3_mux_24_18_g31/inv_sel0, \m21_3_mux_24_18_g31/w_0, \m21_3_mux_24_18_g31/w_1, \m21_3_mux_24_18_g30/inv_sel0, \m21_3_mux_24_18_g30/w_0, \m21_3_mux_24_18_g30/w_1, \m21_3_mux_24_18_g29/inv_sel0, \m21_3_mux_24_18_g29/w_0, \m21_3_mux_24_18_g29/w_1, \m21_3_mux_24_18_g28/inv_sel0, \m21_3_mux_24_18_g28/w_0, \m21_3_mux_24_18_g28/w_1, \m21_3_mux_24_18_g27/inv_sel0, \m21_3_mux_24_18_g27/w_0, \m21_3_mux_24_18_g27/w_1, \m21_3_mux_24_18_g26/inv_sel0, \m21_3_mux_24_18_g26/w_0, \m21_3_mux_24_18_g26/w_1, \m21_3_mux_24_18_g25/inv_sel0, \m21_3_mux_24_18_g25/w_0, \m21_3_mux_24_18_g25/w_1, \m21_3_mux_24_18_g24/inv_sel0, \m21_3_mux_24_18_g24/w_0, \m21_3_mux_24_18_g24/w_1, \m21_3_mux_24_18_g23/inv_sel0, \m21_3_mux_24_18_g23/w_0, \m21_3_mux_24_18_g23/w_1, \m21_3_mux_24_18_g22/inv_sel0, \m21_3_mux_24_18_g22/w_0, \m21_3_mux_24_18_g22/w_1, \m21_3_mux_24_18_g21/inv_sel0, \m21_3_mux_24_18_g21/w_0, \m21_3_mux_24_18_g21/w_1, \m21_3_mux_24_18_g20/inv_sel0, \m21_3_mux_24_18_g20/w_0, \m21_3_mux_24_18_g20/w_1, \m21_3_mux_24_18_g19/inv_sel0, \m21_3_mux_24_18_g19/w_0, \m21_3_mux_24_18_g19/w_1, \m21_3_mux_24_18_g18/inv_sel0, \m21_3_mux_24_18_g18/w_0, \m21_3_mux_24_18_g18/w_1, \m21_3_mux_24_18_g17/inv_sel0, \m21_3_mux_24_18_g17/w_0, \m21_3_mux_24_18_g17/w_1, \m21_3_mux_24_18_g16/inv_sel0, \m21_3_mux_24_18_g16/w_0, \m21_3_mux_24_18_g16/w_1, \m21_3_mux_24_18_g15/inv_sel0, \m21_3_mux_24_18_g15/w_0, \m21_3_mux_24_18_g15/w_1, \m21_3_mux_24_18_g14/inv_sel0, \m21_3_mux_24_18_g14/w_0, \m21_3_mux_24_18_g14/w_1, \m21_3_mux_24_18_g13/inv_sel0, \m21_3_mux_24_18_g13/w_0, \m21_3_mux_24_18_g13/w_1, \m21_3_mux_24_18_g12/inv_sel0, \m21_3_mux_24_18_g12/w_0, \m21_3_mux_24_18_g12/w_1, \m21_3_mux_24_18_g11/inv_sel0, \m21_3_mux_24_18_g11/w_0, \m21_3_mux_24_18_g11/w_1, \m21_3_mux_24_18_g10/inv_sel0, \m21_3_mux_24_18_g10/w_0, \m21_3_mux_24_18_g10/w_1, \m21_2_mux_24_18_g9/inv_sel0, \m21_2_mux_24_18_g9/w_0, \m21_2_mux_24_18_g9/w_1, \m21_2_mux_24_18_g8/inv_sel0, \m21_2_mux_24_18_g8/w_0, \m21_2_mux_24_18_g8/w_1, \m21_2_mux_24_18_g7/inv_sel0, \m21_2_mux_24_18_g7/w_0, \m21_2_mux_24_18_g7/w_1, \m21_2_mux_24_18_g6/inv_sel0, \m21_2_mux_24_18_g6/w_0, \m21_2_mux_24_18_g6/w_1, \m21_2_mux_24_18_g5/inv_sel0, \m21_2_mux_24_18_g5/w_0, \m21_2_mux_24_18_g5/w_1, \m21_2_mux_24_18_g4/inv_sel0, \m21_2_mux_24_18_g4/w_0, \m21_2_mux_24_18_g4/w_1, \m21_2_mux_24_18_g32/inv_sel0, \m21_2_mux_24_18_g32/w_0, \m21_2_mux_24_18_g32/w_1, \m21_2_mux_24_18_g31/inv_sel0, \m21_2_mux_24_18_g31/w_0, \m21_2_mux_24_18_g31/w_1, \m21_2_mux_24_18_g30/inv_sel0, \m21_2_mux_24_18_g30/w_0, \m21_2_mux_24_18_g30/w_1, \m21_2_mux_24_18_g3/inv_sel0, \m21_2_mux_24_18_g3/w_0, \m21_2_mux_24_18_g3/w_1, \m21_2_mux_24_18_g29/inv_sel0, \m21_2_mux_24_18_g29/w_0, \m21_2_mux_24_18_g29/w_1, \m21_2_mux_24_18_g28/inv_sel0, \m21_2_mux_24_18_g28/w_0, \m21_2_mux_24_18_g28/w_1, \m21_2_mux_24_18_g27/inv_sel0, \m21_2_mux_24_18_g27/w_0, \m21_2_mux_24_18_g27/w_1, \m21_2_mux_24_18_g26/inv_sel0, \m21_2_mux_24_18_g26/w_0, \m21_2_mux_24_18_g26/w_1, \m21_2_mux_24_18_g25/inv_sel0, \m21_2_mux_24_18_g25/w_0, \m21_2_mux_24_18_g25/w_1, \m21_2_mux_24_18_g24/inv_sel0, \m21_2_mux_24_18_g24/w_0, \m21_2_mux_24_18_g24/w_1, \m21_2_mux_24_18_g23/inv_sel0, \m21_2_mux_24_18_g23/w_0, \m21_2_mux_24_18_g23/w_1, \m21_2_mux_24_18_g22/inv_sel0, \m21_2_mux_24_18_g22/w_0, \m21_2_mux_24_18_g22/w_1, \m21_2_mux_24_18_g21/inv_sel0, \m21_2_mux_24_18_g21/w_0, \m21_2_mux_24_18_g21/w_1, \m21_2_mux_24_18_g20/inv_sel0, \m21_2_mux_24_18_g20/w_0, \m21_2_mux_24_18_g20/w_1, \m21_2_mux_24_18_g2/inv_sel0, \m21_2_mux_24_18_g2/w_0, \m21_2_mux_24_18_g2/w_1, \m21_2_mux_24_18_g19/inv_sel0, \m21_2_mux_24_18_g19/w_0, \m21_2_mux_24_18_g19/w_1, \m21_2_mux_24_18_g18/inv_sel0, \m21_2_mux_24_18_g18/w_0, \m21_2_mux_24_18_g18/w_1, \m21_2_mux_24_18_g17/inv_sel0, \m21_2_mux_24_18_g17/w_0, \m21_2_mux_24_18_g17/w_1, \m21_2_mux_24_18_g16/inv_sel0, \m21_2_mux_24_18_g16/w_0, \m21_2_mux_24_18_g16/w_1, \m21_2_mux_24_18_g15/inv_sel0, \m21_2_mux_24_18_g15/w_0, \m21_2_mux_24_18_g15/w_1, \m21_2_mux_24_18_g14/inv_sel0, \m21_2_mux_24_18_g14/w_0, \m21_2_mux_24_18_g14/w_1, \m21_2_mux_24_18_g13/inv_sel0, \m21_2_mux_24_18_g13/w_0, \m21_2_mux_24_18_g13/w_1, \m21_2_mux_24_18_g12/inv_sel0, \m21_2_mux_24_18_g12/w_0, \m21_2_mux_24_18_g12/w_1, \m21_2_mux_24_18_g11/inv_sel0, \m21_2_mux_24_18_g11/w_0, \m21_2_mux_24_18_g11/w_1, \m21_2_mux_24_18_g10/inv_sel0, \m21_2_mux_24_18_g10/w_0, \m21_2_mux_24_18_g10/w_1, \m21_2_mux_24_18_g1/inv_sel0, \m21_2_mux_24_18_g1/w_0, \m21_2_mux_24_18_g1/w_1, \m21_1_mux_24_18_g9/inv_sel0, \m21_1_mux_24_18_g9/w_0, \m21_1_mux_24_18_g9/w_1, \m21_1_mux_24_18_g8/inv_sel0, \m21_1_mux_24_18_g8/w_0, \m21_1_mux_24_18_g8/w_1, \m21_1_mux_24_18_g7/inv_sel0, \m21_1_mux_24_18_g7/w_0, \m21_1_mux_24_18_g7/w_1, \m21_1_mux_24_18_g6/inv_sel0, \m21_1_mux_24_18_g6/w_0, \m21_1_mux_24_18_g6/w_1, \m21_1_mux_24_18_g5/inv_sel0, \m21_1_mux_24_18_g5/w_0, \m21_1_mux_24_18_g5/w_1, \m21_1_mux_24_18_g4/inv_sel0, \m21_1_mux_24_18_g4/w_0, \m21_1_mux_24_18_g4/w_1, \m21_1_mux_24_18_g32/inv_sel0, \m21_1_mux_24_18_g32/w_0, \m21_1_mux_24_18_g32/w_1, \m21_1_mux_24_18_g31/inv_sel0, \m21_1_mux_24_18_g31/w_0, \m21_1_mux_24_18_g31/w_1, \m21_1_mux_24_18_g30/inv_sel0, \m21_1_mux_24_18_g30/w_0, \m21_1_mux_24_18_g30/w_1, \m21_1_mux_24_18_g3/inv_sel0, \m21_1_mux_24_18_g3/w_0, \m21_1_mux_24_18_g3/w_1, \m21_1_mux_24_18_g29/inv_sel0, \m21_1_mux_24_18_g29/w_0, \m21_1_mux_24_18_g29/w_1, \m21_1_mux_24_18_g28/inv_sel0, \m21_1_mux_24_18_g28/w_0, \m21_1_mux_24_18_g28/w_1, \m21_1_mux_24_18_g27/inv_sel0, \m21_1_mux_24_18_g27/w_0, \m21_1_mux_24_18_g27/w_1, \m21_1_mux_24_18_g26/inv_sel0, \m21_1_mux_24_18_g26/w_0, \m21_1_mux_24_18_g26/w_1, \m21_1_mux_24_18_g25/inv_sel0, \m21_1_mux_24_18_g25/w_0, \m21_1_mux_24_18_g25/w_1, \m21_1_mux_24_18_g24/inv_sel0, \m21_1_mux_24_18_g24/w_0, \m21_1_mux_24_18_g24/w_1, \m21_1_mux_24_18_g23/inv_sel0, \m21_1_mux_24_18_g23/w_0, \m21_1_mux_24_18_g23/w_1, \m21_1_mux_24_18_g22/inv_sel0, \m21_1_mux_24_18_g22/w_0, \m21_1_mux_24_18_g22/w_1, \m21_1_mux_24_18_g21/inv_sel0, \m21_1_mux_24_18_g21/w_0, \m21_1_mux_24_18_g21/w_1, \m21_1_mux_24_18_g20/inv_sel0, \m21_1_mux_24_18_g20/w_0, \m21_1_mux_24_18_g20/w_1, \m21_1_mux_24_18_g2/inv_sel0, \m21_1_mux_24_18_g2/w_0, \m21_1_mux_24_18_g2/w_1, \m21_1_mux_24_18_g19/inv_sel0, \m21_1_mux_24_18_g19/w_0, \m21_1_mux_24_18_g19/w_1, \m21_1_mux_24_18_g18/inv_sel0, \m21_1_mux_24_18_g18/w_0, \m21_1_mux_24_18_g18/w_1, \m21_1_mux_24_18_g17/inv_sel0, \m21_1_mux_24_18_g17/w_0, \m21_1_mux_24_18_g17/w_1, \m21_1_mux_24_18_g16/inv_sel0, \m21_1_mux_24_18_g16/w_0, \m21_1_mux_24_18_g16/w_1, \m21_1_mux_24_18_g15/inv_sel0, \m21_1_mux_24_18_g15/w_0, \m21_1_mux_24_18_g15/w_1, \m21_1_mux_24_18_g14/inv_sel0, \m21_1_mux_24_18_g14/w_0, \m21_1_mux_24_18_g14/w_1, \m21_1_mux_24_18_g13/inv_sel0, \m21_1_mux_24_18_g13/w_0, \m21_1_mux_24_18_g13/w_1, \m21_1_mux_24_18_g12/inv_sel0, \m21_1_mux_24_18_g12/w_0, \m21_1_mux_24_18_g12/w_1, \m21_1_mux_24_18_g11/inv_sel0, \m21_1_mux_24_18_g11/w_0, \m21_1_mux_24_18_g11/w_1, \m21_1_mux_24_18_g10/inv_sel0, \m21_1_mux_24_18_g10/w_0, \m21_1_mux_24_18_g10/w_1, \m21_0_mux_24_18_g9/inv_sel0, \m21_0_mux_24_18_g9/w_0, \m21_0_mux_24_18_g9/w_1, \m21_0_mux_24_18_g8/inv_sel0, \m21_0_mux_24_18_g8/w_0, \m21_0_mux_24_18_g8/w_1, \m21_0_mux_24_18_g7/inv_sel0, \m21_0_mux_24_18_g7/w_0, \m21_0_mux_24_18_g7/w_1, \m21_0_mux_24_18_g6/inv_sel0, \m21_0_mux_24_18_g6/w_0, \m21_0_mux_24_18_g6/w_1, \m21_0_mux_24_18_g5/inv_sel0, \m21_0_mux_24_18_g5/w_0, \m21_0_mux_24_18_g5/w_1, \m21_0_mux_24_18_g4/inv_sel0, \m21_0_mux_24_18_g4/w_0, \m21_0_mux_24_18_g4/w_1, \m21_0_mux_24_18_g32/inv_sel0, \m21_0_mux_24_18_g32/w_0, \m21_0_mux_24_18_g32/w_1, \m21_0_mux_24_18_g31/inv_sel0, \m21_0_mux_24_18_g31/w_0, \m21_0_mux_24_18_g31/w_1, \m21_0_mux_24_18_g30/inv_sel0, \m21_0_mux_24_18_g30/w_0, \m21_0_mux_24_18_g30/w_1, \m21_0_mux_24_18_g3/inv_sel0, \m21_0_mux_24_18_g3/w_0, \m21_0_mux_24_18_g3/w_1, \m21_0_mux_24_18_g29/inv_sel0, \m21_0_mux_24_18_g29/w_0, \m21_0_mux_24_18_g29/w_1, \m21_0_mux_24_18_g28/inv_sel0, \m21_0_mux_24_18_g28/w_0, \m21_0_mux_24_18_g28/w_1, \m21_0_mux_24_18_g27/inv_sel0, \m21_0_mux_24_18_g27/w_0, \m21_0_mux_24_18_g27/w_1, \m21_0_mux_24_18_g26/inv_sel0, \m21_0_mux_24_18_g26/w_0, \m21_0_mux_24_18_g26/w_1, \m21_0_mux_24_18_g25/inv_sel0, \m21_0_mux_24_18_g25/w_0, \m21_0_mux_24_18_g25/w_1, \m21_0_mux_24_18_g24/inv_sel0, \m21_0_mux_24_18_g24/w_0, \m21_0_mux_24_18_g24/w_1, \m21_0_mux_24_18_g23/inv_sel0, \m21_0_mux_24_18_g23/w_0, \m21_0_mux_24_18_g23/w_1, \m21_0_mux_24_18_g22/inv_sel0, \m21_0_mux_24_18_g22/w_0, \m21_0_mux_24_18_g22/w_1, \m21_0_mux_24_18_g21/inv_sel0, \m21_0_mux_24_18_g21/w_0, \m21_0_mux_24_18_g21/w_1, \m21_0_mux_24_18_g20/inv_sel0, \m21_0_mux_24_18_g20/w_0, \m21_0_mux_24_18_g20/w_1, \m21_0_mux_24_18_g2/inv_sel0, \m21_0_mux_24_18_g2/w_0, \m21_0_mux_24_18_g2/w_1, \m21_0_mux_24_18_g19/inv_sel0, \m21_0_mux_24_18_g19/w_0, \m21_0_mux_24_18_g19/w_1, \m21_0_mux_24_18_g18/inv_sel0, \m21_0_mux_24_18_g18/w_0, \m21_0_mux_24_18_g18/w_1, \m21_0_mux_24_18_g17/inv_sel0, \m21_0_mux_24_18_g17/w_0, \m21_0_mux_24_18_g17/w_1, \m21_0_mux_24_18_g16/inv_sel0, \m21_0_mux_24_18_g16/w_0, \m21_0_mux_24_18_g16/w_1, \m21_0_mux_24_18_g15/inv_sel0, \m21_0_mux_24_18_g15/w_0, \m21_0_mux_24_18_g15/w_1, \m21_0_mux_24_18_g14/inv_sel0, \m21_0_mux_24_18_g14/w_0, \m21_0_mux_24_18_g14/w_1, \m21_0_mux_24_18_g13/inv_sel0, \m21_0_mux_24_18_g13/w_0, \m21_0_mux_24_18_g13/w_1, \m21_0_mux_24_18_g12/inv_sel0, \m21_0_mux_24_18_g12/w_0, \m21_0_mux_24_18_g12/w_1, \m21_0_mux_24_18_g11/inv_sel0, \m21_0_mux_24_18_g11/w_0, \m21_0_mux_24_18_g11/w_1, \m21_0_mux_24_18_g10/inv_sel0, \m21_0_mux_24_18_g10/w_0, \m21_0_mux_24_18_g10/w_1, n_228, n_227, n_224, n_223, n_220, n_219, n_216, n_215, n_212, n_211, n_208, n_207, n_204, n_203, n_200, n_199, n_196, n_195, n_192, n_191, n_188, n_187, n_184, n_183, n_180, n_179, n_176, n_175, n_172, n_171, n_168, n_167, n_166, n_165, n_164, n_163, n_160, n_159, n_156, n_155, n_152, n_151, n_148, n_147, n_144, n_143, n_140, n_139, n_136, n_135, n_134, n_133, m21_4_n_81, m21_4_n_80, m21_4_n_79, m21_4_n_78, m21_4_n_77, m21_4_n_76, m21_4_n_75, m21_4_n_74, m21_4_n_73, m21_4_n_72, m21_4_n_71, m21_4_n_70, m21_4_n_69, m21_4_n_68, m21_4_n_67, m21_4_n_66, m21_3_n_89, m21_3_n_88, m21_3_n_87, m21_3_n_86, m21_3_n_85, m21_3_n_84, m21_3_n_83, m21_3_n_82, m21_3_n_81, m21_3_n_80, m21_3_n_79, m21_3_n_78, m21_3_n_77, m21_3_n_76, m21_3_n_75, m21_3_n_74, m21_3_n_73, m21_3_n_72, m21_3_n_71, m21_3_n_70, m21_3_n_69, m21_3_n_68, m21_3_n_67, m21_3_n_66, m21_2_n_97, m21_2_n_96, m21_2_n_95, m21_2_n_94, m21_2_n_93, m21_2_n_92, m21_2_n_91, m21_2_n_90, m21_2_n_89, m21_2_n_88, m21_2_n_87, m21_2_n_86, m21_2_n_85, m21_2_n_84, m21_2_n_83, m21_2_n_82, m21_2_n_81, m21_2_n_80, m21_2_n_79, m21_2_n_78, m21_2_n_77, m21_2_n_76, m21_2_n_75, m21_2_n_74, m21_2_n_73, m21_2_n_72, m21_2_n_71, m21_2_n_70, m21_2_n_69, m21_2_n_68, m21_2_n_67, m21_2_n_66, m21_1_n_96, m21_1_n_95, m21_1_n_94, m21_1_n_93, m21_1_n_92, m21_1_n_91, m21_1_n_90, m21_1_n_89, m21_1_n_88, m21_1_n_87, m21_1_n_86, m21_1_n_85, m21_1_n_84, m21_1_n_83, m21_1_n_82, m21_1_n_81, m21_1_n_80, m21_1_n_79, m21_1_n_78, m21_1_n_77, m21_1_n_76, m21_1_n_75, m21_1_n_74, m21_1_n_73, m21_1_n_72, m21_1_n_71, m21_1_n_70, m21_1_n_69, m21_1_n_68, m21_1_n_67, m21_1_n_66, m21_0_n_96, m21_0_n_95, m21_0_n_94, m21_0_n_93, m21_0_n_92, m21_0_n_91, m21_0_n_90, m21_0_n_89, m21_0_n_88, m21_0_n_87, m21_0_n_86, m21_0_n_85, m21_0_n_84, m21_0_n_83, m21_0_n_82, m21_0_n_81, m21_0_n_80, m21_0_n_79, m21_0_n_78, m21_0_n_77, m21_0_n_76, m21_0_n_75, m21_0_n_74, m21_0_n_73, m21_0_n_72, m21_0_n_71, m21_0_n_70, m21_0_n_69, m21_0_n_68, m21_0_n_67, m21_0_n_66;
	wire [31:0]d3, d2, d1, d0, z;
	wire [4:0]shiftCnt;
	wire [31:0]a;
	wire sub_wire0, w_eco0, w_eco1, w_eco2;

	or \m21_4_mux_24_18_g32/org(m21_4_n_66, \m21_4_mux_24_18_g32/w_0, \m21_4_mux_24_18_g32/w_1);
	and \m21_4_mux_24_18_g32/a_1(\m21_4_mux_24_18_g32/w_1, shiftCnt[4], d3[16]);
	and \m21_4_mux_24_18_g32/a_0(\m21_4_mux_24_18_g32/w_0, \m21_4_mux_24_18_g32/inv_sel0, d3[0]);
	not \m21_4_mux_24_18_g32/i_0(\m21_4_mux_24_18_g32/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g31/org(m21_4_n_67, \m21_4_mux_24_18_g31/w_0, \m21_4_mux_24_18_g31/w_1);
	and \m21_4_mux_24_18_g31/a_1(\m21_4_mux_24_18_g31/w_1, shiftCnt[4], d3[17]);
	and \m21_4_mux_24_18_g31/a_0(\m21_4_mux_24_18_g31/w_0, \m21_4_mux_24_18_g31/inv_sel0, d3[1]);
	not \m21_4_mux_24_18_g31/i_0(\m21_4_mux_24_18_g31/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g30/org(m21_4_n_68, \m21_4_mux_24_18_g30/w_0, \m21_4_mux_24_18_g30/w_1);
	and \m21_4_mux_24_18_g30/a_1(\m21_4_mux_24_18_g30/w_1, shiftCnt[4], d3[18]);
	and \m21_4_mux_24_18_g30/a_0(\m21_4_mux_24_18_g30/w_0, \m21_4_mux_24_18_g30/inv_sel0, d3[2]);
	not \m21_4_mux_24_18_g30/i_0(\m21_4_mux_24_18_g30/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g29/org(m21_4_n_69, \m21_4_mux_24_18_g29/w_0, \m21_4_mux_24_18_g29/w_1);
	and \m21_4_mux_24_18_g29/a_1(\m21_4_mux_24_18_g29/w_1, shiftCnt[4], d3[19]);
	and \m21_4_mux_24_18_g29/a_0(\m21_4_mux_24_18_g29/w_0, \m21_4_mux_24_18_g29/inv_sel0, d3[3]);
	not \m21_4_mux_24_18_g29/i_0(\m21_4_mux_24_18_g29/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g28/org(m21_4_n_70, \m21_4_mux_24_18_g28/w_0, \m21_4_mux_24_18_g28/w_1);
	and \m21_4_mux_24_18_g28/a_1(\m21_4_mux_24_18_g28/w_1, shiftCnt[4], d3[20]);
	and \m21_4_mux_24_18_g28/a_0(\m21_4_mux_24_18_g28/w_0, \m21_4_mux_24_18_g28/inv_sel0, d3[4]);
	not \m21_4_mux_24_18_g28/i_0(\m21_4_mux_24_18_g28/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g27/org(m21_4_n_71, \m21_4_mux_24_18_g27/w_0, \m21_4_mux_24_18_g27/w_1);
	and \m21_4_mux_24_18_g27/a_1(\m21_4_mux_24_18_g27/w_1, shiftCnt[4], d3[21]);
	and \m21_4_mux_24_18_g27/a_0(\m21_4_mux_24_18_g27/w_0, \m21_4_mux_24_18_g27/inv_sel0, d3[5]);
	not \m21_4_mux_24_18_g27/i_0(\m21_4_mux_24_18_g27/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g26/org(m21_4_n_72, \m21_4_mux_24_18_g26/w_0, \m21_4_mux_24_18_g26/w_1);
	and \m21_4_mux_24_18_g26/a_1(\m21_4_mux_24_18_g26/w_1, shiftCnt[4], d3[22]);
	and \m21_4_mux_24_18_g26/a_0(\m21_4_mux_24_18_g26/w_0, \m21_4_mux_24_18_g26/inv_sel0, d3[6]);
	not \m21_4_mux_24_18_g26/i_0(\m21_4_mux_24_18_g26/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g25/org(m21_4_n_73, \m21_4_mux_24_18_g25/w_0, \m21_4_mux_24_18_g25/w_1);
	and \m21_4_mux_24_18_g25/a_1(\m21_4_mux_24_18_g25/w_1, shiftCnt[4], d3[23]);
	and \m21_4_mux_24_18_g25/a_0(\m21_4_mux_24_18_g25/w_0, \m21_4_mux_24_18_g25/inv_sel0, d3[7]);
	not \m21_4_mux_24_18_g25/i_0(\m21_4_mux_24_18_g25/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g24/org(m21_4_n_74, \m21_4_mux_24_18_g24/w_0, \m21_4_mux_24_18_g24/w_1);
	and \m21_4_mux_24_18_g24/a_1(\m21_4_mux_24_18_g24/w_1, shiftCnt[4], d3[24]);
	and \m21_4_mux_24_18_g24/a_0(\m21_4_mux_24_18_g24/w_0, \m21_4_mux_24_18_g24/inv_sel0, d3[8]);
	not \m21_4_mux_24_18_g24/i_0(\m21_4_mux_24_18_g24/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g23/org(m21_4_n_75, \m21_4_mux_24_18_g23/w_0, \m21_4_mux_24_18_g23/w_1);
	and \m21_4_mux_24_18_g23/a_1(\m21_4_mux_24_18_g23/w_1, shiftCnt[4], d3[25]);
	and \m21_4_mux_24_18_g23/a_0(\m21_4_mux_24_18_g23/w_0, \m21_4_mux_24_18_g23/inv_sel0, d3[9]);
	not \m21_4_mux_24_18_g23/i_0(\m21_4_mux_24_18_g23/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g22/org(m21_4_n_76, \m21_4_mux_24_18_g22/w_0, \m21_4_mux_24_18_g22/w_1);
	and \m21_4_mux_24_18_g22/a_1(\m21_4_mux_24_18_g22/w_1, shiftCnt[4], d3[26]);
	and \m21_4_mux_24_18_g22/a_0(\m21_4_mux_24_18_g22/w_0, \m21_4_mux_24_18_g22/inv_sel0, d3[10]);
	not \m21_4_mux_24_18_g22/i_0(\m21_4_mux_24_18_g22/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g21/org(m21_4_n_77, \m21_4_mux_24_18_g21/w_0, \m21_4_mux_24_18_g21/w_1);
	and \m21_4_mux_24_18_g21/a_1(\m21_4_mux_24_18_g21/w_1, shiftCnt[4], d3[27]);
	and \m21_4_mux_24_18_g21/a_0(\m21_4_mux_24_18_g21/w_0, \m21_4_mux_24_18_g21/inv_sel0, d3[11]);
	not \m21_4_mux_24_18_g21/i_0(\m21_4_mux_24_18_g21/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g20/org(m21_4_n_78, \m21_4_mux_24_18_g20/w_0, \m21_4_mux_24_18_g20/w_1);
	and \m21_4_mux_24_18_g20/a_1(\m21_4_mux_24_18_g20/w_1, shiftCnt[4], d3[28]);
	and \m21_4_mux_24_18_g20/a_0(\m21_4_mux_24_18_g20/w_0, \m21_4_mux_24_18_g20/inv_sel0, d3[12]);
	not \m21_4_mux_24_18_g20/i_0(\m21_4_mux_24_18_g20/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g19/org(m21_4_n_79, \m21_4_mux_24_18_g19/w_0, \m21_4_mux_24_18_g19/w_1);
	and \m21_4_mux_24_18_g19/a_1(\m21_4_mux_24_18_g19/w_1, shiftCnt[4], d3[29]);
	and \m21_4_mux_24_18_g19/a_0(\m21_4_mux_24_18_g19/w_0, \m21_4_mux_24_18_g19/inv_sel0, d3[13]);
	not \m21_4_mux_24_18_g19/i_0(\m21_4_mux_24_18_g19/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g18/org(m21_4_n_80, \m21_4_mux_24_18_g18/w_0, \m21_4_mux_24_18_g18/w_1);
	and \m21_4_mux_24_18_g18/a_1(\m21_4_mux_24_18_g18/w_1, shiftCnt[4], d3[30]);
	and \m21_4_mux_24_18_g18/a_0(\m21_4_mux_24_18_g18/w_0, \m21_4_mux_24_18_g18/inv_sel0, d3[14]);
	not \m21_4_mux_24_18_g18/i_0(\m21_4_mux_24_18_g18/inv_sel0, shiftCnt[4]);
	or \m21_4_mux_24_18_g17/org(m21_4_n_81, \m21_4_mux_24_18_g17/w_0, \m21_4_mux_24_18_g17/w_1);
	and \m21_4_mux_24_18_g17/a_1(\m21_4_mux_24_18_g17/w_1, shiftCnt[4], d3[31]);
	and \m21_4_mux_24_18_g17/a_0(\m21_4_mux_24_18_g17/w_0, \m21_4_mux_24_18_g17/inv_sel0, d3[15]);
	not \m21_4_mux_24_18_g17/i_0(\m21_4_mux_24_18_g17/inv_sel0, shiftCnt[4]);
	or \m21_3_mux_24_18_g9/org(m21_3_n_89, \m21_3_mux_24_18_g9/w_0, \m21_3_mux_24_18_g9/w_1);
	and \m21_3_mux_24_18_g9/a_1(\m21_3_mux_24_18_g9/w_1, shiftCnt[3], d2[31]);
	and \m21_3_mux_24_18_g9/a_0(\m21_3_mux_24_18_g9/w_0, \m21_3_mux_24_18_g9/inv_sel0, d2[23]);
	not \m21_3_mux_24_18_g9/i_0(\m21_3_mux_24_18_g9/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g32/org(m21_3_n_66, \m21_3_mux_24_18_g32/w_0, \m21_3_mux_24_18_g32/w_1);
	and \m21_3_mux_24_18_g32/a_1(\m21_3_mux_24_18_g32/w_1, shiftCnt[3], d2[8]);
	and \m21_3_mux_24_18_g32/a_0(\m21_3_mux_24_18_g32/w_0, \m21_3_mux_24_18_g32/inv_sel0, d2[0]);
	not \m21_3_mux_24_18_g32/i_0(\m21_3_mux_24_18_g32/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g31/org(m21_3_n_67, \m21_3_mux_24_18_g31/w_0, \m21_3_mux_24_18_g31/w_1);
	and \m21_3_mux_24_18_g31/a_1(\m21_3_mux_24_18_g31/w_1, shiftCnt[3], d2[9]);
	and \m21_3_mux_24_18_g31/a_0(\m21_3_mux_24_18_g31/w_0, \m21_3_mux_24_18_g31/inv_sel0, d2[1]);
	not \m21_3_mux_24_18_g31/i_0(\m21_3_mux_24_18_g31/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g30/org(m21_3_n_68, \m21_3_mux_24_18_g30/w_0, \m21_3_mux_24_18_g30/w_1);
	and \m21_3_mux_24_18_g30/a_1(\m21_3_mux_24_18_g30/w_1, shiftCnt[3], d2[10]);
	and \m21_3_mux_24_18_g30/a_0(\m21_3_mux_24_18_g30/w_0, \m21_3_mux_24_18_g30/inv_sel0, d2[2]);
	not \m21_3_mux_24_18_g30/i_0(\m21_3_mux_24_18_g30/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g29/org(m21_3_n_69, \m21_3_mux_24_18_g29/w_0, \m21_3_mux_24_18_g29/w_1);
	and \m21_3_mux_24_18_g29/a_1(\m21_3_mux_24_18_g29/w_1, shiftCnt[3], d2[11]);
	and \m21_3_mux_24_18_g29/a_0(\m21_3_mux_24_18_g29/w_0, \m21_3_mux_24_18_g29/inv_sel0, d2[3]);
	not \m21_3_mux_24_18_g29/i_0(\m21_3_mux_24_18_g29/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g28/org(m21_3_n_70, \m21_3_mux_24_18_g28/w_0, \m21_3_mux_24_18_g28/w_1);
	and \m21_3_mux_24_18_g28/a_1(\m21_3_mux_24_18_g28/w_1, shiftCnt[3], d2[12]);
	and \m21_3_mux_24_18_g28/a_0(\m21_3_mux_24_18_g28/w_0, \m21_3_mux_24_18_g28/inv_sel0, d2[4]);
	not \m21_3_mux_24_18_g28/i_0(\m21_3_mux_24_18_g28/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g27/org(m21_3_n_71, \m21_3_mux_24_18_g27/w_0, \m21_3_mux_24_18_g27/w_1);
	and \m21_3_mux_24_18_g27/a_1(\m21_3_mux_24_18_g27/w_1, shiftCnt[3], d2[13]);
	and \m21_3_mux_24_18_g27/a_0(\m21_3_mux_24_18_g27/w_0, \m21_3_mux_24_18_g27/inv_sel0, d2[5]);
	not \m21_3_mux_24_18_g27/i_0(\m21_3_mux_24_18_g27/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g26/org(m21_3_n_72, \m21_3_mux_24_18_g26/w_0, \m21_3_mux_24_18_g26/w_1);
	and \m21_3_mux_24_18_g26/a_1(\m21_3_mux_24_18_g26/w_1, shiftCnt[3], d2[14]);
	and \m21_3_mux_24_18_g26/a_0(\m21_3_mux_24_18_g26/w_0, \m21_3_mux_24_18_g26/inv_sel0, d2[6]);
	not \m21_3_mux_24_18_g26/i_0(\m21_3_mux_24_18_g26/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g25/org(m21_3_n_73, \m21_3_mux_24_18_g25/w_0, \m21_3_mux_24_18_g25/w_1);
	and \m21_3_mux_24_18_g25/a_1(\m21_3_mux_24_18_g25/w_1, shiftCnt[3], d2[15]);
	and \m21_3_mux_24_18_g25/a_0(\m21_3_mux_24_18_g25/w_0, \m21_3_mux_24_18_g25/inv_sel0, d2[7]);
	not \m21_3_mux_24_18_g25/i_0(\m21_3_mux_24_18_g25/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g24/org(m21_3_n_74, \m21_3_mux_24_18_g24/w_0, \m21_3_mux_24_18_g24/w_1);
	and \m21_3_mux_24_18_g24/a_1(\m21_3_mux_24_18_g24/w_1, shiftCnt[3], d2[16]);
	and \m21_3_mux_24_18_g24/a_0(\m21_3_mux_24_18_g24/w_0, \m21_3_mux_24_18_g24/inv_sel0, d2[8]);
	not \m21_3_mux_24_18_g24/i_0(\m21_3_mux_24_18_g24/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g23/org(m21_3_n_75, \m21_3_mux_24_18_g23/w_0, \m21_3_mux_24_18_g23/w_1);
	and \m21_3_mux_24_18_g23/a_1(\m21_3_mux_24_18_g23/w_1, shiftCnt[3], d2[17]);
	and \m21_3_mux_24_18_g23/a_0(\m21_3_mux_24_18_g23/w_0, \m21_3_mux_24_18_g23/inv_sel0, d2[9]);
	not \m21_3_mux_24_18_g23/i_0(\m21_3_mux_24_18_g23/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g22/org(m21_3_n_76, \m21_3_mux_24_18_g22/w_0, \m21_3_mux_24_18_g22/w_1);
	and \m21_3_mux_24_18_g22/a_1(\m21_3_mux_24_18_g22/w_1, shiftCnt[3], d2[18]);
	and \m21_3_mux_24_18_g22/a_0(\m21_3_mux_24_18_g22/w_0, \m21_3_mux_24_18_g22/inv_sel0, d2[10]);
	not \m21_3_mux_24_18_g22/i_0(\m21_3_mux_24_18_g22/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g21/org(m21_3_n_77, \m21_3_mux_24_18_g21/w_0, \m21_3_mux_24_18_g21/w_1);
	and \m21_3_mux_24_18_g21/a_1(\m21_3_mux_24_18_g21/w_1, shiftCnt[3], d2[19]);
	and \m21_3_mux_24_18_g21/a_0(\m21_3_mux_24_18_g21/w_0, \m21_3_mux_24_18_g21/inv_sel0, d2[11]);
	not \m21_3_mux_24_18_g21/i_0(\m21_3_mux_24_18_g21/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g20/org(m21_3_n_78, \m21_3_mux_24_18_g20/w_0, \m21_3_mux_24_18_g20/w_1);
	and \m21_3_mux_24_18_g20/a_1(\m21_3_mux_24_18_g20/w_1, shiftCnt[3], d2[20]);
	and \m21_3_mux_24_18_g20/a_0(\m21_3_mux_24_18_g20/w_0, \m21_3_mux_24_18_g20/inv_sel0, d2[12]);
	not \m21_3_mux_24_18_g20/i_0(\m21_3_mux_24_18_g20/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g19/org(m21_3_n_79, \m21_3_mux_24_18_g19/w_0, \m21_3_mux_24_18_g19/w_1);
	and \m21_3_mux_24_18_g19/a_1(\m21_3_mux_24_18_g19/w_1, shiftCnt[3], d2[21]);
	and \m21_3_mux_24_18_g19/a_0(\m21_3_mux_24_18_g19/w_0, \m21_3_mux_24_18_g19/inv_sel0, d2[13]);
	not \m21_3_mux_24_18_g19/i_0(\m21_3_mux_24_18_g19/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g18/org(m21_3_n_80, \m21_3_mux_24_18_g18/w_0, \m21_3_mux_24_18_g18/w_1);
	and \m21_3_mux_24_18_g18/a_1(\m21_3_mux_24_18_g18/w_1, shiftCnt[3], d2[22]);
	and \m21_3_mux_24_18_g18/a_0(\m21_3_mux_24_18_g18/w_0, \m21_3_mux_24_18_g18/inv_sel0, d2[14]);
	not \m21_3_mux_24_18_g18/i_0(\m21_3_mux_24_18_g18/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g17/org(m21_3_n_81, \m21_3_mux_24_18_g17/w_0, \m21_3_mux_24_18_g17/w_1);
	and \m21_3_mux_24_18_g17/a_1(\m21_3_mux_24_18_g17/w_1, shiftCnt[3], d2[23]);
	and \m21_3_mux_24_18_g17/a_0(\m21_3_mux_24_18_g17/w_0, \m21_3_mux_24_18_g17/inv_sel0, d2[15]);
	not \m21_3_mux_24_18_g17/i_0(\m21_3_mux_24_18_g17/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g16/org(m21_3_n_82, \m21_3_mux_24_18_g16/w_0, \m21_3_mux_24_18_g16/w_1);
	and \m21_3_mux_24_18_g16/a_1(\m21_3_mux_24_18_g16/w_1, shiftCnt[3], d2[24]);
	and \m21_3_mux_24_18_g16/a_0(\m21_3_mux_24_18_g16/w_0, \m21_3_mux_24_18_g16/inv_sel0, d2[16]);
	not \m21_3_mux_24_18_g16/i_0(\m21_3_mux_24_18_g16/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g15/org(m21_3_n_83, \m21_3_mux_24_18_g15/w_0, \m21_3_mux_24_18_g15/w_1);
	and \m21_3_mux_24_18_g15/a_1(\m21_3_mux_24_18_g15/w_1, shiftCnt[3], d2[25]);
	and \m21_3_mux_24_18_g15/a_0(\m21_3_mux_24_18_g15/w_0, \m21_3_mux_24_18_g15/inv_sel0, d2[17]);
	not \m21_3_mux_24_18_g15/i_0(\m21_3_mux_24_18_g15/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g14/org(m21_3_n_84, \m21_3_mux_24_18_g14/w_0, \m21_3_mux_24_18_g14/w_1);
	and \m21_3_mux_24_18_g14/a_1(\m21_3_mux_24_18_g14/w_1, shiftCnt[3], d2[26]);
	and \m21_3_mux_24_18_g14/a_0(\m21_3_mux_24_18_g14/w_0, \m21_3_mux_24_18_g14/inv_sel0, d2[18]);
	not \m21_3_mux_24_18_g14/i_0(\m21_3_mux_24_18_g14/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g13/org(m21_3_n_85, \m21_3_mux_24_18_g13/w_0, \m21_3_mux_24_18_g13/w_1);
	and \m21_3_mux_24_18_g13/a_1(\m21_3_mux_24_18_g13/w_1, shiftCnt[3], d2[27]);
	and \m21_3_mux_24_18_g13/a_0(\m21_3_mux_24_18_g13/w_0, \m21_3_mux_24_18_g13/inv_sel0, d2[19]);
	not \m21_3_mux_24_18_g13/i_0(\m21_3_mux_24_18_g13/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g12/org(m21_3_n_86, \m21_3_mux_24_18_g12/w_0, \m21_3_mux_24_18_g12/w_1);
	and \m21_3_mux_24_18_g12/a_1(\m21_3_mux_24_18_g12/w_1, shiftCnt[3], d2[28]);
	and \m21_3_mux_24_18_g12/a_0(\m21_3_mux_24_18_g12/w_0, \m21_3_mux_24_18_g12/inv_sel0, d2[20]);
	not \m21_3_mux_24_18_g12/i_0(\m21_3_mux_24_18_g12/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g11/org(m21_3_n_87, \m21_3_mux_24_18_g11/w_0, \m21_3_mux_24_18_g11/w_1);
	and \m21_3_mux_24_18_g11/a_1(\m21_3_mux_24_18_g11/w_1, shiftCnt[3], d2[29]);
	and \m21_3_mux_24_18_g11/a_0(\m21_3_mux_24_18_g11/w_0, \m21_3_mux_24_18_g11/inv_sel0, d2[21]);
	not \m21_3_mux_24_18_g11/i_0(\m21_3_mux_24_18_g11/inv_sel0, shiftCnt[3]);
	or \m21_3_mux_24_18_g10/org(m21_3_n_88, \m21_3_mux_24_18_g10/w_0, \m21_3_mux_24_18_g10/w_1);
	and \m21_3_mux_24_18_g10/a_1(\m21_3_mux_24_18_g10/w_1, shiftCnt[3], d2[30]);
	and \m21_3_mux_24_18_g10/a_0(\m21_3_mux_24_18_g10/w_0, \m21_3_mux_24_18_g10/inv_sel0, d2[22]);
	not \m21_3_mux_24_18_g10/i_0(\m21_3_mux_24_18_g10/inv_sel0, shiftCnt[3]);
	or \m21_2_mux_24_18_g9/org(m21_2_n_89, \m21_2_mux_24_18_g9/w_0, \m21_2_mux_24_18_g9/w_1);
	and \m21_2_mux_24_18_g9/a_1(\m21_2_mux_24_18_g9/w_1, shiftCnt[2], d1[27]);
	and \m21_2_mux_24_18_g9/a_0(\m21_2_mux_24_18_g9/w_0, \m21_2_mux_24_18_g9/inv_sel0, d1[23]);
	not \m21_2_mux_24_18_g9/i_0(\m21_2_mux_24_18_g9/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g8/org(m21_2_n_90, \m21_2_mux_24_18_g8/w_0, \m21_2_mux_24_18_g8/w_1);
	and \m21_2_mux_24_18_g8/a_1(\m21_2_mux_24_18_g8/w_1, shiftCnt[2], d1[28]);
	and \m21_2_mux_24_18_g8/a_0(\m21_2_mux_24_18_g8/w_0, \m21_2_mux_24_18_g8/inv_sel0, d1[24]);
	not \m21_2_mux_24_18_g8/i_0(\m21_2_mux_24_18_g8/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g7/org(m21_2_n_91, \m21_2_mux_24_18_g7/w_0, \m21_2_mux_24_18_g7/w_1);
	and \m21_2_mux_24_18_g7/a_1(\m21_2_mux_24_18_g7/w_1, shiftCnt[2], d1[29]);
	and \m21_2_mux_24_18_g7/a_0(\m21_2_mux_24_18_g7/w_0, \m21_2_mux_24_18_g7/inv_sel0, d1[25]);
	not \m21_2_mux_24_18_g7/i_0(\m21_2_mux_24_18_g7/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g6/org(m21_2_n_92, \m21_2_mux_24_18_g6/w_0, \m21_2_mux_24_18_g6/w_1);
	and \m21_2_mux_24_18_g6/a_1(\m21_2_mux_24_18_g6/w_1, shiftCnt[2], d1[30]);
	and \m21_2_mux_24_18_g6/a_0(\m21_2_mux_24_18_g6/w_0, \m21_2_mux_24_18_g6/inv_sel0, d1[26]);
	not \m21_2_mux_24_18_g6/i_0(\m21_2_mux_24_18_g6/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g5/org(m21_2_n_93, \m21_2_mux_24_18_g5/w_0, \m21_2_mux_24_18_g5/w_1);
	and \m21_2_mux_24_18_g5/a_1(\m21_2_mux_24_18_g5/w_1, shiftCnt[2], d1[31]);
	and \m21_2_mux_24_18_g5/a_0(\m21_2_mux_24_18_g5/w_0, \m21_2_mux_24_18_g5/inv_sel0, d1[27]);
	not \m21_2_mux_24_18_g5/i_0(\m21_2_mux_24_18_g5/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g4/org(m21_2_n_94, \m21_2_mux_24_18_g4/w_0, \m21_2_mux_24_18_g4/w_1);
	and \m21_2_mux_24_18_g4/a_1(\m21_2_mux_24_18_g4/w_1, shiftCnt[2], a[31]);
	and \m21_2_mux_24_18_g4/a_0(\m21_2_mux_24_18_g4/w_0, \m21_2_mux_24_18_g4/inv_sel0, d1[28]);
	not \m21_2_mux_24_18_g4/i_0(\m21_2_mux_24_18_g4/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g32/org(m21_2_n_66, \m21_2_mux_24_18_g32/w_0, \m21_2_mux_24_18_g32/w_1);
	and \m21_2_mux_24_18_g32/a_1(\m21_2_mux_24_18_g32/w_1, shiftCnt[2], d1[4]);
	and \m21_2_mux_24_18_g32/a_0(\m21_2_mux_24_18_g32/w_0, \m21_2_mux_24_18_g32/inv_sel0, d1[0]);
	not \m21_2_mux_24_18_g32/i_0(\m21_2_mux_24_18_g32/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g31/org(m21_2_n_67, \m21_2_mux_24_18_g31/w_0, \m21_2_mux_24_18_g31/w_1);
	and \m21_2_mux_24_18_g31/a_1(\m21_2_mux_24_18_g31/w_1, shiftCnt[2], d1[5]);
	and \m21_2_mux_24_18_g31/a_0(\m21_2_mux_24_18_g31/w_0, \m21_2_mux_24_18_g31/inv_sel0, d1[1]);
	not \m21_2_mux_24_18_g31/i_0(\m21_2_mux_24_18_g31/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g30/org(m21_2_n_68, \m21_2_mux_24_18_g30/w_0, \m21_2_mux_24_18_g30/w_1);
	and \m21_2_mux_24_18_g30/a_1(\m21_2_mux_24_18_g30/w_1, shiftCnt[2], d1[6]);
	and \m21_2_mux_24_18_g30/a_0(\m21_2_mux_24_18_g30/w_0, \m21_2_mux_24_18_g30/inv_sel0, d1[2]);
	not \m21_2_mux_24_18_g30/i_0(\m21_2_mux_24_18_g30/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g3/org(m21_2_n_95, \m21_2_mux_24_18_g3/w_0, \m21_2_mux_24_18_g3/w_1);
	and \m21_2_mux_24_18_g3/a_1(\m21_2_mux_24_18_g3/w_1, shiftCnt[2], a[31]);
	and \m21_2_mux_24_18_g3/a_0(\m21_2_mux_24_18_g3/w_0, \m21_2_mux_24_18_g3/inv_sel0, d1[29]);
	not \m21_2_mux_24_18_g3/i_0(\m21_2_mux_24_18_g3/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g29/org(m21_2_n_69, \m21_2_mux_24_18_g29/w_0, \m21_2_mux_24_18_g29/w_1);
	and \m21_2_mux_24_18_g29/a_1(\m21_2_mux_24_18_g29/w_1, shiftCnt[2], d1[7]);
	and \m21_2_mux_24_18_g29/a_0(\m21_2_mux_24_18_g29/w_0, \m21_2_mux_24_18_g29/inv_sel0, d1[3]);
	not \m21_2_mux_24_18_g29/i_0(\m21_2_mux_24_18_g29/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g28/org(m21_2_n_70, \m21_2_mux_24_18_g28/w_0, \m21_2_mux_24_18_g28/w_1);
	and \m21_2_mux_24_18_g28/a_1(\m21_2_mux_24_18_g28/w_1, shiftCnt[2], d1[8]);
	and \m21_2_mux_24_18_g28/a_0(\m21_2_mux_24_18_g28/w_0, \m21_2_mux_24_18_g28/inv_sel0, d1[4]);
	not \m21_2_mux_24_18_g28/i_0(\m21_2_mux_24_18_g28/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g27/org(m21_2_n_71, \m21_2_mux_24_18_g27/w_0, \m21_2_mux_24_18_g27/w_1);
	and \m21_2_mux_24_18_g27/a_1(\m21_2_mux_24_18_g27/w_1, shiftCnt[2], d1[9]);
	and \m21_2_mux_24_18_g27/a_0(\m21_2_mux_24_18_g27/w_0, \m21_2_mux_24_18_g27/inv_sel0, d1[5]);
	not \m21_2_mux_24_18_g27/i_0(\m21_2_mux_24_18_g27/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g26/org(m21_2_n_72, \m21_2_mux_24_18_g26/w_0, \m21_2_mux_24_18_g26/w_1);
	and \m21_2_mux_24_18_g26/a_1(\m21_2_mux_24_18_g26/w_1, shiftCnt[2], d1[10]);
	and \m21_2_mux_24_18_g26/a_0(\m21_2_mux_24_18_g26/w_0, \m21_2_mux_24_18_g26/inv_sel0, d1[6]);
	not \m21_2_mux_24_18_g26/i_0(\m21_2_mux_24_18_g26/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g25/org(m21_2_n_73, \m21_2_mux_24_18_g25/w_0, \m21_2_mux_24_18_g25/w_1);
	and \m21_2_mux_24_18_g25/a_1(\m21_2_mux_24_18_g25/w_1, shiftCnt[2], d1[11]);
	and \m21_2_mux_24_18_g25/a_0(\m21_2_mux_24_18_g25/w_0, \m21_2_mux_24_18_g25/inv_sel0, d1[7]);
	not \m21_2_mux_24_18_g25/i_0(\m21_2_mux_24_18_g25/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g24/org(m21_2_n_74, \m21_2_mux_24_18_g24/w_0, \m21_2_mux_24_18_g24/w_1);
	and \m21_2_mux_24_18_g24/a_1(\m21_2_mux_24_18_g24/w_1, shiftCnt[2], d1[12]);
	and \m21_2_mux_24_18_g24/a_0(\m21_2_mux_24_18_g24/w_0, \m21_2_mux_24_18_g24/inv_sel0, d1[8]);
	not \m21_2_mux_24_18_g24/i_0(\m21_2_mux_24_18_g24/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g23/org(m21_2_n_75, \m21_2_mux_24_18_g23/w_0, \m21_2_mux_24_18_g23/w_1);
	and \m21_2_mux_24_18_g23/a_1(\m21_2_mux_24_18_g23/w_1, shiftCnt[2], d1[13]);
	and \m21_2_mux_24_18_g23/a_0(\m21_2_mux_24_18_g23/w_0, \m21_2_mux_24_18_g23/inv_sel0, d1[9]);
	not \m21_2_mux_24_18_g23/i_0(\m21_2_mux_24_18_g23/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g22/org(m21_2_n_76, \m21_2_mux_24_18_g22/w_0, \m21_2_mux_24_18_g22/w_1);
	and \m21_2_mux_24_18_g22/a_1(\m21_2_mux_24_18_g22/w_1, shiftCnt[2], d1[14]);
	and \m21_2_mux_24_18_g22/a_0(\m21_2_mux_24_18_g22/w_0, \m21_2_mux_24_18_g22/inv_sel0, d1[10]);
	not \m21_2_mux_24_18_g22/i_0(\m21_2_mux_24_18_g22/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g21/org(m21_2_n_77, \m21_2_mux_24_18_g21/w_0, \m21_2_mux_24_18_g21/w_1);
	and \m21_2_mux_24_18_g21/a_1(\m21_2_mux_24_18_g21/w_1, shiftCnt[2], d1[15]);
	and \m21_2_mux_24_18_g21/a_0(\m21_2_mux_24_18_g21/w_0, \m21_2_mux_24_18_g21/inv_sel0, d1[11]);
	not \m21_2_mux_24_18_g21/i_0(\m21_2_mux_24_18_g21/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g20/org(m21_2_n_78, \m21_2_mux_24_18_g20/w_0, \m21_2_mux_24_18_g20/w_1);
	and \m21_2_mux_24_18_g20/a_1(\m21_2_mux_24_18_g20/w_1, shiftCnt[2], d1[16]);
	and \m21_2_mux_24_18_g20/a_0(\m21_2_mux_24_18_g20/w_0, \m21_2_mux_24_18_g20/inv_sel0, d1[12]);
	not \m21_2_mux_24_18_g20/i_0(\m21_2_mux_24_18_g20/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g2/org(m21_2_n_96, \m21_2_mux_24_18_g2/w_0, \m21_2_mux_24_18_g2/w_1);
	and \m21_2_mux_24_18_g2/a_1(\m21_2_mux_24_18_g2/w_1, shiftCnt[2], a[31]);
	and \m21_2_mux_24_18_g2/a_0(\m21_2_mux_24_18_g2/w_0, \m21_2_mux_24_18_g2/inv_sel0, d1[30]);
	not \m21_2_mux_24_18_g2/i_0(\m21_2_mux_24_18_g2/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g19/org(m21_2_n_79, \m21_2_mux_24_18_g19/w_0, \m21_2_mux_24_18_g19/w_1);
	and \m21_2_mux_24_18_g19/a_1(\m21_2_mux_24_18_g19/w_1, shiftCnt[2], d1[17]);
	and \m21_2_mux_24_18_g19/a_0(\m21_2_mux_24_18_g19/w_0, \m21_2_mux_24_18_g19/inv_sel0, d1[13]);
	not \m21_2_mux_24_18_g19/i_0(\m21_2_mux_24_18_g19/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g18/org(m21_2_n_80, \m21_2_mux_24_18_g18/w_0, \m21_2_mux_24_18_g18/w_1);
	and \m21_2_mux_24_18_g18/a_1(\m21_2_mux_24_18_g18/w_1, shiftCnt[2], d1[18]);
	and \m21_2_mux_24_18_g18/a_0(\m21_2_mux_24_18_g18/w_0, \m21_2_mux_24_18_g18/inv_sel0, d1[14]);
	not \m21_2_mux_24_18_g18/i_0(\m21_2_mux_24_18_g18/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g17/org(m21_2_n_81, \m21_2_mux_24_18_g17/w_0, \m21_2_mux_24_18_g17/w_1);
	and \m21_2_mux_24_18_g17/a_1(\m21_2_mux_24_18_g17/w_1, shiftCnt[2], d1[19]);
	and \m21_2_mux_24_18_g17/a_0(\m21_2_mux_24_18_g17/w_0, \m21_2_mux_24_18_g17/inv_sel0, d1[15]);
	not \m21_2_mux_24_18_g17/i_0(\m21_2_mux_24_18_g17/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g16/org(m21_2_n_82, \m21_2_mux_24_18_g16/w_0, \m21_2_mux_24_18_g16/w_1);
	and \m21_2_mux_24_18_g16/a_1(\m21_2_mux_24_18_g16/w_1, shiftCnt[2], d1[20]);
	and \m21_2_mux_24_18_g16/a_0(\m21_2_mux_24_18_g16/w_0, \m21_2_mux_24_18_g16/inv_sel0, d1[16]);
	not \m21_2_mux_24_18_g16/i_0(\m21_2_mux_24_18_g16/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g15/org(m21_2_n_83, \m21_2_mux_24_18_g15/w_0, \m21_2_mux_24_18_g15/w_1);
	and \m21_2_mux_24_18_g15/a_1(\m21_2_mux_24_18_g15/w_1, shiftCnt[2], d1[21]);
	and \m21_2_mux_24_18_g15/a_0(\m21_2_mux_24_18_g15/w_0, \m21_2_mux_24_18_g15/inv_sel0, d1[17]);
	not \m21_2_mux_24_18_g15/i_0(\m21_2_mux_24_18_g15/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g14/org(m21_2_n_84, \m21_2_mux_24_18_g14/w_0, \m21_2_mux_24_18_g14/w_1);
	and \m21_2_mux_24_18_g14/a_1(\m21_2_mux_24_18_g14/w_1, shiftCnt[2], d1[22]);
	and \m21_2_mux_24_18_g14/a_0(\m21_2_mux_24_18_g14/w_0, \m21_2_mux_24_18_g14/inv_sel0, d1[18]);
	not \m21_2_mux_24_18_g14/i_0(\m21_2_mux_24_18_g14/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g13/org(m21_2_n_85, \m21_2_mux_24_18_g13/w_0, \m21_2_mux_24_18_g13/w_1);
	and \m21_2_mux_24_18_g13/a_1(\m21_2_mux_24_18_g13/w_1, shiftCnt[2], d1[23]);
	and \m21_2_mux_24_18_g13/a_0(\m21_2_mux_24_18_g13/w_0, \m21_2_mux_24_18_g13/inv_sel0, d1[19]);
	not \m21_2_mux_24_18_g13/i_0(\m21_2_mux_24_18_g13/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g12/org(m21_2_n_86, \m21_2_mux_24_18_g12/w_0, \m21_2_mux_24_18_g12/w_1);
	and \m21_2_mux_24_18_g12/a_1(\m21_2_mux_24_18_g12/w_1, shiftCnt[2], d1[24]);
	and \m21_2_mux_24_18_g12/a_0(\m21_2_mux_24_18_g12/w_0, \m21_2_mux_24_18_g12/inv_sel0, d1[20]);
	not \m21_2_mux_24_18_g12/i_0(\m21_2_mux_24_18_g12/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g11/org(m21_2_n_87, \m21_2_mux_24_18_g11/w_0, \m21_2_mux_24_18_g11/w_1);
	and \m21_2_mux_24_18_g11/a_1(\m21_2_mux_24_18_g11/w_1, shiftCnt[2], d1[25]);
	and \m21_2_mux_24_18_g11/a_0(\m21_2_mux_24_18_g11/w_0, \m21_2_mux_24_18_g11/inv_sel0, d1[21]);
	not \m21_2_mux_24_18_g11/i_0(\m21_2_mux_24_18_g11/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g10/org(m21_2_n_88, \m21_2_mux_24_18_g10/w_0, \m21_2_mux_24_18_g10/w_1);
	and \m21_2_mux_24_18_g10/a_1(\m21_2_mux_24_18_g10/w_1, shiftCnt[2], d1[26]);
	and \m21_2_mux_24_18_g10/a_0(\m21_2_mux_24_18_g10/w_0, \m21_2_mux_24_18_g10/inv_sel0, d1[22]);
	not \m21_2_mux_24_18_g10/i_0(\m21_2_mux_24_18_g10/inv_sel0, shiftCnt[2]);
	or \m21_2_mux_24_18_g1/org(m21_2_n_97, \m21_2_mux_24_18_g1/w_0, \m21_2_mux_24_18_g1/w_1);
	and \m21_2_mux_24_18_g1/a_1(\m21_2_mux_24_18_g1/w_1, shiftCnt[2], a[31]);
	and \m21_2_mux_24_18_g1/a_0(\m21_2_mux_24_18_g1/w_0, \m21_2_mux_24_18_g1/inv_sel0, d1[31]);
	not \m21_2_mux_24_18_g1/i_0(\m21_2_mux_24_18_g1/inv_sel0, shiftCnt[2]);
	or \m21_1_mux_24_18_g9/org(m21_1_n_89, \m21_1_mux_24_18_g9/w_0, \m21_1_mux_24_18_g9/w_1);
	and \m21_1_mux_24_18_g9/a_1(\m21_1_mux_24_18_g9/w_1, shiftCnt[1], d0[25]);
	and \m21_1_mux_24_18_g9/a_0(\m21_1_mux_24_18_g9/w_0, \m21_1_mux_24_18_g9/inv_sel0, d0[23]);
	not \m21_1_mux_24_18_g9/i_0(\m21_1_mux_24_18_g9/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g8/org(m21_1_n_90, \m21_1_mux_24_18_g8/w_0, \m21_1_mux_24_18_g8/w_1);
	and \m21_1_mux_24_18_g8/a_1(\m21_1_mux_24_18_g8/w_1, shiftCnt[1], d0[26]);
	and \m21_1_mux_24_18_g8/a_0(\m21_1_mux_24_18_g8/w_0, \m21_1_mux_24_18_g8/inv_sel0, d0[24]);
	not \m21_1_mux_24_18_g8/i_0(\m21_1_mux_24_18_g8/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g7/org(m21_1_n_91, \m21_1_mux_24_18_g7/w_0, \m21_1_mux_24_18_g7/w_1);
	and \m21_1_mux_24_18_g7/a_1(\m21_1_mux_24_18_g7/w_1, shiftCnt[1], d0[27]);
	and \m21_1_mux_24_18_g7/a_0(\m21_1_mux_24_18_g7/w_0, \m21_1_mux_24_18_g7/inv_sel0, d0[25]);
	not \m21_1_mux_24_18_g7/i_0(\m21_1_mux_24_18_g7/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g6/org(m21_1_n_92, \m21_1_mux_24_18_g6/w_0, \m21_1_mux_24_18_g6/w_1);
	and \m21_1_mux_24_18_g6/a_1(\m21_1_mux_24_18_g6/w_1, shiftCnt[1], d0[28]);
	and \m21_1_mux_24_18_g6/a_0(\m21_1_mux_24_18_g6/w_0, \m21_1_mux_24_18_g6/inv_sel0, d0[26]);
	not \m21_1_mux_24_18_g6/i_0(\m21_1_mux_24_18_g6/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g5/org(m21_1_n_93, \m21_1_mux_24_18_g5/w_0, \m21_1_mux_24_18_g5/w_1);
	and \m21_1_mux_24_18_g5/a_1(\m21_1_mux_24_18_g5/w_1, shiftCnt[1], d0[29]);
	and \m21_1_mux_24_18_g5/a_0(\m21_1_mux_24_18_g5/w_0, \m21_1_mux_24_18_g5/inv_sel0, d0[27]);
	not \m21_1_mux_24_18_g5/i_0(\m21_1_mux_24_18_g5/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g4/org(m21_1_n_94, \m21_1_mux_24_18_g4/w_0, \m21_1_mux_24_18_g4/w_1);
	and \m21_1_mux_24_18_g4/a_1(\m21_1_mux_24_18_g4/w_1, shiftCnt[1], d0[30]);
	and \m21_1_mux_24_18_g4/a_0(\m21_1_mux_24_18_g4/w_0, \m21_1_mux_24_18_g4/inv_sel0, d0[28]);
	not \m21_1_mux_24_18_g4/i_0(\m21_1_mux_24_18_g4/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g32/org(m21_1_n_66, \m21_1_mux_24_18_g32/w_0, \m21_1_mux_24_18_g32/w_1);
	and \m21_1_mux_24_18_g32/a_1(\m21_1_mux_24_18_g32/w_1, shiftCnt[1], d0[2]);
	and \m21_1_mux_24_18_g32/a_0(\m21_1_mux_24_18_g32/w_0, \m21_1_mux_24_18_g32/inv_sel0, d0[0]);
	not \m21_1_mux_24_18_g32/i_0(\m21_1_mux_24_18_g32/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g31/org(m21_1_n_67, \m21_1_mux_24_18_g31/w_0, \m21_1_mux_24_18_g31/w_1);
	and \m21_1_mux_24_18_g31/a_1(\m21_1_mux_24_18_g31/w_1, shiftCnt[1], d0[3]);
	and \m21_1_mux_24_18_g31/a_0(\m21_1_mux_24_18_g31/w_0, \m21_1_mux_24_18_g31/inv_sel0, d0[1]);
	not \m21_1_mux_24_18_g31/i_0(\m21_1_mux_24_18_g31/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g30/org(m21_1_n_68, \m21_1_mux_24_18_g30/w_0, \m21_1_mux_24_18_g30/w_1);
	and \m21_1_mux_24_18_g30/a_1(\m21_1_mux_24_18_g30/w_1, shiftCnt[1], d0[4]);
	and \m21_1_mux_24_18_g30/a_0(\m21_1_mux_24_18_g30/w_0, \m21_1_mux_24_18_g30/inv_sel0, d0[2]);
	not \m21_1_mux_24_18_g30/i_0(\m21_1_mux_24_18_g30/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g3/org(m21_1_n_95, \m21_1_mux_24_18_g3/w_0, \m21_1_mux_24_18_g3/w_1);
	and \m21_1_mux_24_18_g3/a_1(\m21_1_mux_24_18_g3/w_1, shiftCnt[1], d0[31]);
	and \m21_1_mux_24_18_g3/a_0(\m21_1_mux_24_18_g3/w_0, \m21_1_mux_24_18_g3/inv_sel0, d0[29]);
	not \m21_1_mux_24_18_g3/i_0(\m21_1_mux_24_18_g3/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g29/org(m21_1_n_69, \m21_1_mux_24_18_g29/w_0, \m21_1_mux_24_18_g29/w_1);
	and \m21_1_mux_24_18_g29/a_1(\m21_1_mux_24_18_g29/w_1, shiftCnt[1], d0[5]);
	and \m21_1_mux_24_18_g29/a_0(\m21_1_mux_24_18_g29/w_0, \m21_1_mux_24_18_g29/inv_sel0, d0[3]);
	not \m21_1_mux_24_18_g29/i_0(\m21_1_mux_24_18_g29/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g28/org(m21_1_n_70, \m21_1_mux_24_18_g28/w_0, \m21_1_mux_24_18_g28/w_1);
	and \m21_1_mux_24_18_g28/a_1(\m21_1_mux_24_18_g28/w_1, shiftCnt[1], d0[6]);
	and \m21_1_mux_24_18_g28/a_0(\m21_1_mux_24_18_g28/w_0, \m21_1_mux_24_18_g28/inv_sel0, d0[4]);
	not \m21_1_mux_24_18_g28/i_0(\m21_1_mux_24_18_g28/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g27/org(m21_1_n_71, \m21_1_mux_24_18_g27/w_0, \m21_1_mux_24_18_g27/w_1);
	and \m21_1_mux_24_18_g27/a_1(\m21_1_mux_24_18_g27/w_1, shiftCnt[1], d0[7]);
	and \m21_1_mux_24_18_g27/a_0(\m21_1_mux_24_18_g27/w_0, \m21_1_mux_24_18_g27/inv_sel0, d0[5]);
	not \m21_1_mux_24_18_g27/i_0(\m21_1_mux_24_18_g27/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g26/org(m21_1_n_72, \m21_1_mux_24_18_g26/w_0, \m21_1_mux_24_18_g26/w_1);
	and \m21_1_mux_24_18_g26/a_1(\m21_1_mux_24_18_g26/w_1, shiftCnt[1], d0[8]);
	and \m21_1_mux_24_18_g26/a_0(\m21_1_mux_24_18_g26/w_0, \m21_1_mux_24_18_g26/inv_sel0, d0[6]);
	not \m21_1_mux_24_18_g26/i_0(\m21_1_mux_24_18_g26/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g25/org(m21_1_n_73, \m21_1_mux_24_18_g25/w_0, \m21_1_mux_24_18_g25/w_1);
	and \m21_1_mux_24_18_g25/a_1(\m21_1_mux_24_18_g25/w_1, shiftCnt[1], d0[9]);
	and \m21_1_mux_24_18_g25/a_0(\m21_1_mux_24_18_g25/w_0, \m21_1_mux_24_18_g25/inv_sel0, d0[7]);
	not \m21_1_mux_24_18_g25/i_0(\m21_1_mux_24_18_g25/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g24/org(m21_1_n_74, \m21_1_mux_24_18_g24/w_0, \m21_1_mux_24_18_g24/w_1);
	and \m21_1_mux_24_18_g24/a_1(\m21_1_mux_24_18_g24/w_1, shiftCnt[1], d0[10]);
	and \m21_1_mux_24_18_g24/a_0(\m21_1_mux_24_18_g24/w_0, \m21_1_mux_24_18_g24/inv_sel0, d0[8]);
	not \m21_1_mux_24_18_g24/i_0(\m21_1_mux_24_18_g24/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g23/org(m21_1_n_75, \m21_1_mux_24_18_g23/w_0, \m21_1_mux_24_18_g23/w_1);
	and \m21_1_mux_24_18_g23/a_1(\m21_1_mux_24_18_g23/w_1, shiftCnt[1], d0[11]);
	and \m21_1_mux_24_18_g23/a_0(\m21_1_mux_24_18_g23/w_0, \m21_1_mux_24_18_g23/inv_sel0, d0[9]);
	not \m21_1_mux_24_18_g23/i_0(\m21_1_mux_24_18_g23/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g22/org(m21_1_n_76, \m21_1_mux_24_18_g22/w_0, \m21_1_mux_24_18_g22/w_1);
	and \m21_1_mux_24_18_g22/a_1(\m21_1_mux_24_18_g22/w_1, shiftCnt[1], d0[12]);
	and \m21_1_mux_24_18_g22/a_0(\m21_1_mux_24_18_g22/w_0, \m21_1_mux_24_18_g22/inv_sel0, d0[10]);
	not \m21_1_mux_24_18_g22/i_0(\m21_1_mux_24_18_g22/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g21/org(m21_1_n_77, \m21_1_mux_24_18_g21/w_0, \m21_1_mux_24_18_g21/w_1);
	and \m21_1_mux_24_18_g21/a_1(\m21_1_mux_24_18_g21/w_1, shiftCnt[1], d0[13]);
	and \m21_1_mux_24_18_g21/a_0(\m21_1_mux_24_18_g21/w_0, \m21_1_mux_24_18_g21/inv_sel0, d0[11]);
	not \m21_1_mux_24_18_g21/i_0(\m21_1_mux_24_18_g21/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g20/org(m21_1_n_78, \m21_1_mux_24_18_g20/w_0, \m21_1_mux_24_18_g20/w_1);
	and \m21_1_mux_24_18_g20/a_1(\m21_1_mux_24_18_g20/w_1, shiftCnt[1], d0[14]);
	and \m21_1_mux_24_18_g20/a_0(\m21_1_mux_24_18_g20/w_0, \m21_1_mux_24_18_g20/inv_sel0, d0[12]);
	not \m21_1_mux_24_18_g20/i_0(\m21_1_mux_24_18_g20/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g2/org(m21_1_n_96, \m21_1_mux_24_18_g2/w_0, \m21_1_mux_24_18_g2/w_1);
	and \m21_1_mux_24_18_g2/a_1(\m21_1_mux_24_18_g2/w_1, shiftCnt[1], a[31]);
	and \m21_1_mux_24_18_g2/a_0(\m21_1_mux_24_18_g2/w_0, \m21_1_mux_24_18_g2/inv_sel0, d0[30]);
	not \m21_1_mux_24_18_g2/i_0(\m21_1_mux_24_18_g2/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g19/org(m21_1_n_79, \m21_1_mux_24_18_g19/w_0, \m21_1_mux_24_18_g19/w_1);
	and \m21_1_mux_24_18_g19/a_1(\m21_1_mux_24_18_g19/w_1, shiftCnt[1], d0[15]);
	and \m21_1_mux_24_18_g19/a_0(\m21_1_mux_24_18_g19/w_0, \m21_1_mux_24_18_g19/inv_sel0, d0[13]);
	not \m21_1_mux_24_18_g19/i_0(\m21_1_mux_24_18_g19/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g18/org(m21_1_n_80, \m21_1_mux_24_18_g18/w_0, \m21_1_mux_24_18_g18/w_1);
	and \m21_1_mux_24_18_g18/a_1(\m21_1_mux_24_18_g18/w_1, shiftCnt[1], d0[16]);
	and \m21_1_mux_24_18_g18/a_0(\m21_1_mux_24_18_g18/w_0, \m21_1_mux_24_18_g18/inv_sel0, d0[14]);
	not \m21_1_mux_24_18_g18/i_0(\m21_1_mux_24_18_g18/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g17/org(m21_1_n_81, \m21_1_mux_24_18_g17/w_0, \m21_1_mux_24_18_g17/w_1);
	and \m21_1_mux_24_18_g17/a_1(\m21_1_mux_24_18_g17/w_1, shiftCnt[1], d0[17]);
	and \m21_1_mux_24_18_g17/a_0(\m21_1_mux_24_18_g17/w_0, \m21_1_mux_24_18_g17/inv_sel0, d0[15]);
	not \m21_1_mux_24_18_g17/i_0(\m21_1_mux_24_18_g17/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g16/org(m21_1_n_82, \m21_1_mux_24_18_g16/w_0, \m21_1_mux_24_18_g16/w_1);
	and \m21_1_mux_24_18_g16/a_1(\m21_1_mux_24_18_g16/w_1, shiftCnt[1], d0[18]);
	and \m21_1_mux_24_18_g16/a_0(\m21_1_mux_24_18_g16/w_0, \m21_1_mux_24_18_g16/inv_sel0, d0[16]);
	not \m21_1_mux_24_18_g16/i_0(\m21_1_mux_24_18_g16/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g15/org(m21_1_n_83, \m21_1_mux_24_18_g15/w_0, \m21_1_mux_24_18_g15/w_1);
	and \m21_1_mux_24_18_g15/a_1(\m21_1_mux_24_18_g15/w_1, shiftCnt[1], d0[19]);
	and \m21_1_mux_24_18_g15/a_0(\m21_1_mux_24_18_g15/w_0, \m21_1_mux_24_18_g15/inv_sel0, d0[17]);
	not \m21_1_mux_24_18_g15/i_0(\m21_1_mux_24_18_g15/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g14/org(m21_1_n_84, \m21_1_mux_24_18_g14/w_0, \m21_1_mux_24_18_g14/w_1);
	and \m21_1_mux_24_18_g14/a_1(\m21_1_mux_24_18_g14/w_1, shiftCnt[1], d0[20]);
	and \m21_1_mux_24_18_g14/a_0(\m21_1_mux_24_18_g14/w_0, \m21_1_mux_24_18_g14/inv_sel0, d0[18]);
	not \m21_1_mux_24_18_g14/i_0(\m21_1_mux_24_18_g14/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g13/org(m21_1_n_85, \m21_1_mux_24_18_g13/w_0, \m21_1_mux_24_18_g13/w_1);
	and \m21_1_mux_24_18_g13/a_1(\m21_1_mux_24_18_g13/w_1, shiftCnt[1], d0[21]);
	and \m21_1_mux_24_18_g13/a_0(\m21_1_mux_24_18_g13/w_0, \m21_1_mux_24_18_g13/inv_sel0, d0[19]);
	not \m21_1_mux_24_18_g13/i_0(\m21_1_mux_24_18_g13/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g12/org(m21_1_n_86, \m21_1_mux_24_18_g12/w_0, \m21_1_mux_24_18_g12/w_1);
	and \m21_1_mux_24_18_g12/a_1(\m21_1_mux_24_18_g12/w_1, shiftCnt[1], d0[22]);
	and \m21_1_mux_24_18_g12/a_0(\m21_1_mux_24_18_g12/w_0, \m21_1_mux_24_18_g12/inv_sel0, d0[20]);
	not \m21_1_mux_24_18_g12/i_0(\m21_1_mux_24_18_g12/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g11/org(m21_1_n_87, \m21_1_mux_24_18_g11/w_0, \m21_1_mux_24_18_g11/w_1);
	and \m21_1_mux_24_18_g11/a_1(\m21_1_mux_24_18_g11/w_1, shiftCnt[1], d0[23]);
	and \m21_1_mux_24_18_g11/a_0(\m21_1_mux_24_18_g11/w_0, \m21_1_mux_24_18_g11/inv_sel0, d0[21]);
	not \m21_1_mux_24_18_g11/i_0(\m21_1_mux_24_18_g11/inv_sel0, shiftCnt[1]);
	or \m21_1_mux_24_18_g10/org(m21_1_n_88, \m21_1_mux_24_18_g10/w_0, \m21_1_mux_24_18_g10/w_1);
	and \m21_1_mux_24_18_g10/a_1(\m21_1_mux_24_18_g10/w_1, shiftCnt[1], d0[24]);
	and \m21_1_mux_24_18_g10/a_0(\m21_1_mux_24_18_g10/w_0, \m21_1_mux_24_18_g10/inv_sel0, d0[22]);
	not \m21_1_mux_24_18_g10/i_0(\m21_1_mux_24_18_g10/inv_sel0, shiftCnt[1]);
	or \m21_0_mux_24_18_g9/org(m21_0_n_89, \m21_0_mux_24_18_g9/w_0, \m21_0_mux_24_18_g9/w_1);
	and \m21_0_mux_24_18_g9/a_1(\m21_0_mux_24_18_g9/w_1, shiftCnt[0], a[24]);
	and \m21_0_mux_24_18_g9/a_0(\m21_0_mux_24_18_g9/w_0, \m21_0_mux_24_18_g9/inv_sel0, a[23]);
	not \m21_0_mux_24_18_g9/i_0(\m21_0_mux_24_18_g9/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g8/org(m21_0_n_90, \m21_0_mux_24_18_g8/w_0, \m21_0_mux_24_18_g8/w_1);
	and \m21_0_mux_24_18_g8/a_1(\m21_0_mux_24_18_g8/w_1, shiftCnt[0], a[25]);
	and \m21_0_mux_24_18_g8/a_0(\m21_0_mux_24_18_g8/w_0, \m21_0_mux_24_18_g8/inv_sel0, a[24]);
	not \m21_0_mux_24_18_g8/i_0(\m21_0_mux_24_18_g8/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g7/org(m21_0_n_91, \m21_0_mux_24_18_g7/w_0, \m21_0_mux_24_18_g7/w_1);
	and \m21_0_mux_24_18_g7/a_1(\m21_0_mux_24_18_g7/w_1, shiftCnt[0], a[26]);
	and \m21_0_mux_24_18_g7/a_0(\m21_0_mux_24_18_g7/w_0, \m21_0_mux_24_18_g7/inv_sel0, a[25]);
	not \m21_0_mux_24_18_g7/i_0(\m21_0_mux_24_18_g7/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g6/org(m21_0_n_92, \m21_0_mux_24_18_g6/w_0, \m21_0_mux_24_18_g6/w_1);
	and \m21_0_mux_24_18_g6/a_1(\m21_0_mux_24_18_g6/w_1, shiftCnt[0], a[27]);
	and \m21_0_mux_24_18_g6/a_0(\m21_0_mux_24_18_g6/w_0, \m21_0_mux_24_18_g6/inv_sel0, a[26]);
	not \m21_0_mux_24_18_g6/i_0(\m21_0_mux_24_18_g6/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g5/org(m21_0_n_93, \m21_0_mux_24_18_g5/w_0, \m21_0_mux_24_18_g5/w_1);
	and \m21_0_mux_24_18_g5/a_1(\m21_0_mux_24_18_g5/w_1, shiftCnt[0], a[28]);
	and \m21_0_mux_24_18_g5/a_0(\m21_0_mux_24_18_g5/w_0, \m21_0_mux_24_18_g5/inv_sel0, a[27]);
	not \m21_0_mux_24_18_g5/i_0(\m21_0_mux_24_18_g5/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g4/org(m21_0_n_94, \m21_0_mux_24_18_g4/w_0, \m21_0_mux_24_18_g4/w_1);
	and \m21_0_mux_24_18_g4/a_1(\m21_0_mux_24_18_g4/w_1, shiftCnt[0], a[29]);
	and \m21_0_mux_24_18_g4/a_0(\m21_0_mux_24_18_g4/w_0, \m21_0_mux_24_18_g4/inv_sel0, a[28]);
	not \m21_0_mux_24_18_g4/i_0(\m21_0_mux_24_18_g4/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g32/org(m21_0_n_66, \m21_0_mux_24_18_g32/w_0, \m21_0_mux_24_18_g32/w_1);
	and \m21_0_mux_24_18_g32/a_1(\m21_0_mux_24_18_g32/w_1, shiftCnt[0], a[1]);
	and \m21_0_mux_24_18_g32/a_0(\m21_0_mux_24_18_g32/w_0, \m21_0_mux_24_18_g32/inv_sel0, a[0]);
	not \m21_0_mux_24_18_g32/i_0(\m21_0_mux_24_18_g32/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g31/org(m21_0_n_67, \m21_0_mux_24_18_g31/w_0, \m21_0_mux_24_18_g31/w_1);
	and \m21_0_mux_24_18_g31/a_1(\m21_0_mux_24_18_g31/w_1, shiftCnt[0], a[2]);
	and \m21_0_mux_24_18_g31/a_0(\m21_0_mux_24_18_g31/w_0, \m21_0_mux_24_18_g31/inv_sel0, a[1]);
	not \m21_0_mux_24_18_g31/i_0(\m21_0_mux_24_18_g31/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g30/org(m21_0_n_68, \m21_0_mux_24_18_g30/w_0, \m21_0_mux_24_18_g30/w_1);
	and \m21_0_mux_24_18_g30/a_1(\m21_0_mux_24_18_g30/w_1, shiftCnt[0], a[3]);
	and \m21_0_mux_24_18_g30/a_0(\m21_0_mux_24_18_g30/w_0, \m21_0_mux_24_18_g30/inv_sel0, a[2]);
	not \m21_0_mux_24_18_g30/i_0(\m21_0_mux_24_18_g30/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g3/org(m21_0_n_95, \m21_0_mux_24_18_g3/w_0, \m21_0_mux_24_18_g3/w_1);
	and \m21_0_mux_24_18_g3/a_1(\m21_0_mux_24_18_g3/w_1, shiftCnt[0], a[30]);
	and \m21_0_mux_24_18_g3/a_0(\m21_0_mux_24_18_g3/w_0, \m21_0_mux_24_18_g3/inv_sel0, a[29]);
	not \m21_0_mux_24_18_g3/i_0(\m21_0_mux_24_18_g3/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g29/org(m21_0_n_69, \m21_0_mux_24_18_g29/w_0, \m21_0_mux_24_18_g29/w_1);
	and \m21_0_mux_24_18_g29/a_1(\m21_0_mux_24_18_g29/w_1, shiftCnt[0], a[4]);
	and \m21_0_mux_24_18_g29/a_0(\m21_0_mux_24_18_g29/w_0, \m21_0_mux_24_18_g29/inv_sel0, a[3]);
	not \m21_0_mux_24_18_g29/i_0(\m21_0_mux_24_18_g29/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g28/org(m21_0_n_70, \m21_0_mux_24_18_g28/w_0, \m21_0_mux_24_18_g28/w_1);
	and \m21_0_mux_24_18_g28/a_1(\m21_0_mux_24_18_g28/w_1, shiftCnt[0], a[5]);
	and \m21_0_mux_24_18_g28/a_0(\m21_0_mux_24_18_g28/w_0, \m21_0_mux_24_18_g28/inv_sel0, a[4]);
	not \m21_0_mux_24_18_g28/i_0(\m21_0_mux_24_18_g28/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g27/org(m21_0_n_71, \m21_0_mux_24_18_g27/w_0, \m21_0_mux_24_18_g27/w_1);
	and \m21_0_mux_24_18_g27/a_1(\m21_0_mux_24_18_g27/w_1, shiftCnt[0], a[6]);
	and \m21_0_mux_24_18_g27/a_0(\m21_0_mux_24_18_g27/w_0, \m21_0_mux_24_18_g27/inv_sel0, a[5]);
	not \m21_0_mux_24_18_g27/i_0(\m21_0_mux_24_18_g27/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g26/org(m21_0_n_72, \m21_0_mux_24_18_g26/w_0, \m21_0_mux_24_18_g26/w_1);
	and \m21_0_mux_24_18_g26/a_1(\m21_0_mux_24_18_g26/w_1, shiftCnt[0], a[7]);
	and \m21_0_mux_24_18_g26/a_0(\m21_0_mux_24_18_g26/w_0, \m21_0_mux_24_18_g26/inv_sel0, a[6]);
	not \m21_0_mux_24_18_g26/i_0(\m21_0_mux_24_18_g26/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g25/org(m21_0_n_73, \m21_0_mux_24_18_g25/w_0, \m21_0_mux_24_18_g25/w_1);
	and \m21_0_mux_24_18_g25/a_1(\m21_0_mux_24_18_g25/w_1, shiftCnt[0], a[8]);
	and \m21_0_mux_24_18_g25/a_0(\m21_0_mux_24_18_g25/w_0, \m21_0_mux_24_18_g25/inv_sel0, a[7]);
	not \m21_0_mux_24_18_g25/i_0(\m21_0_mux_24_18_g25/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g24/org(m21_0_n_74, \m21_0_mux_24_18_g24/w_0, \m21_0_mux_24_18_g24/w_1);
	and \m21_0_mux_24_18_g24/a_1(\m21_0_mux_24_18_g24/w_1, shiftCnt[0], a[9]);
	and \m21_0_mux_24_18_g24/a_0(\m21_0_mux_24_18_g24/w_0, \m21_0_mux_24_18_g24/inv_sel0, a[8]);
	not \m21_0_mux_24_18_g24/i_0(\m21_0_mux_24_18_g24/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g23/org(m21_0_n_75, \m21_0_mux_24_18_g23/w_0, \m21_0_mux_24_18_g23/w_1);
	and \m21_0_mux_24_18_g23/a_1(\m21_0_mux_24_18_g23/w_1, shiftCnt[0], a[10]);
	and \m21_0_mux_24_18_g23/a_0(\m21_0_mux_24_18_g23/w_0, \m21_0_mux_24_18_g23/inv_sel0, a[9]);
	not \m21_0_mux_24_18_g23/i_0(\m21_0_mux_24_18_g23/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g22/org(m21_0_n_76, \m21_0_mux_24_18_g22/w_0, \m21_0_mux_24_18_g22/w_1);
	and \m21_0_mux_24_18_g22/a_1(\m21_0_mux_24_18_g22/w_1, shiftCnt[0], a[11]);
	and \m21_0_mux_24_18_g22/a_0(\m21_0_mux_24_18_g22/w_0, \m21_0_mux_24_18_g22/inv_sel0, a[10]);
	not \m21_0_mux_24_18_g22/i_0(\m21_0_mux_24_18_g22/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g21/org(m21_0_n_77, \m21_0_mux_24_18_g21/w_0, \m21_0_mux_24_18_g21/w_1);
	and \m21_0_mux_24_18_g21/a_1(\m21_0_mux_24_18_g21/w_1, shiftCnt[0], a[12]);
	and \m21_0_mux_24_18_g21/a_0(\m21_0_mux_24_18_g21/w_0, \m21_0_mux_24_18_g21/inv_sel0, a[11]);
	not \m21_0_mux_24_18_g21/i_0(\m21_0_mux_24_18_g21/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g20/org(m21_0_n_78, \m21_0_mux_24_18_g20/w_0, \m21_0_mux_24_18_g20/w_1);
	and \m21_0_mux_24_18_g20/a_1(\m21_0_mux_24_18_g20/w_1, shiftCnt[0], a[13]);
	and \m21_0_mux_24_18_g20/a_0(\m21_0_mux_24_18_g20/w_0, \m21_0_mux_24_18_g20/inv_sel0, a[12]);
	not \m21_0_mux_24_18_g20/i_0(\m21_0_mux_24_18_g20/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g2/org(m21_0_n_96, \m21_0_mux_24_18_g2/w_0, \m21_0_mux_24_18_g2/w_1);
	and \m21_0_mux_24_18_g2/a_1(\m21_0_mux_24_18_g2/w_1, shiftCnt[0], a[31]);
	and \m21_0_mux_24_18_g2/a_0(\m21_0_mux_24_18_g2/w_0, \m21_0_mux_24_18_g2/inv_sel0, a[30]);
	not \m21_0_mux_24_18_g2/i_0(\m21_0_mux_24_18_g2/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g19/org(m21_0_n_79, \m21_0_mux_24_18_g19/w_0, \m21_0_mux_24_18_g19/w_1);
	and \m21_0_mux_24_18_g19/a_1(\m21_0_mux_24_18_g19/w_1, shiftCnt[0], a[14]);
	and \m21_0_mux_24_18_g19/a_0(\m21_0_mux_24_18_g19/w_0, \m21_0_mux_24_18_g19/inv_sel0, a[13]);
	not \m21_0_mux_24_18_g19/i_0(\m21_0_mux_24_18_g19/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g18/org(m21_0_n_80, \m21_0_mux_24_18_g18/w_0, \m21_0_mux_24_18_g18/w_1);
	and \m21_0_mux_24_18_g18/a_1(\m21_0_mux_24_18_g18/w_1, shiftCnt[0], a[15]);
	and \m21_0_mux_24_18_g18/a_0(\m21_0_mux_24_18_g18/w_0, \m21_0_mux_24_18_g18/inv_sel0, a[14]);
	not \m21_0_mux_24_18_g18/i_0(\m21_0_mux_24_18_g18/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g17/org(m21_0_n_81, \m21_0_mux_24_18_g17/w_0, \m21_0_mux_24_18_g17/w_1);
	and \m21_0_mux_24_18_g17/a_1(\m21_0_mux_24_18_g17/w_1, shiftCnt[0], a[16]);
	and \m21_0_mux_24_18_g17/a_0(\m21_0_mux_24_18_g17/w_0, \m21_0_mux_24_18_g17/inv_sel0, a[15]);
	not \m21_0_mux_24_18_g17/i_0(\m21_0_mux_24_18_g17/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g16/org(m21_0_n_82, \m21_0_mux_24_18_g16/w_0, \m21_0_mux_24_18_g16/w_1);
	and \m21_0_mux_24_18_g16/a_1(\m21_0_mux_24_18_g16/w_1, shiftCnt[0], a[17]);
	and \m21_0_mux_24_18_g16/a_0(\m21_0_mux_24_18_g16/w_0, \m21_0_mux_24_18_g16/inv_sel0, a[16]);
	not \m21_0_mux_24_18_g16/i_0(\m21_0_mux_24_18_g16/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g15/org(m21_0_n_83, \m21_0_mux_24_18_g15/w_0, \m21_0_mux_24_18_g15/w_1);
	and \m21_0_mux_24_18_g15/a_1(\m21_0_mux_24_18_g15/w_1, shiftCnt[0], a[18]);
	and \m21_0_mux_24_18_g15/a_0(\m21_0_mux_24_18_g15/w_0, \m21_0_mux_24_18_g15/inv_sel0, a[17]);
	not \m21_0_mux_24_18_g15/i_0(\m21_0_mux_24_18_g15/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g14/org(m21_0_n_84, \m21_0_mux_24_18_g14/w_0, \m21_0_mux_24_18_g14/w_1);
	and \m21_0_mux_24_18_g14/a_1(\m21_0_mux_24_18_g14/w_1, shiftCnt[0], a[19]);
	and \m21_0_mux_24_18_g14/a_0(\m21_0_mux_24_18_g14/w_0, \m21_0_mux_24_18_g14/inv_sel0, a[18]);
	not \m21_0_mux_24_18_g14/i_0(\m21_0_mux_24_18_g14/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g13/org(m21_0_n_85, \m21_0_mux_24_18_g13/w_0, \m21_0_mux_24_18_g13/w_1);
	and \m21_0_mux_24_18_g13/a_1(\m21_0_mux_24_18_g13/w_1, shiftCnt[0], a[20]);
	and \m21_0_mux_24_18_g13/a_0(\m21_0_mux_24_18_g13/w_0, \m21_0_mux_24_18_g13/inv_sel0, a[19]);
	not \m21_0_mux_24_18_g13/i_0(\m21_0_mux_24_18_g13/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g12/org(m21_0_n_86, \m21_0_mux_24_18_g12/w_0, \m21_0_mux_24_18_g12/w_1);
	and \m21_0_mux_24_18_g12/a_1(\m21_0_mux_24_18_g12/w_1, shiftCnt[0], a[21]);
	and \m21_0_mux_24_18_g12/a_0(\m21_0_mux_24_18_g12/w_0, \m21_0_mux_24_18_g12/inv_sel0, a[20]);
	not \m21_0_mux_24_18_g12/i_0(\m21_0_mux_24_18_g12/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g11/org(m21_0_n_87, \m21_0_mux_24_18_g11/w_0, \m21_0_mux_24_18_g11/w_1);
	and \m21_0_mux_24_18_g11/a_1(\m21_0_mux_24_18_g11/w_1, shiftCnt[0], a[22]);
	and \m21_0_mux_24_18_g11/a_0(\m21_0_mux_24_18_g11/w_0, \m21_0_mux_24_18_g11/inv_sel0, a[21]);
	not \m21_0_mux_24_18_g11/i_0(\m21_0_mux_24_18_g11/inv_sel0, shiftCnt[0]);
	or \m21_0_mux_24_18_g10/org(m21_0_n_88, \m21_0_mux_24_18_g10/w_0, \m21_0_mux_24_18_g10/w_1);
	and \m21_0_mux_24_18_g10/a_1(\m21_0_mux_24_18_g10/w_1, shiftCnt[0], a[23]);
	and \m21_0_mux_24_18_g10/a_0(\m21_0_mux_24_18_g10/w_0, \m21_0_mux_24_18_g10/inv_sel0, a[22]);
	not \m21_0_mux_24_18_g10/i_0(\m21_0_mux_24_18_g10/inv_sel0, shiftCnt[0]);
	not m21_0_g1_g1(d0[31], a[31]);
	not m21_0_g1_g10(d0[22], m21_0_n_88);
	not m21_0_g1_g11(d0[21], m21_0_n_87);
	not m21_0_g1_g12(d0[20], m21_0_n_86);
	not m21_0_g1_g13(d0[19], m21_0_n_85);
	not m21_0_g1_g14(d0[18], m21_0_n_84);
	not m21_0_g1_g15(d0[17], m21_0_n_83);
	not m21_0_g1_g16(d0[16], m21_0_n_82);
	not m21_0_g1_g17(d0[15], m21_0_n_81);
	not m21_0_g1_g18(d0[14], m21_0_n_80);
	not m21_0_g1_g19(d0[13], m21_0_n_79);
	not m21_0_g1_g2(d0[30], m21_0_n_96);
	not m21_0_g1_g20(d0[12], m21_0_n_78);
	not m21_0_g1_g21(d0[11], m21_0_n_77);
	not m21_0_g1_g22(d0[10], m21_0_n_76);
	not m21_0_g1_g23(d0[9], m21_0_n_75);
	not m21_0_g1_g24(d0[8], m21_0_n_74);
	not m21_0_g1_g25(d0[7], m21_0_n_73);
	not m21_0_g1_g26(d0[6], m21_0_n_72);
	not m21_0_g1_g27(d0[5], m21_0_n_71);
	not m21_0_g1_g28(d0[4], m21_0_n_70);
	not m21_0_g1_g29(d0[3], m21_0_n_69);
	not m21_0_g1_g3(d0[29], m21_0_n_95);
	not m21_0_g1_g30(d0[2], m21_0_n_68);
	not m21_0_g1_g31(d0[1], m21_0_n_67);
	not m21_0_g1_g32(d0[0], m21_0_n_66);
	not m21_0_g1_g4(d0[28], m21_0_n_94);
	not m21_0_g1_g5(d0[27], m21_0_n_93);
	not m21_0_g1_g6(d0[26], m21_0_n_92);
	not m21_0_g1_g7(d0[25], m21_0_n_91);
	not m21_0_g1_g8(d0[24], m21_0_n_90);
	not m21_0_g1_g9(d0[23], m21_0_n_89);
	not m21_1_g1_g10(d1[22], m21_1_n_88);
	not m21_1_g1_g11(d1[21], m21_1_n_87);
	not m21_1_g1_g12(d1[20], m21_1_n_86);
	not m21_1_g1_g13(d1[19], m21_1_n_85);
	not m21_1_g1_g14(d1[18], m21_1_n_84);
	not m21_1_g1_g15(d1[17], m21_1_n_83);
	not m21_1_g1_g16(d1[16], m21_1_n_82);
	not m21_1_g1_g17(d1[15], m21_1_n_81);
	not m21_1_g1_g18(d1[14], m21_1_n_80);
	not m21_1_g1_g19(d1[13], m21_1_n_79);
	not m21_1_g1_g2(d1[30], m21_1_n_96);
	not m21_1_g1_g20(d1[12], m21_1_n_78);
	not m21_1_g1_g21(d1[11], m21_1_n_77);
	not m21_1_g1_g22(d1[10], m21_1_n_76);
	not m21_1_g1_g23(d1[9], m21_1_n_75);
	not m21_1_g1_g24(d1[8], m21_1_n_74);
	not m21_1_g1_g25(d1[7], m21_1_n_73);
	not m21_1_g1_g26(d1[6], m21_1_n_72);
	not m21_1_g1_g27(d1[5], m21_1_n_71);
	not m21_1_g1_g28(d1[4], m21_1_n_70);
	not m21_1_g1_g29(d1[3], m21_1_n_69);
	not m21_1_g1_g3(d1[29], m21_1_n_95);
	not m21_1_g1_g30(d1[2], m21_1_n_68);
	not m21_1_g1_g31(d1[1], m21_1_n_67);
	not m21_1_g1_g32(d1[0], m21_1_n_66);
	not m21_1_g1_g4(d1[28], m21_1_n_94);
	not m21_1_g1_g5(d1[27], m21_1_n_93);
	not m21_1_g1_g6(d1[26], m21_1_n_92);
	not m21_1_g1_g7(d1[25], m21_1_n_91);
	not m21_1_g1_g8(d1[24], m21_1_n_90);
	not m21_1_g1_g9(d1[23], m21_1_n_89);
	not m21_2_g1_g1(d2[31], m21_2_n_97);
	not m21_2_g1_g10(d2[22], m21_2_n_88);
	not m21_2_g1_g11(d2[21], m21_2_n_87);
	not m21_2_g1_g12(d2[20], m21_2_n_86);
	not m21_2_g1_g13(d2[19], m21_2_n_85);
	not m21_2_g1_g14(d2[18], m21_2_n_84);
	not m21_2_g1_g15(d2[17], m21_2_n_83);
	not m21_2_g1_g16(d2[16], m21_2_n_82);
	not m21_2_g1_g17(d2[15], m21_2_n_81);
	not m21_2_g1_g18(d2[14], m21_2_n_80);
	not m21_2_g1_g19(d2[13], m21_2_n_79);
	not m21_2_g1_g2(d2[30], m21_2_n_96);
	not m21_2_g1_g20(d2[12], m21_2_n_78);
	not m21_2_g1_g21(d2[11], m21_2_n_77);
	not m21_2_g1_g22(d2[10], m21_2_n_76);
	not m21_2_g1_g23(d2[9], m21_2_n_75);
	not m21_2_g1_g24(d2[8], m21_2_n_74);
	not m21_2_g1_g25(d2[7], m21_2_n_73);
	not m21_2_g1_g26(d2[6], m21_2_n_72);
	not m21_2_g1_g27(d2[5], m21_2_n_71);
	not m21_2_g1_g28(d2[4], m21_2_n_70);
	not m21_2_g1_g29(d2[3], m21_2_n_69);
	not m21_2_g1_g3(d2[29], m21_2_n_95);
	not m21_2_g1_g30(d2[2], m21_2_n_68);
	not m21_2_g1_g31(d2[1], m21_2_n_67);
	not m21_2_g1_g32(d2[0], m21_2_n_66);
	not m21_2_g1_g4(d2[28], m21_2_n_94);
	not m21_2_g1_g5(d2[27], m21_2_n_93);
	not m21_2_g1_g6(d2[26], m21_2_n_92);
	not m21_2_g1_g7(d2[25], m21_2_n_91);
	not m21_2_g1_g8(d2[24], m21_2_n_90);
	not m21_2_g1_g9(d2[23], m21_2_n_89);
	not m21_3_g1_g1(d3[31], n_136);
	not m21_3_g1_g10(d3[22], m21_3_n_88);
	not m21_3_g1_g11(d3[21], m21_3_n_87);
	not m21_3_g1_g12(d3[20], m21_3_n_86);
	not m21_3_g1_g13(d3[19], m21_3_n_85);
	not m21_3_g1_g14(d3[18], m21_3_n_84);
	not m21_3_g1_g15(d3[17], m21_3_n_83);
	not m21_3_g1_g16(d3[16], m21_3_n_82);
	not m21_3_g1_g17(d3[15], m21_3_n_81);
	not m21_3_g1_g18(d3[14], m21_3_n_80);
	not m21_3_g1_g19(d3[13], m21_3_n_79);
	not m21_3_g1_g2(d3[30], n_140);
	not m21_3_g1_g20(d3[12], m21_3_n_78);
	not m21_3_g1_g21(d3[11], m21_3_n_77);
	not m21_3_g1_g22(d3[10], m21_3_n_76);
	not m21_3_g1_g23(d3[9], m21_3_n_75);
	not m21_3_g1_g24(d3[8], m21_3_n_74);
	not m21_3_g1_g25(d3[7], m21_3_n_73);
	not m21_3_g1_g26(d3[6], m21_3_n_72);
	not m21_3_g1_g27(d3[5], m21_3_n_71);
	not m21_3_g1_g28(d3[4], m21_3_n_70);
	not m21_3_g1_g29(d3[3], m21_3_n_69);
	not m21_3_g1_g3(d3[29], n_144);
	not m21_3_g1_g30(d3[2], m21_3_n_68);
	not m21_3_g1_g31(d3[1], m21_3_n_67);
	not m21_3_g1_g32(d3[0], m21_3_n_66);
	not m21_3_g1_g4(d3[28], n_148);
	not m21_3_g1_g5(d3[27], n_152);
	not m21_3_g1_g6(d3[26], n_156);
	not m21_3_g1_g7(d3[25], n_160);
	not m21_3_g1_g8(d3[24], n_164);
	not m21_3_g1_g9(d3[23], m21_3_n_89);
	not m21_4_g1_g1(z[31], n_168);
	not m21_4_g1_g10(z[22], n_172);
	not m21_4_g1_g11(sub_wire0, n_176);
	not m21_4_g1_g12(z[20], n_180);
	not m21_4_g1_g13(z[19], n_184);
	not m21_4_g1_g14(z[18], n_188);
	not m21_4_g1_g15(z[17], n_192);
	not m21_4_g1_g16(z[16], n_196);
	not m21_4_g1_g17(z[15], m21_4_n_81);
	not m21_4_g1_g18(z[14], m21_4_n_80);
	not m21_4_g1_g19(z[13], m21_4_n_79);
	not m21_4_g1_g2(z[30], n_200);
	not m21_4_g1_g20(z[12], m21_4_n_78);
	not m21_4_g1_g21(z[11], m21_4_n_77);
	not m21_4_g1_g22(z[10], m21_4_n_76);
	not m21_4_g1_g23(z[9], m21_4_n_75);
	not m21_4_g1_g24(z[8], m21_4_n_74);
	not m21_4_g1_g25(z[7], m21_4_n_73);
	not m21_4_g1_g26(z[6], m21_4_n_72);
	not m21_4_g1_g27(z[5], m21_4_n_71);
	not m21_4_g1_g28(z[4], m21_4_n_70);
	not m21_4_g1_g29(z[3], m21_4_n_69);
	not m21_4_g1_g3(z[29], n_204);
	not m21_4_g1_g30(z[2], m21_4_n_68);
	not m21_4_g1_g31(z[1], m21_4_n_67);
	not m21_4_g1_g32(z[0], m21_4_n_66);
	not m21_4_g1_g4(z[28], n_208);
	not m21_4_g1_g5(z[27], n_212);
	not m21_4_g1_g6(z[26], n_216);
	not m21_4_g1_g7(z[25], n_220);
	not m21_4_g1_g8(z[24], n_224);
	not m21_4_g1_g9(z[23], n_228);
	xor g34(d1[31], a[31], shiftCnt[1]);
	and g35(n_134, shiftCnt[3], a[31]);
	not g36(n_133, shiftCnt[3]);
	and g37(n_135, n_133, d2[31]);
	or g38(n_136, n_134, n_135);
	and g41(n_139, n_133, d2[30]);
	or g42(n_140, n_134, n_139);
	and g45(n_143, n_133, d2[29]);
	or g46(n_144, n_134, n_143);
	and g49(n_147, n_133, d2[28]);
	or g50(n_148, n_134, n_147);
	and g53(n_151, n_133, d2[27]);
	or g54(n_152, n_134, n_151);
	and g57(n_155, n_133, d2[26]);
	or g58(n_156, n_134, n_155);
	and g61(n_159, n_133, d2[25]);
	or g62(n_160, n_134, n_159);
	and g65(n_163, n_133, d2[24]);
	or g66(n_164, n_134, n_163);
	and g67(n_166, shiftCnt[4], a[31]);
	not g68(n_165, shiftCnt[4]);
	and g69(n_167, n_165, d3[31]);
	or g70(n_168, n_166, n_167);
	and g73(n_171, n_165, d3[22]);
	or g74(n_172, n_166, n_171);
	and g77(n_175, n_165, d3[21]);
	or g78(n_176, n_166, n_175);
	and g81(n_179, n_165, d3[20]);
	or g82(n_180, n_166, n_179);
	and g85(n_183, n_165, d3[19]);
	or g86(n_184, n_166, n_183);
	and g89(n_187, n_165, d3[18]);
	or g90(n_188, n_166, n_187);
	and g93(n_191, n_165, d3[17]);
	or g94(n_192, n_166, n_191);
	and g97(n_195, n_165, d3[16]);
	or g98(n_196, n_166, n_195);
	and g101(n_199, n_165, d3[30]);
	or g102(n_200, n_166, n_199);
	and g105(n_203, n_165, d3[29]);
	or g106(n_204, n_166, n_203);
	and g109(n_207, n_165, d3[28]);
	or g110(n_208, n_166, n_207);
	and g113(n_211, n_165, d3[27]);
	or g114(n_212, n_166, n_211);
	and g117(n_215, n_165, d3[26]);
	or g118(n_216, n_166, n_215);
	and g121(n_219, n_165, d3[25]);
	or g122(n_220, n_166, n_219);
	and g125(n_223, n_165, d3[24]);
	or g126(n_224, n_166, n_223);
	and g129(n_227, n_165, d3[23]);
	or g130(n_228, n_166, n_227);
	assign w_eco0 = !shiftCnt[4];
	assign w_eco1 = !a[31];
	or _ECO_2(w_eco2, w_eco0, w_eco1);
	xor _ECO_out0(z[21], sub_wire0, w_eco2);

endmodule