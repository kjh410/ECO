module top(parity,overflow,greater,is_eq,less,y,a,b,op);
	input [7:0]a, b;
	input [1:0]op;
	output parity, overflow, greater, is_eq, less;
	output [7:0]y;
	wire \mux_44_12_g156/w_0, \mux_44_12_g156/w_1, \mux_44_12_g156/w_2, \mux_temp_y_21_12_g792/w_0, \mux_temp_y_21_12_g792/w_1, \mux_temp_y_21_12_g19/w_0, \mux_temp_y_21_12_g19/w_1, \mux_temp_y_21_12_g19/w_2, \mux_temp_y_21_12_g19/w_3, \mux_temp_y_21_12_g18/w_0, \mux_temp_y_21_12_g18/w_1, \mux_temp_y_21_12_g18/w_2, \mux_temp_y_21_12_g18/w_3, \mux_temp_y_21_12_g17/w_0, \mux_temp_y_21_12_g17/w_1, \mux_temp_y_21_12_g17/w_2, \mux_temp_y_21_12_g17/w_3, \mux_temp_y_21_12_g16/w_0, \mux_temp_y_21_12_g16/w_1, \mux_temp_y_21_12_g16/w_2, \mux_temp_y_21_12_g16/w_3, \mux_temp_y_21_12_g15/w_0, \mux_temp_y_21_12_g15/w_1, \mux_temp_y_21_12_g15/w_2, \mux_temp_y_21_12_g15/w_3, \mux_temp_y_21_12_g10/w_0, \mux_temp_y_21_12_g10/w_1, \mux_temp_y_21_12_g10/w_2, \mux_temp_y_21_12_g10/w_3, sub_29_29_n_1105, sub_29_29_n_1103, sub_29_29_n_320, sub_29_29_n_69, sub_29_29_n_66, sub_29_29_n_63, sub_29_29_n_59, sub_29_29_n_54, sub_29_29_n_37, sub_29_29_n_32, n_1123, n_1114, n_1113, n_1112, n_1111, n_1106, n_1104, n_1102, n_1101, n_1099, n_1098, n_1097, n_1096, n_1095, n_988, n_987, n_986, n_985, n_984, n_983, n_982, n_981, n_980, n_979, n_978, n_977, n_976, n_975, n_974, n_973, n_972, n_971, n_970, n_969, n_968, n_967, n_966, n_965, n_964, n_963, n_962, n_961, n_960, n_959, n_958, n_957, n_956, n_955, n_954, n_953, n_952, n_951, n_950, n_949, n_948, n_947, n_946, n_945, n_944, n_943, n_942, n_940, n_939, n_938, n_937, n_936, n_935, n_934, n_933, n_932, n_931, n_930, n_929, n_928, n_927, n_926, n_925, n_924, n_923, n_922, n_921, n_920, n_919, n_918, n_917, n_916, n_915, n_914, n_913, n_912, n_911, n_910, n_909, n_908, n_907, n_906, n_905, n_904, n_903, n_902, n_901, n_900, n_898, n_897, n_895, n_894, n_892, n_891, n_890, n_889, n_888, n_887, n_886, n_885, n_884, n_883, n_882, n_881, n_880, n_878, n_877, n_876, n_875, n_874, n_873, n_872, n_871, n_870, n_869, n_867, n_866, n_865, n_864, n_863, n_862, n_861, n_860, n_859, n_858, n_857, n_856, n_840, n_827, n_806, n_805, n_620, n_619, n_618, n_617, n_616, n_615, n_437, n_436, n_435, n_431, n_429, n_428, n_419, n_416, n_415, n_397, n_395, n_379, n_367, n_323, n_318, n_308, n_301, n_300, n_298, n_136, n_135, n_133, n_132, n_131, n_130, n_129, n_77, n_76, n_75, n_74, n_73, n_43, n_41, n_39, n_38, n_37, n_35, n_34, n_33, n_31, n_30, n_29, n_26, n_25, n_23, n_22, n_21, n_19, n_18, n_17, n_16, gt_39_12_n_57, gt_39_12_n_52, gt_39_12_n_46, gt_25_24_n_35, add_24_29_n_1115, add_24_29_n_57, add_24_29_n_55, add_24_29_n_53, add_24_29_n_51, add_24_29_n_50, add_24_29_n_49, add_24_29_n_48, add_24_29_n_47, add_24_29_n_43, add_24_29_n_39, add_24_29_n_37, add_24_29_n_33, add_24_29_n_27, less, is_eq, greater, overflow, parity, \mux_44_12_g156/data0;
	wire [7:0]y;
	wire [1:0]op;
	wire [7:0]b, a;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388;

	assign \mux_44_12_g156/data0 = 0;
	or \mux_44_12_g156/org(sub_wire0, \mux_44_12_g156/w_0, \mux_44_12_g156/w_1, \mux_44_12_g156/w_2);
	and \mux_44_12_g156/a_2(\mux_44_12_g156/w_2, n_988, n_43);
	and \mux_44_12_g156/a_1(\mux_44_12_g156/w_1, n_987, n_41);
	and \mux_44_12_g156/a_0(\mux_44_12_g156/w_0, n_986, n_43);
	or \mux_temp_y_21_12_g792/org(n_129, \mux_temp_y_21_12_g792/w_0, \mux_temp_y_21_12_g792/w_1);
	and \mux_temp_y_21_12_g792/a_1(\mux_temp_y_21_12_g792/w_1, n_805, n_16);
	and \mux_temp_y_21_12_g792/a_0(\mux_temp_y_21_12_g792/w_0, n_318, n_1114);
	or \mux_temp_y_21_12_g19/org(n_136, \mux_temp_y_21_12_g19/w_0, \mux_temp_y_21_12_g19/w_1, \mux_temp_y_21_12_g19/w_2, \mux_temp_y_21_12_g19/w_3);
	and \mux_temp_y_21_12_g19/a_3(\mux_temp_y_21_12_g19/w_3, n_301, n_616);
	and \mux_temp_y_21_12_g19/a_2(\mux_temp_y_21_12_g19/w_2, n_318, n_35);
	and \mux_temp_y_21_12_g19/a_1(\mux_temp_y_21_12_g19/w_1, n_1095, n_34);
	and \mux_temp_y_21_12_g19/a_0(\mux_temp_y_21_12_g19/w_0, n_1111, n_33);
	or \mux_temp_y_21_12_g18/org(n_135, \mux_temp_y_21_12_g18/w_0, \mux_temp_y_21_12_g18/w_1, \mux_temp_y_21_12_g18/w_2, \mux_temp_y_21_12_g18/w_3);
	and \mux_temp_y_21_12_g18/a_3(\mux_temp_y_21_12_g18/w_3, n_301, n_615);
	and \mux_temp_y_21_12_g18/a_2(\mux_temp_y_21_12_g18/w_2, n_318, n_39);
	and \mux_temp_y_21_12_g18/a_1(\mux_temp_y_21_12_g18/w_1, n_1095, n_38);
	and \mux_temp_y_21_12_g18/a_0(\mux_temp_y_21_12_g18/w_0, n_1111, n_37);
	or \mux_temp_y_21_12_g17/org(n_133, \mux_temp_y_21_12_g17/w_0, \mux_temp_y_21_12_g17/w_1, \mux_temp_y_21_12_g17/w_2, \mux_temp_y_21_12_g17/w_3);
	and \mux_temp_y_21_12_g17/a_3(\mux_temp_y_21_12_g17/w_3, n_301, n_620);
	and \mux_temp_y_21_12_g17/a_2(\mux_temp_y_21_12_g17/w_2, n_318, n_1113);
	and \mux_temp_y_21_12_g17/a_1(\mux_temp_y_21_12_g17/w_1, n_1095, n_26);
	and \mux_temp_y_21_12_g17/a_0(\mux_temp_y_21_12_g17/w_0, n_1111, n_25);
	or \mux_temp_y_21_12_g16/org(n_132, \mux_temp_y_21_12_g16/w_0, \mux_temp_y_21_12_g16/w_1, \mux_temp_y_21_12_g16/w_2, \mux_temp_y_21_12_g16/w_3);
	and \mux_temp_y_21_12_g16/a_3(\mux_temp_y_21_12_g16/w_3, n_301, n_619);
	and \mux_temp_y_21_12_g16/a_2(\mux_temp_y_21_12_g16/w_2, n_318, n_31);
	and \mux_temp_y_21_12_g16/a_1(\mux_temp_y_21_12_g16/w_1, n_1095, n_30);
	and \mux_temp_y_21_12_g16/a_0(\mux_temp_y_21_12_g16/w_0, n_1111, n_29);
	or \mux_temp_y_21_12_g15/org(n_131, \mux_temp_y_21_12_g15/w_0, \mux_temp_y_21_12_g15/w_1, \mux_temp_y_21_12_g15/w_2, \mux_temp_y_21_12_g15/w_3);
	and \mux_temp_y_21_12_g15/a_3(\mux_temp_y_21_12_g15/w_3, n_301, n_618);
	and \mux_temp_y_21_12_g15/a_2(\mux_temp_y_21_12_g15/w_2, n_318, n_23);
	and \mux_temp_y_21_12_g15/a_1(\mux_temp_y_21_12_g15/w_1, n_1095, n_22);
	and \mux_temp_y_21_12_g15/a_0(\mux_temp_y_21_12_g15/w_0, n_1111, n_21);
	or \mux_temp_y_21_12_g10/org(n_130, \mux_temp_y_21_12_g10/w_0, \mux_temp_y_21_12_g10/w_1, \mux_temp_y_21_12_g10/w_2, \mux_temp_y_21_12_g10/w_3);
	and \mux_temp_y_21_12_g10/a_3(\mux_temp_y_21_12_g10/w_3, n_301, n_617);
	and \mux_temp_y_21_12_g10/a_2(\mux_temp_y_21_12_g10/w_2, n_318, n_19);
	and \mux_temp_y_21_12_g10/a_1(\mux_temp_y_21_12_g10/w_1, n_1095, n_18);
	and \mux_temp_y_21_12_g10/a_0(\mux_temp_y_21_12_g10/w_0, n_1111, n_17);
	nor add_24_29_g10(add_24_29_n_33, a[3], b[3]);
	nor add_24_29_g12(add_24_29_n_43, a[4], b[4]);
	nor add_24_29_g14(add_24_29_n_39, a[5], b[5]);
	nor add_24_29_g16(add_24_29_n_50, a[6], b[6]);
	nor add_24_29_g23(add_24_29_n_48, n_880, n_1113);
	nor add_24_29_g24(add_24_29_n_47, add_24_29_n_37, add_24_29_n_33);
	nor add_24_29_g27(add_24_29_n_51, n_884, n_35);
	nor add_24_29_g28(add_24_29_n_55, add_24_29_n_43, add_24_29_n_39);
	nand add_24_29_g32(add_24_29_n_49, add_24_29_n_47, add_24_29_n_1115);
	nand add_24_29_g33(add_24_29_n_57, add_24_29_n_48, add_24_29_n_49);
	nor add_24_29_g34(add_24_29_n_53, add_24_29_n_50, add_24_29_n_51);
	xnor add_24_29_g48(n_17, n_1114, n_965);
	xnor add_24_29_g50(n_21, add_24_29_n_1115, n_966);
	xnor add_24_29_g53(n_25, n_972, n_970);
	xnor add_24_29_g55(n_29, add_24_29_n_57, n_969);
	xnor add_24_29_g58(n_33, n_979, n_968);
	nor add_24_29_g6(add_24_29_n_27, a[1], b[1]);
	xnor add_24_29_g60(n_37, n_978, n_967);
	nor add_24_29_g8(add_24_29_n_37, a[2], b[2]);
	xor g15(n_16, a[0], b[0]);
	xor g21(n_74, n_129, n_135);
	xor g22(n_75, n_136, n_130);
	xor g23(n_76, n_131, n_73);
	xor g24(n_77, n_74, n_75);
	xor g25(parity, n_76, n_77);
	xor g3(n_73, n_132, n_133);
	not gt_39_12_g10(greater, n_840);
	nand sub_29_29_g38(sub_29_29_n_54, sub_29_29_n_320, n_1104);
	nand sub_29_29_g46(sub_29_29_n_69, sub_29_29_n_63, n_300);
	xnor sub_29_29_g56(n_18, sub_29_29_n_37, n_617);
	xnor sub_29_29_g58(n_22, sub_29_29_n_320, n_618);
	xnor sub_29_29_g61(n_26, n_977, n_620);
	xnor sub_29_29_g63(n_30, sub_29_29_n_1105, n_619);
	xnor sub_29_29_g66(n_34, n_985, n_616);
	xnor sub_29_29_g68(n_38, n_984, n_615);
	not sub_29_29_g9(n_43, sub_29_29_n_32);
	nor g251(n_395, n_916, n_1096, gt_39_12_n_57);
	nor g287(n_419, n_1102, a[0]);
	nor g298(n_429, n_1096, gt_39_12_n_57, n_397);
	nor g299(n_428, gt_39_12_n_57, n_323, n_397);
	nor g303(n_431, n_1104, gt_39_12_n_46);
	not g793(n_805, n_318);
	not g904(n_872, a[7]);
	not g907(n_875, add_24_29_n_33);
	not g915(n_881, n_1113);
	not g916(n_882, add_24_29_n_37);
	not g931(n_891, gt_39_12_n_52);
	not g933(n_892, n_308);
	nor g936(gt_39_12_n_57, n_872, b[7]);
	not g937(n_894, gt_39_12_n_57);
	nand g938(n_895, n_891, n_892, n_1097, n_894);
	not g942(n_897, n_431);
	not g949(n_901, n_419);
	nor g952(n_903, n_1102, n_871);
	not g953(n_904, n_903);
	nand g954(n_905, n_901, sub_29_29_n_1103, n_904);
	nand g955(n_906, n_1098, n_1101, n_905);
	nand g956(n_907, n_897, n_1099, n_906);
	not g957(n_908, n_907);
	nor g958(n_909, n_895, n_908);
	not g959(n_910, n_909);
	not g965(n_913, sub_29_29_n_63);
	nor g966(n_914, n_891, n_911);
	not g967(n_915, n_914);
	nand g968(n_916, n_913, n_915);
	nand g971(n_323, n_872, b[7]);
	not g972(n_918, n_323);
	nor g973(n_919, n_395, n_917, n_918);
	not g974(n_920, n_919);
	nor g975(n_921, n_395, n_894, n_918);
	not g976(n_922, n_921);
	nand g977(n_923, n_920, n_922);
	nand g978(n_840, n_910, n_923);
	not g985(n_928, sub_29_29_n_69);
	nor g992(n_397, n_918, n_932);
	not g993(n_933, n_429);
	not g994(n_934, n_428);
	nand g995(n_367, n_933, n_934);
	not g996(n_935, n_367);
	nor g997(n_936, greater, n_367);
	not g998(n_937, n_936);
	nand g1004(n_379, n_928, n_323, sub_29_29_n_1105);
	not g1005(n_942, n_379);
	nor g1006(n_943, greater, n_379);
	not g1007(n_944, n_943);
	nand g1008(is_eq, n_937, n_944);
	nor g1009(less, greater, n_935, n_942);
	nor g1036(n_318, n_1123, op[0]);
	nor g1037(n_301, n_1123, n_869);
	nand g1038(n_965, n_888, n_887);
	nand g1039(n_966, n_882, n_1112);
	nand g1041(n_615, n_300, n_1097);
	nand g1043(n_616, n_891, n_298);
	nand g1044(n_617, n_900, sub_29_29_n_1103);
	nand g1045(n_618, n_1101, n_1104);
	nand g1047(n_619, n_892, sub_29_29_n_66);
	nand g1048(n_970, n_875, n_881);
	nand g1049(n_620, n_1098, n_1099);
	nand g1050(n_971, n_882, add_24_29_n_1115);
	nand g1051(n_972, n_1112, n_971);
	nand g1056(n_977, sub_29_29_n_54, n_1101);
	nor g1059(n_980, n_913, n_1106);
	not g1060(n_981, n_980);
	nor g1061(n_982, n_912, n_1106);
	not g1062(n_983, n_982);
	nand g1063(n_984, sub_29_29_n_59, n_981);
	nand g1064(n_985, n_892, n_983);
	not g901(n_869, op[0]);
	nor g1029(n_1095, op[1], n_869);
	not g1030(n_960, n_1095);
	not g895(n_863, a[6]);
	nor g934(n_1096, n_863, b[6]);
	not g935(n_1097, n_1096);
	nand g969(n_300, n_863, b[6]);
	not g970(n_917, n_300);
	not g893(n_861, a[5]);
	nor g930(gt_39_12_n_52, n_861, b[5]);
	nand g960(n_298, n_861, b[5]);
	nor g282(n_416, gt_39_12_n_52, n_298);
	not g987(n_930, n_416);
	not g891(n_859, a[4]);
	nor g932(n_308, n_859, b[4]);
	nor g283(n_415, gt_39_12_n_52, n_308);
	not g988(n_931, n_415);
	nand g989(sub_29_29_n_59, n_930, n_931);
	nor g990(n_827, n_917, sub_29_29_n_59);
	not g991(n_932, n_827);
	not g961(n_911, n_298);
	nand g962(sub_29_29_n_66, n_859, b[4]);
	not g963(n_912, sub_29_29_n_66);
	nor g964(sub_29_29_n_63, n_911, n_912);
	not g889(n_857, a[3]);
	nor g940(gt_39_12_n_46, n_857, b[3]);
	not g941(n_1098, gt_39_12_n_46);
	nand g943(n_1099, n_857, b[3]);
	not g944(n_898, n_1099);
	not g899(n_867, a[2]);
	nor g945(n_806, n_867, b[2]);
	not g946(n_1101, n_806);
	nor g999(n_938, n_898, n_1101);
	not g1000(n_939, n_938);
	not g897(n_865, a[1]);
	nor g947(n_1102, n_865, b[1]);
	not g948(n_900, n_1102);
	nand g950(sub_29_29_n_1103, n_865, b[1]);
	not g951(n_902, sub_29_29_n_1103);
	not g902(n_870, a[0]);
	nand g979(sub_29_29_n_37, n_870, b[0]);
	not g980(n_924, sub_29_29_n_37);
	nor g981(n_925, n_902, n_924);
	not g982(n_926, n_925);
	nand g983(sub_29_29_n_320, n_900, n_926);
	nand g939(n_1104, n_867, b[2]);
	not g984(n_927, sub_29_29_n_54);
	nand g1001(n_940, n_927, n_1099);
	nand g1002(sub_29_29_n_1105, n_1098, n_939, n_940);
	not g1003(n_1106, sub_29_29_n_1105);
	nor g1010(n_945, sub_29_29_n_69, n_1106);
	not g1011(n_946, n_945);
	nand g1012(sub_29_29_n_32, n_1097, n_932, n_946);
	nor g1031(n_961, n_960, sub_29_29_n_32);
	not g1032(n_962, n_961);
	nor g108(n_1111, op[0], op[1]);
	not g986(n_929, n_1111);
	not g890(n_858, b[4]);
	nor g917(n_31, n_859, n_858);
	not g918(n_883, n_31);
	nor g919(n_884, add_24_29_n_39, n_883);
	not g892(n_860, b[5]);
	nor g920(n_35, n_861, n_860);
	not g922(n_886, add_24_29_n_55);
	not g898(n_866, b[2]);
	nor g911(n_23, n_867, n_866);
	not g912(n_1112, n_23);
	nor g913(n_880, add_24_29_n_33, n_1112);
	not g888(n_856, b[3]);
	nor g914(n_1113, n_857, n_856);
	not g896(n_864, b[1]);
	nor g923(n_19, n_865, n_864);
	not g924(n_887, n_19);
	not g925(n_888, add_24_29_n_27);
	not g903(n_871, b[0]);
	nor g926(n_1114, n_870, n_871);
	nand g927(n_889, n_888, n_1114);
	nand g928(add_24_29_n_1115, n_887, n_889);
	not g1013(n_947, add_24_29_n_57);
	nor g1052(n_973, n_886, n_947);
	not g1053(n_974, n_973);
	nand g1057(n_978, add_24_29_n_51, n_974);
	not g910(n_878, add_24_29_n_50);
	not g894(n_862, b[6]);
	nor g1014(n_39, n_863, n_862);
	not g1015(n_948, n_39);
	nand g1040(n_967, n_878, n_948);
	not g905(n_873, n_37);
	not g908(n_876, add_24_29_n_43);
	nand g1046(n_969, n_876, n_883);
	not g929(n_890, add_24_29_n_53);
	nand g1016(n_949, n_878, add_24_29_n_55);
	nor g1017(n_950, n_947, n_949);
	not g1018(n_951, n_950);
	nand g1019(n_41, n_890, n_948, n_951);
	nor g307(n_436, n_29, n_41);
	not g1021(n_953, n_436);
	nor g1054(n_975, add_24_29_n_43, n_947);
	not g1055(n_976, n_975);
	nand g1058(n_979, n_883, n_976);
	not g909(n_877, add_24_29_n_39);
	not g921(n_885, n_35);
	nand g1042(n_968, n_877, n_885);
	nor g308(n_435, n_33, n_41);
	not g1022(n_954, n_435);
	nand g1023(n_437, n_953, n_954);
	nor g1024(n_955, n_873, n_437);
	not g1025(n_956, n_955);
	not g1020(n_952, n_41);
	nor g1026(n_957, n_952, n_437);
	not g1027(n_958, n_957);
	nand g1028(n_959, n_956, n_958);
	nand g498(gt_25_24_n_35, n_959, n_41);
	nor g1033(n_963, n_929, gt_25_24_n_35);
	not g1034(n_964, n_963);
	nand g1035(overflow, n_962, n_964);
	not g900(n_1123, op[1]);
	nand g1065(n_986, overflow, n_1123);
	not g906(n_874, overflow);
	nor g1066(n_987, n_874, n_929);
	nor g1067(n_988, n_874, n_960);
	and g1068(y[6], overflow, n_135);
	and g1069(y[5], overflow, n_136);
	and g1070(y[4], overflow, n_132);
	and g1071(y[3], overflow, n_133);
	and g1072(y[2], overflow, n_131);
	and g1073(y[1], overflow, n_130);
	and g1074(y[0], overflow, n_129);
	and _ECO_0(w_eco0, !a[4], !b[4], a[5], b[5], b[6]);
	and _ECO_1(w_eco1, !a[4], !b[4], !a[5], a[6], b[6]);
	and _ECO_2(w_eco2, !a[4], !a[5], !a[6], op[0]);
	and _ECO_3(w_eco3, b[4], !a[5], !b[5], a[6], b[6]);
	and _ECO_4(w_eco4, b[4], b[5], b[6], op[0]);
	and _ECO_5(w_eco5, b[4], b[5], !a[6], op[0]);
	and _ECO_6(w_eco6, !a[4], b[5], !a[6], op[0]);
	and _ECO_7(w_eco7, !a[6], b[6], op[0]);
	and _ECO_8(w_eco8, !a[5], b[5], !a[6], op[0]);
	and _ECO_9(w_eco9, !a[4], !a[5], !a[6], op[1]);
	and _ECO_10(w_eco10, b[4], !a[5], !a[6], op[0]);
	and _ECO_11(w_eco11, b[4], b[5], b[6], op[1]);
	and _ECO_12(w_eco12, b[4], b[5], !a[6], op[1]);
	and _ECO_13(w_eco13, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[2]);
	and _ECO_14(w_eco14, !a[4], b[5], !a[6], op[1]);
	and _ECO_15(w_eco15, !a[5], b[5], b[6], op[0]);
	and _ECO_16(w_eco16, !a[6], b[6], op[1]);
	and _ECO_17(w_eco17, !a[5], b[5], !a[6], op[1]);
	and _ECO_18(w_eco18, !a[3], a[4], a[5], !a[2], op[0]);
	and _ECO_19(w_eco19, !a[3], !a[4], !b[4], a[6], b[6], !a[2]);
	and _ECO_20(w_eco20, !a[3], !b[4], a[5], !a[2], op[0]);
	and _ECO_21(w_eco21, b[4], !a[5], !a[6], op[1]);
	and _ECO_22(w_eco22, !a[3], !a[5], !b[5], a[6], b[6], !a[2]);
	and _ECO_23(w_eco23, !a[3], a[4], !b[5], !a[2], op[0]);
	and _ECO_24(w_eco24, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6]);
	and _ECO_25(w_eco25, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2]);
	and _ECO_26(w_eco26, !a[5], b[5], b[6], op[1]);
	and _ECO_27(w_eco27, !a[3], b[3], a[4], a[5], op[0]);
	and _ECO_28(w_eco28, b[3], a[4], a[5], !a[2], op[0]);
	and _ECO_29(w_eco29, !a[3], a[4], a[5], !a[2], op[1]);
	and _ECO_30(w_eco30, !a[3], b[3], !a[4], !b[4], a[6], b[6]);
	and _ECO_31(w_eco31, b[3], !a[4], !b[4], a[6], b[6], !a[2]);
	and _ECO_32(w_eco32, !a[3], b[3], !b[4], a[5], op[0]);
	and _ECO_33(w_eco33, b[3], !b[4], a[5], !a[2], op[0]);
	and _ECO_34(w_eco34, !a[3], !b[4], a[5], !a[2], op[1]);
	and _ECO_35(w_eco35, !a[3], b[3], !a[5], !b[5], a[6], b[6]);
	and _ECO_36(w_eco36, b[3], !a[5], !b[5], a[6], b[6], !a[2]);
	and _ECO_37(w_eco37, !a[3], b[3], a[4], !b[5], op[0]);
	and _ECO_38(w_eco38, b[3], a[4], !b[5], !a[2], op[0]);
	and _ECO_39(w_eco39, !a[3], a[4], !b[5], !a[2], op[1]);
	and _ECO_40(w_eco40, !a[3], !b[4], !b[5], !a[2], op[0]);
	and _ECO_41(w_eco41, !a[3], !b[3], a[4], b[4], b[5], b[6]);
	and _ECO_42(w_eco42, !a[3], !b[3], !a[4], a[5], b[5], b[6]);
	and _ECO_43(w_eco43, !a[3], b[3], a[4], a[5], op[1]);
	and _ECO_44(w_eco44, b[3], a[4], a[5], !a[2], op[1]);
	and _ECO_45(w_eco45, !a[3], b[3], !b[4], a[5], op[1]);
	and _ECO_46(w_eco46, b[3], !b[4], a[5], !a[2], op[1]);
	and _ECO_47(w_eco47, !a[3], b[3], a[4], !b[5], op[1]);
	and _ECO_48(w_eco48, b[3], a[4], !b[5], !a[2], op[1]);
	and _ECO_49(w_eco49, !a[3], b[3], !b[4], !b[5], op[0]);
	and _ECO_50(w_eco50, b[3], !b[4], !b[5], !a[2], op[0]);
	and _ECO_51(w_eco51, !a[3], !b[4], !b[5], !a[2], op[1]);
	and _ECO_52(w_eco52, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[2]);
	and _ECO_53(w_eco53, !a[3], !b[3], a[4], a[6], b[6], !a[2]);
	and _ECO_54(w_eco54, !a[3], !b[3], a[5], b[5], !a[6], b[6]);
	and _ECO_55(w_eco55, !a[3], !b[3], a[4], a[5], b[5], a[6], !a[2]);
	and _ECO_56(w_eco56, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[0]);
	and _ECO_57(w_eco57, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[0]);
	and _ECO_58(w_eco58, !a[3], !b[3], !a[4], !a[5], a[6], b[6]);
	and _ECO_59(w_eco59, !a[3], !b[3], !a[5], b[5], a[6], b[6]);
	and _ECO_60(w_eco60, !a[3], !b[3], a[4], b[4], a[5], !a[6], b[6]);
	and _ECO_61(w_eco61, b[3], a[4], a[5], !b[1], !b[0], op[0]);
	and _ECO_62(w_eco62, a[4], a[5], !b[1], a[2], !b[0], op[0]);
	and _ECO_63(w_eco63, b[3], !a[4], !b[4], a[6], b[6], !b[1], !b[0]);
	and _ECO_64(w_eco64, !a[4], !b[4], a[6], b[6], !b[1], a[2], !b[0]);
	and _ECO_65(w_eco65, b[3], !b[4], a[5], !b[1], !b[0], op[0]);
	and _ECO_66(w_eco66, !b[4], a[5], !b[1], a[2], !b[0], op[0]);
	and _ECO_67(w_eco67, b[3], !a[5], !b[5], a[6], b[6], !b[1], !b[0]);
	and _ECO_68(w_eco68, !a[5], !b[5], a[6], b[6], !b[1], a[2], !b[0]);
	and _ECO_69(w_eco69, b[3], a[4], !b[5], !b[1], !b[0], op[0]);
	and _ECO_70(w_eco70, a[4], !b[5], !b[1], a[2], !b[0], op[0]);
	and _ECO_71(w_eco71, !a[3], b[3], !b[4], !b[5], op[1]);
	and _ECO_72(w_eco72, b[3], !b[4], !b[5], !a[2], op[1]);
	and _ECO_73(w_eco73, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0]);
	and _ECO_74(w_eco74, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0]);
	and _ECO_75(w_eco75, !b[3], !a[4], a[5], b[5], b[6], !b[1], !a[2], !b[0]);
	and _ECO_76(w_eco76, !a[3], a[5], b[5], b[6], !b[1], !a[2], !b[0]);
	and _ECO_77(w_eco77, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[0]);
	and _ECO_78(w_eco78, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[0]);
	and _ECO_79(w_eco79, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], a[0]);
	and _ECO_80(w_eco80, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[0]);
	and _ECO_81(w_eco81, !b[3], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0]);
	and _ECO_82(w_eco82, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0]);
	and _ECO_83(w_eco83, b[3], a[4], a[5], !b[1], a[0], op[0]);
	and _ECO_84(w_eco84, b[3], a[4], a[5], a[1], !b[0], op[0]);
	and _ECO_85(w_eco85, a[4], a[5], !b[1], a[2], a[0], op[0]);
	and _ECO_86(w_eco86, a[4], a[5], a[1], a[2], !b[0], op[0]);
	and _ECO_87(w_eco87, b[3], a[4], a[5], !b[1], !b[0], op[1]);
	and _ECO_88(w_eco88, a[4], a[5], !b[1], a[2], !b[0], op[1]);
	and _ECO_89(w_eco89, a[4], a[5], !b[1], !b[2], !b[0], op[0]);
	and _ECO_90(w_eco90, b[3], !a[4], !b[4], a[6], b[6], !b[1], a[0]);
	and _ECO_91(w_eco91, b[3], !a[4], !b[4], a[6], b[6], a[1], !b[0]);
	and _ECO_92(w_eco92, !a[4], !b[4], a[6], b[6], !b[1], a[2], a[0]);
	and _ECO_93(w_eco93, !a[4], !b[4], a[6], b[6], a[1], a[2], !b[0]);
	and _ECO_94(w_eco94, !b[3], !b[4], a[6], b[6], !b[1], !b[2], !b[0]);
	and _ECO_95(w_eco95, b[3], !b[4], a[5], !b[1], a[0], op[0]);
	and _ECO_96(w_eco96, b[3], !b[4], a[5], a[1], !b[0], op[0]);
	and _ECO_97(w_eco97, !b[4], a[5], !b[1], a[2], a[0], op[0]);
	and _ECO_98(w_eco98, !b[4], a[5], a[1], a[2], !b[0], op[0]);
	and _ECO_99(w_eco99, b[3], !b[4], a[5], !b[1], !b[0], op[1]);
	and _ECO_100(w_eco100, !b[4], a[5], !b[1], a[2], !b[0], op[1]);
	and _ECO_101(w_eco101, !b[4], a[5], !b[1], !b[2], !b[0], op[0]);
	and _ECO_102(w_eco102, b[3], !a[5], !b[5], a[6], b[6], !b[1], a[0]);
	and _ECO_103(w_eco103, b[3], !a[5], !b[5], a[6], b[6], a[1], !b[0]);
	and _ECO_104(w_eco104, !a[5], !b[5], a[6], b[6], !b[1], a[2], a[0]);
	and _ECO_105(w_eco105, !a[5], !b[5], a[6], b[6], a[1], a[2], !b[0]);
	and _ECO_106(w_eco106, b[3], a[4], !b[5], !b[1], a[0], op[0]);
	and _ECO_107(w_eco107, b[3], a[4], !b[5], a[1], !b[0], op[0]);
	and _ECO_108(w_eco108, a[4], !b[5], !b[1], a[2], a[0], op[0]);
	and _ECO_109(w_eco109, a[4], !b[5], a[1], a[2], !b[0], op[0]);
	and _ECO_110(w_eco110, b[3], a[4], !b[5], !b[1], !b[0], op[1]);
	and _ECO_111(w_eco111, a[4], !b[5], !b[1], a[2], !b[0], op[1]);
	and _ECO_112(w_eco112, a[4], !b[5], !b[1], !b[2], !b[0], op[0]);
	and _ECO_113(w_eco113, b[3], !b[4], !b[5], !b[1], !b[0], op[0]);
	and _ECO_114(w_eco114, !b[4], !b[5], !b[1], a[2], !b[0], op[0]);
	and _ECO_115(w_eco115, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_116(w_eco116, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_117(w_eco117, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0]);
	and _ECO_118(w_eco118, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0]);
	and _ECO_119(w_eco119, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0]);
	and _ECO_120(w_eco120, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0]);
	and _ECO_121(w_eco121, !a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !b[0]);
	and _ECO_122(w_eco122, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0]);
	and _ECO_123(w_eco123, !b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_124(w_eco124, !a[3], a[5], b[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_125(w_eco125, !b[3], !a[4], a[5], b[5], b[6], !b[1], !a[2], !a[0]);
	and _ECO_126(w_eco126, !b[3], !a[4], a[5], b[5], b[6], !a[1], !a[2], !b[0]);
	and _ECO_127(w_eco127, !a[3], a[5], b[5], b[6], !b[1], !a[2], !a[0]);
	and _ECO_128(w_eco128, !a[3], a[5], b[5], b[6], !a[1], !a[2], !b[0]);
	and _ECO_129(w_eco129, !a[3], a[4], a[5], b[5], a[6], !b[1], !a[2], !b[0]);
	and _ECO_130(w_eco130, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[0]);
	and _ECO_131(w_eco131, b[3], !a[4], !b[4], a[5], b[5], a[6], b[2]);
	and _ECO_132(w_eco132, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0]);
	and _ECO_133(w_eco133, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2]);
	and _ECO_134(w_eco134, !a[3], !b[3], !b[4], a[5], b[5], a[6], b[2]);
	and _ECO_135(w_eco135, !b[3], !b[4], a[5], b[5], a[6], !b[1], !a[2], !b[2], a[0]);
	and _ECO_136(w_eco136, !b[3], !b[4], a[5], b[5], a[6], a[1], !a[2], !b[2], !b[0]);
	and _ECO_137(w_eco137, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_138(w_eco138, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0]);
	and _ECO_139(w_eco139, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0]);
	and _ECO_140(w_eco140, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0]);
	and _ECO_141(w_eco141, !b[3], !a[4], !a[5], a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_142(w_eco142, !a[3], !a[5], a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_143(w_eco143, !a[3], a[4], a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_144(w_eco144, b[3], a[4], a[5], a[1], a[0], op[0]);
	and _ECO_145(w_eco145, b[3], a[4], a[5], b[2], op[0]);
	and _ECO_146(w_eco146, a[4], a[5], a[1], a[2], a[0], op[0]);
	and _ECO_147(w_eco147, a[4], a[5], a[1], !b[1], a[2], op[0]);
	and _ECO_148(w_eco148, !a[3], a[4], a[5], b[2], op[0]);
	and _ECO_149(w_eco149, b[3], a[4], a[5], !b[1], a[0], op[1]);
	and _ECO_150(w_eco150, b[3], a[4], a[5], a[1], !b[0], op[1]);
	and _ECO_151(w_eco151, a[4], a[5], !b[1], a[2], a[0], op[1]);
	and _ECO_152(w_eco152, a[4], a[5], a[1], a[2], !b[0], op[1]);
	and _ECO_153(w_eco153, a[4], a[5], !b[1], !b[2], a[0], op[0]);
	and _ECO_154(w_eco154, a[4], a[5], a[1], !b[2], !b[0], op[0]);
	and _ECO_155(w_eco155, a[4], a[5], !b[1], !b[2], !b[0], op[1]);
	and _ECO_156(w_eco156, b[3], !a[4], !b[4], a[6], b[6], a[1], a[0]);
	and _ECO_157(w_eco157, b[3], !a[4], !b[4], a[6], b[6], b[2]);
	and _ECO_158(w_eco158, !a[4], !b[4], a[6], b[6], a[1], a[2], a[0]);
	and _ECO_159(w_eco159, !a[4], !b[4], a[6], b[6], a[1], !b[1], a[2]);
	and _ECO_160(w_eco160, !a[3], !b[3], !b[4], a[6], b[6], b[2]);
	and _ECO_161(w_eco161, !b[3], !b[4], a[6], b[6], !b[1], !a[2], !b[2], a[0]);
	and _ECO_162(w_eco162, !b[3], !b[4], a[6], b[6], a[1], !a[2], !b[2], !b[0]);
	and _ECO_163(w_eco163, b[3], !b[4], a[5], a[1], a[0], op[0]);
	and _ECO_164(w_eco164, b[3], !b[4], a[5], b[2], op[0]);
	and _ECO_165(w_eco165, !b[4], a[5], a[1], a[2], a[0], op[0]);
	and _ECO_166(w_eco166, !b[4], a[5], a[1], !b[1], a[2], op[0]);
	and _ECO_167(w_eco167, !a[3], !b[4], a[5], b[2], op[0]);
	and _ECO_168(w_eco168, b[3], !b[4], a[5], !b[1], a[0], op[1]);
	and _ECO_169(w_eco169, b[3], !b[4], a[5], a[1], !b[0], op[1]);
	and _ECO_170(w_eco170, !b[4], a[5], !b[1], a[2], a[0], op[1]);
	and _ECO_171(w_eco171, !b[4], a[5], a[1], a[2], !b[0], op[1]);
	and _ECO_172(w_eco172, !b[4], a[5], !b[1], !b[2], a[0], op[0]);
	and _ECO_173(w_eco173, !b[4], a[5], a[1], !b[2], !b[0], op[0]);
	and _ECO_174(w_eco174, !b[4], a[5], !b[1], !b[2], !b[0], op[1]);
	and _ECO_175(w_eco175, b[3], !a[5], !b[5], a[6], b[6], a[1], a[0]);
	and _ECO_176(w_eco176, b[3], !a[5], !b[5], a[6], b[6], b[2]);
	and _ECO_177(w_eco177, !a[5], !b[5], a[6], b[6], a[1], a[2], a[0]);
	and _ECO_178(w_eco178, !a[5], !b[5], a[6], b[6], a[1], !b[1], a[2]);
	and _ECO_179(w_eco179, b[3], a[4], !b[5], a[1], a[0], op[0]);
	and _ECO_180(w_eco180, b[3], a[4], !b[5], b[2], op[0]);
	and _ECO_181(w_eco181, a[4], !b[5], a[1], a[2], a[0], op[0]);
	and _ECO_182(w_eco182, a[4], !b[5], a[1], !b[1], a[2], op[0]);
	and _ECO_183(w_eco183, !a[3], a[4], !b[5], b[2], op[0]);
	and _ECO_184(w_eco184, b[3], a[4], !b[5], !b[1], a[0], op[1]);
	and _ECO_185(w_eco185, b[3], a[4], !b[5], a[1], !b[0], op[1]);
	and _ECO_186(w_eco186, a[4], !b[5], !b[1], a[2], a[0], op[1]);
	and _ECO_187(w_eco187, a[4], !b[5], a[1], a[2], !b[0], op[1]);
	and _ECO_188(w_eco188, a[4], !b[5], !b[1], !b[2], a[0], op[0]);
	and _ECO_189(w_eco189, a[4], !b[5], a[1], !b[2], !b[0], op[0]);
	and _ECO_190(w_eco190, a[4], !b[5], !b[1], !b[2], !b[0], op[1]);
	and _ECO_191(w_eco191, b[3], !b[4], !b[5], !b[1], a[0], op[0]);
	and _ECO_192(w_eco192, b[3], !b[4], !b[5], a[1], !b[0], op[0]);
	and _ECO_193(w_eco193, !b[4], !b[5], !b[1], a[2], a[0], op[0]);
	and _ECO_194(w_eco194, !b[4], !b[5], a[1], a[2], !b[0], op[0]);
	and _ECO_195(w_eco195, b[3], !b[4], !b[5], !b[1], !b[0], op[1]);
	and _ECO_196(w_eco196, !b[4], !b[5], !b[1], a[2], !b[0], op[1]);
	and _ECO_197(w_eco197, !b[4], !b[5], !b[1], !b[2], !b[0], op[0]);
	and _ECO_198(w_eco198, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0]);
	and _ECO_199(w_eco199, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0]);
	and _ECO_200(w_eco200, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0]);
	and _ECO_201(w_eco201, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0]);
	and _ECO_202(w_eco202, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2]);
	and _ECO_203(w_eco203, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2]);
	and _ECO_204(w_eco204, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0]);
	and _ECO_205(w_eco205, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0]);
	and _ECO_206(w_eco206, !a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], a[0]);
	and _ECO_207(w_eco207, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !b[0]);
	and _ECO_208(w_eco208, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0]);
	and _ECO_209(w_eco209, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0]);
	and _ECO_210(w_eco210, !b[3], !a[4], a[5], b[5], b[6], !b[1], !b[2], !a[0]);
	and _ECO_211(w_eco211, !b[3], !a[4], a[5], b[5], b[6], !a[1], !b[2], !b[0]);
	and _ECO_212(w_eco212, !a[3], b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0]);
	and _ECO_213(w_eco213, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[2], !b[0]);
	and _ECO_214(w_eco214, !b[3], !a[4], a[5], b[5], b[6], !a[2], !b[2]);
	and _ECO_215(w_eco215, !a[3], a[5], b[5], b[6], !a[2], !b[2]);
	and _ECO_216(w_eco216, !b[3], a[5], b[5], !a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_217(w_eco217, !b[3], a[5], b[5], !a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_218(w_eco218, !a[3], a[4], a[5], b[5], a[6], !b[1], !b[2], !b[0]);
	and _ECO_219(w_eco219, !a[3], a[4], a[5], b[5], a[6], !b[1], !a[2], !a[0]);
	and _ECO_220(w_eco220, !a[3], a[4], a[5], b[5], a[6], !a[1], !a[2], !b[0]);
	and _ECO_221(w_eco221, !b[3], !b[4], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0]);
	and _ECO_222(w_eco222, !b[3], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0]);
	and _ECO_223(w_eco223, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0]);
	and _ECO_224(w_eco224, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0]);
	and _ECO_225(w_eco225, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2]);
	and _ECO_226(w_eco226, !b[3], !a[5], a[6], b[6], !b[1], !b[2], !b[0]);
	and _ECO_227(w_eco227, !a[3], !a[5], a[6], b[6], !b[1], !b[2], !b[0]);
	and _ECO_228(w_eco228, !b[3], !a[4], !a[5], a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_229(w_eco229, !b[3], !a[4], !a[5], a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_230(w_eco230, !a[3], !a[5], a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_231(w_eco231, !a[3], !a[5], a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_232(w_eco232, !b[3], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_233(w_eco233, !b[3], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_234(w_eco234, !b[3], a[4], b[4], a[5], !a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_235(w_eco235, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_236(w_eco236, !a[3], a[4], a[6], b[6], !b[1], !b[2], !b[0]);
	and _ECO_237(w_eco237, !a[3], a[4], a[6], b[6], !b[1], !a[2], !a[0]);
	and _ECO_238(w_eco238, !a[3], a[4], a[6], b[6], !a[1], !a[2], !b[0]);
	and _ECO_239(w_eco239, b[3], a[4], a[5], a[1], a[0], op[1]);
	and _ECO_240(w_eco240, b[3], a[4], a[5], b[2], op[1]);
	and _ECO_241(w_eco241, a[4], a[5], a[1], a[2], a[0], op[1]);
	and _ECO_242(w_eco242, a[4], a[5], a[1], !b[1], a[2], op[1]);
	and _ECO_243(w_eco243, !a[3], a[4], a[5], b[2], op[1]);
	and _ECO_244(w_eco244, a[4], a[5], a[1], !b[2], a[0], op[0]);
	and _ECO_245(w_eco245, a[4], a[5], a[1], !b[1], !b[2], op[0]);
	and _ECO_246(w_eco246, a[4], a[5], !b[1], !b[2], a[0], op[1]);
	and _ECO_247(w_eco247, a[4], a[5], a[1], !b[2], !b[0], op[1]);
	and _ECO_248(w_eco248, !b[3], !b[4], a[6], b[6], a[1], !a[2], !b[2], a[0]);
	and _ECO_249(w_eco249, !b[3], !b[4], a[6], b[6], a[1], !b[1], !b[2], !a[0]);
	and _ECO_250(w_eco250, b[3], !b[4], a[5], a[1], a[0], op[1]);
	and _ECO_251(w_eco251, b[3], !b[4], a[5], b[2], op[1]);
	and _ECO_252(w_eco252, !b[4], a[5], a[1], a[2], a[0], op[1]);
	and _ECO_253(w_eco253, !b[4], a[5], a[1], !b[1], a[2], op[1]);
	and _ECO_254(w_eco254, !a[3], !b[4], a[5], b[2], op[1]);
	and _ECO_255(w_eco255, !b[4], a[5], a[1], !b[2], a[0], op[0]);
	and _ECO_256(w_eco256, !b[4], a[5], a[1], !b[1], !b[2], op[0]);
	and _ECO_257(w_eco257, !b[4], a[5], !b[1], !b[2], a[0], op[1]);
	and _ECO_258(w_eco258, !b[4], a[5], a[1], !b[2], !b[0], op[1]);
	and _ECO_259(w_eco259, b[3], a[4], !b[5], a[1], a[0], op[1]);
	and _ECO_260(w_eco260, b[3], a[4], !b[5], b[2], op[1]);
	and _ECO_261(w_eco261, a[4], !b[5], a[1], a[2], a[0], op[1]);
	and _ECO_262(w_eco262, a[4], !b[5], a[1], !b[1], a[2], op[1]);
	and _ECO_263(w_eco263, !a[3], a[4], !b[5], b[2], op[1]);
	and _ECO_264(w_eco264, a[4], !b[5], a[1], !b[2], a[0], op[0]);
	and _ECO_265(w_eco265, a[4], !b[5], a[1], !b[1], !b[2], op[0]);
	and _ECO_266(w_eco266, a[4], !b[5], !b[1], !b[2], a[0], op[1]);
	and _ECO_267(w_eco267, a[4], !b[5], a[1], !b[2], !b[0], op[1]);
	and _ECO_268(w_eco268, b[3], !b[4], !b[5], a[1], a[0], op[0]);
	and _ECO_269(w_eco269, b[3], !b[4], !b[5], b[2], op[0]);
	and _ECO_270(w_eco270, !b[4], !b[5], a[1], a[2], a[0], op[0]);
	and _ECO_271(w_eco271, !b[4], !b[5], a[1], !b[1], a[2], op[0]);
	and _ECO_272(w_eco272, !a[3], !b[4], !b[5], b[2], op[0]);
	and _ECO_273(w_eco273, b[3], !b[4], !b[5], !b[1], a[0], op[1]);
	and _ECO_274(w_eco274, b[3], !b[4], !b[5], a[1], !b[0], op[1]);
	and _ECO_275(w_eco275, !b[4], !b[5], !b[1], a[2], a[0], op[1]);
	and _ECO_276(w_eco276, !b[4], !b[5], a[1], a[2], !b[0], op[1]);
	and _ECO_277(w_eco277, !b[4], !b[5], !b[1], !b[2], a[0], op[0]);
	and _ECO_278(w_eco278, !b[4], !b[5], a[1], !b[2], !b[0], op[0]);
	and _ECO_279(w_eco279, !b[4], !b[5], !b[1], !b[2], !b[0], op[1]);
	and _ECO_280(w_eco280, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0]);
	and _ECO_281(w_eco281, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_282(w_eco282, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0]);
	and _ECO_283(w_eco283, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_284(w_eco284, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0]);
	and _ECO_285(w_eco285, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2]);
	and _ECO_286(w_eco286, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0]);
	and _ECO_287(w_eco287, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2]);
	and _ECO_288(w_eco288, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0]);
	and _ECO_289(w_eco289, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0]);
	and _ECO_290(w_eco290, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], a[0]);
	and _ECO_291(w_eco291, !a[3], !b[3], a[4], b[4], a[5], a[6], b[2]);
	and _ECO_292(w_eco292, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[2], a[0]);
	and _ECO_293(w_eco293, !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], !b[0]);
	and _ECO_294(w_eco294, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2]);
	and _ECO_295(w_eco295, !b[3], !a[4], a[5], b[5], b[6], !a[1], !b[2], !a[0]);
	and _ECO_296(w_eco296, !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_297(w_eco297, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0]);
	and _ECO_298(w_eco298, !a[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_299(w_eco299, !b[3], !a[4], a[5], b[5], b[6], !a[1], !a[2], !a[0]);
	and _ECO_300(w_eco300, !b[3], !a[4], a[5], b[5], b[6], !a[1], !b[1], !a[2]);
	and _ECO_301(w_eco301, !a[3], a[5], b[5], b[6], !a[1], !a[2], !a[0]);
	and _ECO_302(w_eco302, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2]);
	and _ECO_303(w_eco303, !a[3], !b[3], a[4], a[6], b[6], a[1], a[0]);
	and _ECO_304(w_eco304, !b[3], a[5], b[5], !a[6], b[6], !b[1], !b[2], !a[0]);
	and _ECO_305(w_eco305, !b[3], a[5], b[5], !a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_306(w_eco306, !b[3], a[5], b[5], !a[6], b[6], !a[2], !b[2]);
	and _ECO_307(w_eco307, !a[3], b[3], a[4], a[5], b[5], a[6], !b[1], !b[2], !a[0]);
	and _ECO_308(w_eco308, !a[3], b[3], a[4], a[5], b[5], a[6], !a[1], !b[2], !b[0]);
	and _ECO_309(w_eco309, !a[3], !b[3], a[4], a[5], b[5], a[6], !b[1], a[0]);
	and _ECO_310(w_eco310, !a[3], !b[3], a[4], a[5], b[5], a[6], a[1], !b[0]);
	and _ECO_311(w_eco311, !a[3], a[4], a[5], b[5], a[6], !a[2], !b[2]);
	and _ECO_312(w_eco312, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2]);
	and _ECO_313(w_eco313, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0]);
	and _ECO_314(w_eco314, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2]);
	and _ECO_315(w_eco315, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0]);
	and _ECO_316(w_eco316, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2]);
	and _ECO_317(w_eco317, !b[3], !a[4], !a[5], a[6], b[6], !b[1], !b[2], !a[0]);
	and _ECO_318(w_eco318, !b[3], !a[4], !a[5], a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_319(w_eco319, !a[3], b[3], !a[5], a[6], b[6], !b[1], !b[2], !a[0]);
	and _ECO_320(w_eco320, !a[3], b[3], !a[5], a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_321(w_eco321, !b[3], !a[4], !a[5], a[6], b[6], !a[2], !b[2]);
	and _ECO_322(w_eco322, !a[3], !a[5], a[6], b[6], !a[2], !b[2]);
	and _ECO_323(w_eco323, !b[3], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2]);
	and _ECO_324(w_eco324, !b[3], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_325(w_eco325, !b[3], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0]);
	and _ECO_326(w_eco326, !b[3], a[4], a[6], b[6], a[1], !b[1], !b[2], !a[0]);
	and _ECO_327(w_eco327, !b[3], a[4], a[6], b[6], a[1], !a[2], !b[2], a[0]);
	and _ECO_328(w_eco328, !b[3], a[4], b[4], a[5], !a[6], b[6], !b[1], !b[2], !a[0]);
	and _ECO_329(w_eco329, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_330(w_eco330, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[2], !b[2]);
	and _ECO_331(w_eco331, !a[3], b[3], a[4], a[6], b[6], !b[1], !b[2], !a[0]);
	and _ECO_332(w_eco332, !a[3], b[3], a[4], a[6], b[6], !a[1], !b[2], !b[0]);
	and _ECO_333(w_eco333, !a[3], a[4], a[6], b[6], !a[2], !b[2]);
	and _ECO_334(w_eco334, a[4], a[5], a[1], !b[2], a[0], op[1]);
	and _ECO_335(w_eco335, a[4], a[5], a[1], !b[1], !b[2], op[1]);
	and _ECO_336(w_eco336, !b[4], a[5], a[1], !b[2], a[0], op[1]);
	and _ECO_337(w_eco337, !b[4], a[5], a[1], !b[1], !b[2], op[1]);
	and _ECO_338(w_eco338, a[4], !b[5], a[1], !b[2], a[0], op[1]);
	and _ECO_339(w_eco339, a[4], !b[5], a[1], !b[1], !b[2], op[1]);
	and _ECO_340(w_eco340, b[3], !b[4], !b[5], a[1], a[0], op[1]);
	and _ECO_341(w_eco341, b[3], !b[4], !b[5], b[2], op[1]);
	and _ECO_342(w_eco342, !b[4], !b[5], a[1], a[2], a[0], op[1]);
	and _ECO_343(w_eco343, !b[4], !b[5], a[1], !b[1], a[2], op[1]);
	and _ECO_344(w_eco344, !a[3], !b[4], !b[5], b[2], op[1]);
	and _ECO_345(w_eco345, !b[4], !b[5], a[1], !b[2], a[0], op[0]);
	and _ECO_346(w_eco346, !b[4], !b[5], a[1], !b[1], !b[2], op[0]);
	and _ECO_347(w_eco347, !b[4], !b[5], !b[1], !b[2], a[0], op[1]);
	and _ECO_348(w_eco348, !b[4], !b[5], a[1], !b[2], !b[0], op[1]);
	and _ECO_349(w_eco349, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_350(w_eco350, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !a[0]);
	and _ECO_351(w_eco351, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0]);
	and _ECO_352(w_eco352, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_353(w_eco353, !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0]);
	and _ECO_354(w_eco354, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0]);
	and _ECO_355(w_eco355, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2]);
	and _ECO_356(w_eco356, !b[3], a[5], b[5], !a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_357(w_eco357, !b[3], a[5], b[5], !a[6], b[6], !a[1], !a[2], !a[0]);
	and _ECO_358(w_eco358, !b[3], a[5], b[5], !a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_359(w_eco359, !b[3], a[5], b[5], !a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_360(w_eco360, !b[3], a[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_361(w_eco361, !a[3], b[3], a[4], a[5], b[5], a[6], !a[1], !b[2], !a[0]);
	and _ECO_362(w_eco362, !a[3], a[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_363(w_eco363, !a[3], !b[3], a[4], a[5], b[5], a[6], a[1], a[0]);
	and _ECO_364(w_eco364, !a[3], a[4], a[5], b[5], a[6], !a[1], !a[2], !a[0]);
	and _ECO_365(w_eco365, !a[3], a[4], a[5], b[5], a[6], !a[1], !b[1], !a[2]);
	and _ECO_366(w_eco366, !b[3], !a[4], !a[5], a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_367(w_eco367, !a[3], b[3], !a[5], a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_368(w_eco368, !a[3], !a[5], a[6], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_369(w_eco369, !b[3], !a[4], !a[5], a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_370(w_eco370, !a[3], !a[5], a[6], b[6], !a[1], !a[2], !a[0]);
	and _ECO_371(w_eco371, !a[3], !a[5], a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_372(w_eco372, !b[3], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_373(w_eco373, !b[3], !a[5], b[5], a[6], b[6], !a[2], !b[2]);
	and _ECO_374(w_eco374, !b[3], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_375(w_eco375, !b[3], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_376(w_eco376, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_377(w_eco377, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[1], !a[2], !a[0]);
	and _ECO_378(w_eco378, !b[3], a[4], b[4], a[5], !a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_379(w_eco379, !b[3], a[4], b[4], a[5], !a[6], b[6], !b[1], !a[2], !b[0]);
	and _ECO_380(w_eco380, !b[3], a[4], a[6], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_381(w_eco381, !a[3], b[3], a[4], a[6], b[6], !a[1], !b[2], !a[0]);
	and _ECO_382(w_eco382, !a[3], a[4], a[6], b[6], !a[1], !b[1], !b[2], a[0]);
	and _ECO_383(w_eco383, !a[3], !b[3], a[4], a[6], b[6], a[1], !b[0]);
	and _ECO_384(w_eco384, !a[3], a[4], a[6], b[6], !a[1], !a[2], !a[0]);
	and _ECO_385(w_eco385, !a[3], a[4], a[6], b[6], !a[1], !b[1], !a[2]);
	and _ECO_386(w_eco386, !b[4], !b[5], a[1], !b[2], a[0], op[1]);
	and _ECO_387(w_eco387, !b[4], !b[5], a[1], !b[1], !b[2], op[1]);
	or _ECO_388(w_eco388, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387);
	xor _ECO_out0(y[7], sub_wire0, w_eco388);

endmodule