//
// Conformal-LEC: Version 11.10-d208 (10-Mar-2012) (64 bit executable)
//
module top(scr_out, scr_in, scr_init, scr_run, clk, reset, scr_out_p, set);
input  scr_init, scr_run, clk, reset, set;
input   [31:0] scr_out;
input   [31:0] scr_in;
output  [31:0] scr_out_p;
wire  \scr_ff_mux_state_427_13_g758/w_0 , \scr_ff_mux_state_427_13_g758/w_1 , 
    \scr_ff_mux_state_427_13_g758/w_2 , \scr_ff_mux_state_427_13_g758/w_3 , 
    \scr_ff_mux_state_427_13_g758/w_4 , \scr_ff_mux_state_427_13_g746/w_0 , 
    \scr_ff_mux_state_427_13_g746/w_1 , \scr_ff_mux_state_427_13_g746/w_2 , 
    \scr_ff_mux_state_427_13_g746/w_3 , \scr_ff_mux_state_427_13_g746/w_4 , 
    \scr_ff_mux_state_427_13_g730/w_0 , \scr_ff_mux_state_427_13_g730/w_1 , 
    \scr_ff_mux_state_427_13_g730/w_2 , \scr_ff_mux_state_427_13_g730/w_3 , 
    \scr_ff_mux_state_427_13_g730/w_4 , \scr_ff_mux_state_427_13_g718/w_0 , 
    \scr_ff_mux_state_427_13_g718/w_1 , \scr_ff_mux_state_427_13_g718/w_2 , 
    \scr_ff_mux_state_427_13_g718/w_3 , \scr_ff_mux_state_427_13_g718/w_4 , 
    \scr_ff_mux_state_427_13_g702/w_0 , \scr_ff_mux_state_427_13_g702/w_1 , 
    \scr_ff_mux_state_427_13_g702/w_2 , \scr_ff_mux_state_427_13_g702/w_3 , 
    \scr_ff_mux_state_427_13_g702/w_4 , \scr_ff_mux_state_427_13_g690/w_0 , 
    \scr_ff_mux_state_427_13_g690/w_1 , \scr_ff_mux_state_427_13_g690/w_2 , 
    \scr_ff_mux_state_427_13_g690/w_3 , \scr_ff_mux_state_427_13_g690/w_4 , 
    \scr_ff_mux_state_427_13_g674/w_0 , \scr_ff_mux_state_427_13_g674/w_1 , 
    \scr_ff_mux_state_427_13_g674/w_2 , \scr_ff_mux_state_427_13_g674/w_3 , 
    \scr_ff_mux_state_427_13_g674/w_4 , \scr_ff_mux_state_427_13_g662/w_0 , 
    \scr_ff_mux_state_427_13_g662/w_1 , \scr_ff_mux_state_427_13_g662/w_2 , 
    \scr_ff_mux_state_427_13_g662/w_3 , \scr_ff_mux_state_427_13_g662/w_4 , 
    \scr_ff_mux_state_427_13_g646/w_0 , \scr_ff_mux_state_427_13_g646/w_1 , 
    \scr_ff_mux_state_427_13_g646/w_2 , \scr_ff_mux_state_427_13_g646/w_3 , 
    \scr_ff_mux_state_427_13_g646/w_4 , \scr_ff_mux_state_427_13_g634/w_0 , 
    \scr_ff_mux_state_427_13_g634/w_1 , \scr_ff_mux_state_427_13_g634/w_2 , 
    \scr_ff_mux_state_427_13_g634/w_3 , \scr_ff_mux_state_427_13_g634/w_4 , 
    \scr_ff_mux_state_427_13_g618/w_0 , \scr_ff_mux_state_427_13_g618/w_1 , 
    \scr_ff_mux_state_427_13_g618/w_2 , \scr_ff_mux_state_427_13_g618/w_3 , 
    \scr_ff_mux_state_427_13_g618/w_4 , \scr_ff_mux_state_427_13_g606/w_0 , 
    \scr_ff_mux_state_427_13_g606/w_1 , \scr_ff_mux_state_427_13_g606/w_2 , 
    \scr_ff_mux_state_427_13_g606/w_3 , \scr_ff_mux_state_427_13_g606/w_4 , 
    \scr_ff_mux_state_427_13_g590/w_0 , \scr_ff_mux_state_427_13_g590/w_1 , 
    \scr_ff_mux_state_427_13_g590/w_2 , \scr_ff_mux_state_427_13_g590/w_3 , 
    \scr_ff_mux_state_427_13_g590/w_4 , \scr_ff_mux_state_427_13_g578/w_0 , 
    \scr_ff_mux_state_427_13_g578/w_1 , \scr_ff_mux_state_427_13_g578/w_2 , 
    \scr_ff_mux_state_427_13_g578/w_3 , \scr_ff_mux_state_427_13_g578/w_4 , 
    \scr_ff_mux_state_427_13_g562/w_0 , \scr_ff_mux_state_427_13_g562/w_1 , 
    \scr_ff_mux_state_427_13_g562/w_2 , \scr_ff_mux_state_427_13_g562/w_3 , 
    \scr_ff_mux_state_427_13_g562/w_4 , \scr_ff_mux_state_427_13_g550/w_0 , 
    \scr_ff_mux_state_427_13_g550/w_1 , \scr_ff_mux_state_427_13_g550/w_2 , 
    \scr_ff_mux_state_427_13_g550/w_3 , \scr_ff_mux_state_427_13_g550/w_4 , 
    \scr_ff_mux_state_427_13_g534/w_0 , \scr_ff_mux_state_427_13_g534/w_1 , 
    \scr_ff_mux_state_427_13_g534/w_2 , \scr_ff_mux_state_427_13_g534/w_3 , 
    \scr_ff_mux_state_427_13_g534/w_4 , \scr_ff_mux_state_427_13_g522/w_0 , 
    \scr_ff_mux_state_427_13_g522/w_1 , \scr_ff_mux_state_427_13_g522/w_2 , 
    \scr_ff_mux_state_427_13_g522/w_3 , \scr_ff_mux_state_427_13_g522/w_4 , 
    \scr_ff_mux_state_427_13_g506/w_0 , \scr_ff_mux_state_427_13_g506/w_1 , 
    \scr_ff_mux_state_427_13_g506/w_2 , \scr_ff_mux_state_427_13_g506/w_3 , 
    \scr_ff_mux_state_427_13_g506/w_4 , \scr_ff_mux_state_427_13_g494/w_0 , 
    \scr_ff_mux_state_427_13_g494/w_1 , \scr_ff_mux_state_427_13_g494/w_2 , 
    \scr_ff_mux_state_427_13_g494/w_3 , \scr_ff_mux_state_427_13_g494/w_4 , 
    \scr_ff_mux_state_427_13_g478/w_0 , \scr_ff_mux_state_427_13_g478/w_1 , 
    \scr_ff_mux_state_427_13_g478/w_2 , \scr_ff_mux_state_427_13_g478/w_3 , 
    \scr_ff_mux_state_427_13_g478/w_4 , \scr_ff_mux_state_427_13_g466/w_0 , 
    \scr_ff_mux_state_427_13_g466/w_1 , \scr_ff_mux_state_427_13_g466/w_2 , 
    \scr_ff_mux_state_427_13_g466/w_3 , \scr_ff_mux_state_427_13_g466/w_4 , 
    \scr_ff_mux_state_427_13_g450/w_0 , \scr_ff_mux_state_427_13_g450/w_1 , 
    \scr_ff_mux_state_427_13_g450/w_2 , \scr_ff_mux_state_427_13_g450/w_3 , 
    \scr_ff_mux_state_427_13_g450/w_4 , \scr_ff_mux_state_427_13_g438/w_0 , 
    \scr_ff_mux_state_427_13_g438/w_1 , \scr_ff_mux_state_427_13_g438/w_2 , 
    \scr_ff_mux_state_427_13_g438/w_3 , \scr_ff_mux_state_427_13_g438/w_4 , 
    \scr_ff_mux_state_427_13_g422/w_0 , \scr_ff_mux_state_427_13_g422/w_1 , 
    \scr_ff_mux_state_427_13_g422/w_2 , \scr_ff_mux_state_427_13_g422/w_3 , 
    \scr_ff_mux_state_427_13_g422/w_4 , \scr_ff_mux_state_427_13_g410/w_0 , 
    \scr_ff_mux_state_427_13_g410/w_1 , \scr_ff_mux_state_427_13_g410/w_2 , 
    \scr_ff_mux_state_427_13_g410/w_3 , \scr_ff_mux_state_427_13_g410/w_4 , 
    \scr_ff_mux_state_427_13_g394/w_0 , \scr_ff_mux_state_427_13_g394/w_1 , 
    \scr_ff_mux_state_427_13_g394/w_2 , \scr_ff_mux_state_427_13_g394/w_3 , 
    \scr_ff_mux_state_427_13_g394/w_4 , \scr_ff_mux_state_427_13_g382/w_0 , 
    \scr_ff_mux_state_427_13_g382/w_1 , \scr_ff_mux_state_427_13_g382/w_2 , 
    \scr_ff_mux_state_427_13_g382/w_3 , \scr_ff_mux_state_427_13_g382/w_4 , 
    \scr_ff_mux_state_427_13_g366/w_0 , \scr_ff_mux_state_427_13_g366/w_1 , 
    \scr_ff_mux_state_427_13_g366/w_2 , \scr_ff_mux_state_427_13_g366/w_3 , 
    \scr_ff_mux_state_427_13_g366/w_4 , \scr_ff_mux_state_427_13_g354/w_0 , 
    \scr_ff_mux_state_427_13_g354/w_1 , \scr_ff_mux_state_427_13_g354/w_2 , 
    \scr_ff_mux_state_427_13_g354/w_3 , \scr_ff_mux_state_427_13_g354/w_4 , 
    \scr_ff_mux_state_427_13_g338/w_0 , \scr_ff_mux_state_427_13_g338/w_1 , 
    \scr_ff_mux_state_427_13_g338/w_2 , \scr_ff_mux_state_427_13_g338/w_3 , 
    \scr_ff_mux_state_427_13_g338/w_4 , \scr_ff_mux_state_427_13_g326/w_0 , 
    \scr_ff_mux_state_427_13_g326/w_1 , \scr_ff_mux_state_427_13_g326/w_2 , 
    \scr_ff_mux_state_427_13_g326/w_3 , \scr_ff_mux_state_427_13_g326/w_4 , 
    n_1120, n_1119, n_1118, n_392, n_391, n_390, n_389, n_370, n_369, n_367, 
    n_366, n_363, n_362, n_361, n_358, n_357, n_356, n_353, n_352, n_351, 
    n_348, n_347, n_346, n_344, n_343, n_342, n_341, n_338, n_337, n_336, 
    n_335, n_334, n_331, n_330, n_329, n_328, n_327, n_326, n_325, n_324, 
    n_323, n_322, n_321, n_320, n_318, n_317, n_316, n_315, n_314, n_312, 
    n_311, n_310, n_309, n_308, n_307, n_305, n_304, n_303, n_302, n_301, 
    n_300, n_299, n_298, n_297, n_296, n_295, n_294, n_293, n_292, n_291, 
    n_290, n_287, n_286, n_285, n_284, n_283, n_282, n_281, n_280, n_279, 
    n_278, n_277, n_276, n_275, n_274, n_273, n_272, n_271, n_270, n_269, 
    n_268, n_267, n_266, n_219, n_214, n_209, n_199, n_198, n_192, n_191, 
    n_185, n_184, n_178, n_177, n_171, n_170, n_111, n_101, n_100, n_96, n_95, 
    n_94, n_93, n_90, n_89, n_88, n_87, n_84, n_81, n_80, n_76, n_75, n_74, 
    n_73, n_72, a15, \a14[0] , \a13[0] , \a12[0] , \a11[0] , \a10[0] , \a9[0] , 
    \a8[0] , \a7[0] , \a6[0] , \a5[0] , \a4[0] , set, reset, clk, scr_run, 
    scr_init;
wire  \scr_ff_mux_state_427_13_g758/data3 , \scr_ff_mux_state_427_13_g758/data4 , 
    \scr_ff_mux_state_427_13_g746/data3 , \scr_ff_mux_state_427_13_g746/data4 , 
    \scr_ff_mux_state_427_13_g730/data3 , \scr_ff_mux_state_427_13_g730/data4 , 
    \scr_ff_mux_state_427_13_g718/data3 , \scr_ff_mux_state_427_13_g718/data4 , 
    \scr_ff_mux_state_427_13_g702/data3 , \scr_ff_mux_state_427_13_g702/data4 , 
    \scr_ff_mux_state_427_13_g690/data3 , \scr_ff_mux_state_427_13_g690/data4 , 
    \scr_ff_mux_state_427_13_g674/data3 , \scr_ff_mux_state_427_13_g674/data4 , 
    \scr_ff_mux_state_427_13_g662/data3 , \scr_ff_mux_state_427_13_g662/data4 , 
    \scr_ff_mux_state_427_13_g646/data3 , \scr_ff_mux_state_427_13_g646/data4 , 
    \scr_ff_mux_state_427_13_g634/data3 , \scr_ff_mux_state_427_13_g634/data4 , 
    \scr_ff_mux_state_427_13_g618/data3 , \scr_ff_mux_state_427_13_g618/data4 , 
    \scr_ff_mux_state_427_13_g606/data3 , \scr_ff_mux_state_427_13_g606/data4 , 
    \scr_ff_mux_state_427_13_g590/data3 , \scr_ff_mux_state_427_13_g590/data4 , 
    \scr_ff_mux_state_427_13_g578/data3 , \scr_ff_mux_state_427_13_g578/data4 , 
    \scr_ff_mux_state_427_13_g562/data3 , \scr_ff_mux_state_427_13_g562/data4 , 
    \scr_ff_mux_state_427_13_g550/data3 , \scr_ff_mux_state_427_13_g550/data4 , 
    \scr_ff_mux_state_427_13_g534/data3 , \scr_ff_mux_state_427_13_g534/data4 , 
    \scr_ff_mux_state_427_13_g522/data3 , \scr_ff_mux_state_427_13_g522/data4 , 
    \scr_ff_mux_state_427_13_g506/data3 , \scr_ff_mux_state_427_13_g506/data4 , 
    \scr_ff_mux_state_427_13_g494/data3 , \scr_ff_mux_state_427_13_g494/data4 , 
    \scr_ff_mux_state_427_13_g478/data3 , \scr_ff_mux_state_427_13_g478/data4 , 
    \scr_ff_mux_state_427_13_g466/data3 , \scr_ff_mux_state_427_13_g466/data4 , 
    \scr_ff_mux_state_427_13_g450/data3 , \scr_ff_mux_state_427_13_g450/data4 , 
    \scr_ff_mux_state_427_13_g438/data3 , \scr_ff_mux_state_427_13_g438/data4 , 
    \scr_ff_mux_state_427_13_g422/data3 , \scr_ff_mux_state_427_13_g422/data4 , 
    \scr_ff_mux_state_427_13_g410/data3 , \scr_ff_mux_state_427_13_g410/data4 , 
    \scr_ff_mux_state_427_13_g394/data3 , \scr_ff_mux_state_427_13_g394/data4 , 
    \scr_ff_mux_state_427_13_g382/data3 , \scr_ff_mux_state_427_13_g382/data4 , 
    \scr_ff_mux_state_427_13_g366/data3 , \scr_ff_mux_state_427_13_g366/data4 , 
    \scr_ff_mux_state_427_13_g354/data3 , \scr_ff_mux_state_427_13_g354/data4 , 
    \scr_ff_mux_state_427_13_g338/data3 , \scr_ff_mux_state_427_13_g338/data4 , 
    \scr_ff_mux_state_427_13_g326/data3 , \scr_ff_mux_state_427_13_g326/data4 ;
wire   [31:0] scram;
wire   [31:0] scr_out_p;
wire   [31:0] scr_in;
wire   [31:0] scr_out;
  assign \scr_ff_mux_state_427_13_g758/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g746/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g730/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g718/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g702/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g690/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g674/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g662/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g646/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g634/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g618/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g606/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g590/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g578/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g562/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g550/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g534/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g522/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g506/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g494/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g478/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g466/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g450/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g438/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g422/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g410/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g394/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g382/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g366/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g354/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g338/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g326/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g758/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g746/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g730/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g718/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g702/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g690/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g674/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g662/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g646/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g634/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g618/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g606/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g590/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g578/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g562/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g550/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g534/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g522/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g506/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g494/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g478/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g466/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g450/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g438/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g422/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g410/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g394/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g382/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g366/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g354/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g338/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g326/data3  = 1'b1;
  or \scr_ff_mux_state_427_13_g758/org (scr_out_p[16], 
    \scr_ff_mux_state_427_13_g758/w_0 , \scr_ff_mux_state_427_13_g758/w_1 , 
    \scr_ff_mux_state_427_13_g758/w_2 , \scr_ff_mux_state_427_13_g758/w_3 , 
    \scr_ff_mux_state_427_13_g758/w_4 );
  and \scr_ff_mux_state_427_13_g758/a_4 (\scr_ff_mux_state_427_13_g758/w_4 , set, 
    \scr_ff_mux_state_427_13_g758/data4 );
  and \scr_ff_mux_state_427_13_g758/a_3 (\scr_ff_mux_state_427_13_g758/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g758/data3 );
  and \scr_ff_mux_state_427_13_g758/a_2 (\scr_ff_mux_state_427_13_g758/w_2 , 
    n_391, scr_in[16]);
  and \scr_ff_mux_state_427_13_g758/a_1 (\scr_ff_mux_state_427_13_g758/w_1 , 
    n_390, n_347);
  and \scr_ff_mux_state_427_13_g758/a_0 (\scr_ff_mux_state_427_13_g758/w_0 , 
    n_389, scr_out[16]);
  or \scr_ff_mux_state_427_13_g746/org (scr_out_p[15], 
    \scr_ff_mux_state_427_13_g746/w_0 , \scr_ff_mux_state_427_13_g746/w_1 , 
    \scr_ff_mux_state_427_13_g746/w_2 , \scr_ff_mux_state_427_13_g746/w_3 , 
    \scr_ff_mux_state_427_13_g746/w_4 );
  and \scr_ff_mux_state_427_13_g746/a_4 (\scr_ff_mux_state_427_13_g746/w_4 , set, 
    \scr_ff_mux_state_427_13_g746/data4 );
  and \scr_ff_mux_state_427_13_g746/a_3 (\scr_ff_mux_state_427_13_g746/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g746/data3 );
  and \scr_ff_mux_state_427_13_g746/a_2 (\scr_ff_mux_state_427_13_g746/w_2 , 
    n_391, scr_in[15]);
  and \scr_ff_mux_state_427_13_g746/a_1 (\scr_ff_mux_state_427_13_g746/w_1 , 
    n_390, n_352);
  and \scr_ff_mux_state_427_13_g746/a_0 (\scr_ff_mux_state_427_13_g746/w_0 , 
    n_389, scr_out[15]);
  or \scr_ff_mux_state_427_13_g730/org (scr_out_p[26], 
    \scr_ff_mux_state_427_13_g730/w_0 , \scr_ff_mux_state_427_13_g730/w_1 , 
    \scr_ff_mux_state_427_13_g730/w_2 , \scr_ff_mux_state_427_13_g730/w_3 , 
    \scr_ff_mux_state_427_13_g730/w_4 );
  and \scr_ff_mux_state_427_13_g730/a_4 (\scr_ff_mux_state_427_13_g730/w_4 , set, 
    \scr_ff_mux_state_427_13_g730/data4 );
  and \scr_ff_mux_state_427_13_g730/a_3 (\scr_ff_mux_state_427_13_g730/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g730/data3 );
  and \scr_ff_mux_state_427_13_g730/a_2 (\scr_ff_mux_state_427_13_g730/w_2 , 
    n_391, scr_in[26]);
  and \scr_ff_mux_state_427_13_g730/a_1 (\scr_ff_mux_state_427_13_g730/w_1 , 
    n_390, n_286);
  and \scr_ff_mux_state_427_13_g730/a_0 (\scr_ff_mux_state_427_13_g730/w_0 , 
    n_389, scr_out[26]);
  or \scr_ff_mux_state_427_13_g718/org (scr_out_p[27], 
    \scr_ff_mux_state_427_13_g718/w_0 , \scr_ff_mux_state_427_13_g718/w_1 , 
    \scr_ff_mux_state_427_13_g718/w_2 , \scr_ff_mux_state_427_13_g718/w_3 , 
    \scr_ff_mux_state_427_13_g718/w_4 );
  and \scr_ff_mux_state_427_13_g718/a_4 (\scr_ff_mux_state_427_13_g718/w_4 , set, 
    \scr_ff_mux_state_427_13_g718/data4 );
  and \scr_ff_mux_state_427_13_g718/a_3 (\scr_ff_mux_state_427_13_g718/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g718/data3 );
  and \scr_ff_mux_state_427_13_g718/a_2 (\scr_ff_mux_state_427_13_g718/w_2 , 
    n_391, scr_in[27]);
  and \scr_ff_mux_state_427_13_g718/a_1 (\scr_ff_mux_state_427_13_g718/w_1 , 
    n_390, n_282);
  and \scr_ff_mux_state_427_13_g718/a_0 (\scr_ff_mux_state_427_13_g718/w_0 , 
    n_389, scr_out[27]);
  or \scr_ff_mux_state_427_13_g702/org (scr_out_p[28], 
    \scr_ff_mux_state_427_13_g702/w_0 , \scr_ff_mux_state_427_13_g702/w_1 , 
    \scr_ff_mux_state_427_13_g702/w_2 , \scr_ff_mux_state_427_13_g702/w_3 , 
    \scr_ff_mux_state_427_13_g702/w_4 );
  and \scr_ff_mux_state_427_13_g702/a_4 (\scr_ff_mux_state_427_13_g702/w_4 , set, 
    \scr_ff_mux_state_427_13_g702/data4 );
  and \scr_ff_mux_state_427_13_g702/a_3 (\scr_ff_mux_state_427_13_g702/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g702/data3 );
  and \scr_ff_mux_state_427_13_g702/a_2 (\scr_ff_mux_state_427_13_g702/w_2 , 
    n_391, scr_in[28]);
  and \scr_ff_mux_state_427_13_g702/a_1 (\scr_ff_mux_state_427_13_g702/w_1 , 
    n_390, n_278);
  and \scr_ff_mux_state_427_13_g702/a_0 (\scr_ff_mux_state_427_13_g702/w_0 , 
    n_389, scr_out[28]);
  or \scr_ff_mux_state_427_13_g690/org (scr_out_p[29], 
    \scr_ff_mux_state_427_13_g690/w_0 , \scr_ff_mux_state_427_13_g690/w_1 , 
    \scr_ff_mux_state_427_13_g690/w_2 , \scr_ff_mux_state_427_13_g690/w_3 , 
    \scr_ff_mux_state_427_13_g690/w_4 );
  and \scr_ff_mux_state_427_13_g690/a_4 (\scr_ff_mux_state_427_13_g690/w_4 , set, 
    \scr_ff_mux_state_427_13_g690/data4 );
  and \scr_ff_mux_state_427_13_g690/a_3 (\scr_ff_mux_state_427_13_g690/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g690/data3 );
  and \scr_ff_mux_state_427_13_g690/a_2 (\scr_ff_mux_state_427_13_g690/w_2 , 
    n_391, scr_in[29]);
  and \scr_ff_mux_state_427_13_g690/a_1 (\scr_ff_mux_state_427_13_g690/w_1 , 
    n_390, n_275);
  and \scr_ff_mux_state_427_13_g690/a_0 (\scr_ff_mux_state_427_13_g690/w_0 , 
    n_389, scr_out[29]);
  or \scr_ff_mux_state_427_13_g674/org (scr_out_p[9], 
    \scr_ff_mux_state_427_13_g674/w_0 , \scr_ff_mux_state_427_13_g674/w_1 , 
    \scr_ff_mux_state_427_13_g674/w_2 , \scr_ff_mux_state_427_13_g674/w_3 , 
    \scr_ff_mux_state_427_13_g674/w_4 );
  and \scr_ff_mux_state_427_13_g674/a_4 (\scr_ff_mux_state_427_13_g674/w_4 , set, 
    \scr_ff_mux_state_427_13_g674/data4 );
  and \scr_ff_mux_state_427_13_g674/a_3 (\scr_ff_mux_state_427_13_g674/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g674/data3 );
  and \scr_ff_mux_state_427_13_g674/a_2 (\scr_ff_mux_state_427_13_g674/w_2 , 
    n_391, scr_in[9]);
  and \scr_ff_mux_state_427_13_g674/a_1 (\scr_ff_mux_state_427_13_g674/w_1 , 
    n_390, scram[9]);
  and \scr_ff_mux_state_427_13_g674/a_0 (\scr_ff_mux_state_427_13_g674/w_0 , 
    n_389, scr_out[9]);
  or \scr_ff_mux_state_427_13_g662/org (scr_out_p[10], 
    \scr_ff_mux_state_427_13_g662/w_0 , \scr_ff_mux_state_427_13_g662/w_1 , 
    \scr_ff_mux_state_427_13_g662/w_2 , \scr_ff_mux_state_427_13_g662/w_3 , 
    \scr_ff_mux_state_427_13_g662/w_4 );
  and \scr_ff_mux_state_427_13_g662/a_4 (\scr_ff_mux_state_427_13_g662/w_4 , set, 
    \scr_ff_mux_state_427_13_g662/data4 );
  and \scr_ff_mux_state_427_13_g662/a_3 (\scr_ff_mux_state_427_13_g662/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g662/data3 );
  and \scr_ff_mux_state_427_13_g662/a_2 (\scr_ff_mux_state_427_13_g662/w_2 , 
    n_391, scr_in[10]);
  and \scr_ff_mux_state_427_13_g662/a_1 (\scr_ff_mux_state_427_13_g662/w_1 , 
    n_390, scram[10]);
  and \scr_ff_mux_state_427_13_g662/a_0 (\scr_ff_mux_state_427_13_g662/w_0 , 
    n_389, scr_out[10]);
  or \scr_ff_mux_state_427_13_g646/org (scr_out_p[11], 
    \scr_ff_mux_state_427_13_g646/w_0 , \scr_ff_mux_state_427_13_g646/w_1 , 
    \scr_ff_mux_state_427_13_g646/w_2 , \scr_ff_mux_state_427_13_g646/w_3 , 
    \scr_ff_mux_state_427_13_g646/w_4 );
  and \scr_ff_mux_state_427_13_g646/a_4 (\scr_ff_mux_state_427_13_g646/w_4 , set, 
    \scr_ff_mux_state_427_13_g646/data4 );
  and \scr_ff_mux_state_427_13_g646/a_3 (\scr_ff_mux_state_427_13_g646/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g646/data3 );
  and \scr_ff_mux_state_427_13_g646/a_2 (\scr_ff_mux_state_427_13_g646/w_2 , 
    n_391, scr_in[11]);
  and \scr_ff_mux_state_427_13_g646/a_1 (\scr_ff_mux_state_427_13_g646/w_1 , 
    n_390, scram[11]);
  and \scr_ff_mux_state_427_13_g646/a_0 (\scr_ff_mux_state_427_13_g646/w_0 , 
    n_389, scr_out[11]);
  or \scr_ff_mux_state_427_13_g634/org (scr_out_p[12], 
    \scr_ff_mux_state_427_13_g634/w_0 , \scr_ff_mux_state_427_13_g634/w_1 , 
    \scr_ff_mux_state_427_13_g634/w_2 , \scr_ff_mux_state_427_13_g634/w_3 , 
    \scr_ff_mux_state_427_13_g634/w_4 );
  and \scr_ff_mux_state_427_13_g634/a_4 (\scr_ff_mux_state_427_13_g634/w_4 , set, 
    \scr_ff_mux_state_427_13_g634/data4 );
  and \scr_ff_mux_state_427_13_g634/a_3 (\scr_ff_mux_state_427_13_g634/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g634/data3 );
  and \scr_ff_mux_state_427_13_g634/a_2 (\scr_ff_mux_state_427_13_g634/w_2 , 
    n_391, scr_in[12]);
  and \scr_ff_mux_state_427_13_g634/a_1 (\scr_ff_mux_state_427_13_g634/w_1 , 
    n_390, n_367);
  and \scr_ff_mux_state_427_13_g634/a_0 (\scr_ff_mux_state_427_13_g634/w_0 , 
    n_389, scr_out[12]);
  or \scr_ff_mux_state_427_13_g618/org (scr_out_p[30], 
    \scr_ff_mux_state_427_13_g618/w_0 , \scr_ff_mux_state_427_13_g618/w_1 , 
    \scr_ff_mux_state_427_13_g618/w_2 , \scr_ff_mux_state_427_13_g618/w_3 , 
    \scr_ff_mux_state_427_13_g618/w_4 );
  and \scr_ff_mux_state_427_13_g618/a_4 (\scr_ff_mux_state_427_13_g618/w_4 , set, 
    \scr_ff_mux_state_427_13_g618/data4 );
  and \scr_ff_mux_state_427_13_g618/a_3 (\scr_ff_mux_state_427_13_g618/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g618/data3 );
  and \scr_ff_mux_state_427_13_g618/a_2 (\scr_ff_mux_state_427_13_g618/w_2 , 
    n_391, scr_in[30]);
  and \scr_ff_mux_state_427_13_g618/a_1 (\scr_ff_mux_state_427_13_g618/w_1 , 
    n_390, n_272);
  and \scr_ff_mux_state_427_13_g618/a_0 (\scr_ff_mux_state_427_13_g618/w_0 , 
    n_389, scr_out[30]);
  or \scr_ff_mux_state_427_13_g606/org (scr_out_p[13], 
    \scr_ff_mux_state_427_13_g606/w_0 , \scr_ff_mux_state_427_13_g606/w_1 , 
    \scr_ff_mux_state_427_13_g606/w_2 , \scr_ff_mux_state_427_13_g606/w_3 , 
    \scr_ff_mux_state_427_13_g606/w_4 );
  and \scr_ff_mux_state_427_13_g606/a_4 (\scr_ff_mux_state_427_13_g606/w_4 , set, 
    \scr_ff_mux_state_427_13_g606/data4 );
  and \scr_ff_mux_state_427_13_g606/a_3 (\scr_ff_mux_state_427_13_g606/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g606/data3 );
  and \scr_ff_mux_state_427_13_g606/a_2 (\scr_ff_mux_state_427_13_g606/w_2 , 
    n_391, scr_in[13]);
  and \scr_ff_mux_state_427_13_g606/a_1 (\scr_ff_mux_state_427_13_g606/w_1 , 
    n_390, n_362);
  and \scr_ff_mux_state_427_13_g606/a_0 (\scr_ff_mux_state_427_13_g606/w_0 , 
    n_389, scr_out[13]);
  or \scr_ff_mux_state_427_13_g590/org (scr_out_p[14], 
    \scr_ff_mux_state_427_13_g590/w_0 , \scr_ff_mux_state_427_13_g590/w_1 , 
    \scr_ff_mux_state_427_13_g590/w_2 , \scr_ff_mux_state_427_13_g590/w_3 , 
    \scr_ff_mux_state_427_13_g590/w_4 );
  and \scr_ff_mux_state_427_13_g590/a_4 (\scr_ff_mux_state_427_13_g590/w_4 , set, 
    \scr_ff_mux_state_427_13_g590/data4 );
  and \scr_ff_mux_state_427_13_g590/a_3 (\scr_ff_mux_state_427_13_g590/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g590/data3 );
  and \scr_ff_mux_state_427_13_g590/a_2 (\scr_ff_mux_state_427_13_g590/w_2 , 
    n_391, scr_in[14]);
  and \scr_ff_mux_state_427_13_g590/a_1 (\scr_ff_mux_state_427_13_g590/w_1 , 
    n_390, n_357);
  and \scr_ff_mux_state_427_13_g590/a_0 (\scr_ff_mux_state_427_13_g590/w_0 , 
    n_389, scr_out[14]);
  or \scr_ff_mux_state_427_13_g578/org (scr_out_p[31], 
    \scr_ff_mux_state_427_13_g578/w_0 , \scr_ff_mux_state_427_13_g578/w_1 , 
    \scr_ff_mux_state_427_13_g578/w_2 , \scr_ff_mux_state_427_13_g578/w_3 , 
    \scr_ff_mux_state_427_13_g578/w_4 );
  and \scr_ff_mux_state_427_13_g578/a_4 (\scr_ff_mux_state_427_13_g578/w_4 , set, 
    \scr_ff_mux_state_427_13_g578/data4 );
  and \scr_ff_mux_state_427_13_g578/a_3 (\scr_ff_mux_state_427_13_g578/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g578/data3 );
  and \scr_ff_mux_state_427_13_g578/a_2 (\scr_ff_mux_state_427_13_g578/w_2 , 
    n_391, scr_in[31]);
  and \scr_ff_mux_state_427_13_g578/a_1 (\scr_ff_mux_state_427_13_g578/w_1 , 
    n_390, n_269);
  and \scr_ff_mux_state_427_13_g578/a_0 (\scr_ff_mux_state_427_13_g578/w_0 , 
    n_389, scr_out[31]);
  or \scr_ff_mux_state_427_13_g562/org (scr_out_p[23], 
    \scr_ff_mux_state_427_13_g562/w_0 , \scr_ff_mux_state_427_13_g562/w_1 , 
    \scr_ff_mux_state_427_13_g562/w_2 , \scr_ff_mux_state_427_13_g562/w_3 , 
    \scr_ff_mux_state_427_13_g562/w_4 );
  and \scr_ff_mux_state_427_13_g562/a_4 (\scr_ff_mux_state_427_13_g562/w_4 , set, 
    \scr_ff_mux_state_427_13_g562/data4 );
  and \scr_ff_mux_state_427_13_g562/a_3 (\scr_ff_mux_state_427_13_g562/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g562/data3 );
  and \scr_ff_mux_state_427_13_g562/a_2 (\scr_ff_mux_state_427_13_g562/w_2 , 
    n_391, scr_in[23]);
  and \scr_ff_mux_state_427_13_g562/a_1 (\scr_ff_mux_state_427_13_g562/w_1 , 
    n_390, n_302);
  and \scr_ff_mux_state_427_13_g562/a_0 (\scr_ff_mux_state_427_13_g562/w_0 , 
    n_389, scr_out[23]);
  or \scr_ff_mux_state_427_13_g550/org (scr_out_p[24], 
    \scr_ff_mux_state_427_13_g550/w_0 , \scr_ff_mux_state_427_13_g550/w_1 , 
    \scr_ff_mux_state_427_13_g550/w_2 , \scr_ff_mux_state_427_13_g550/w_3 , 
    \scr_ff_mux_state_427_13_g550/w_4 );
  and \scr_ff_mux_state_427_13_g550/a_4 (\scr_ff_mux_state_427_13_g550/w_4 , set, 
    \scr_ff_mux_state_427_13_g550/data4 );
  and \scr_ff_mux_state_427_13_g550/a_3 (\scr_ff_mux_state_427_13_g550/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g550/data3 );
  and \scr_ff_mux_state_427_13_g550/a_2 (\scr_ff_mux_state_427_13_g550/w_2 , 
    n_391, scr_in[24]);
  and \scr_ff_mux_state_427_13_g550/a_1 (\scr_ff_mux_state_427_13_g550/w_1 , 
    n_390, n_296);
  and \scr_ff_mux_state_427_13_g550/a_0 (\scr_ff_mux_state_427_13_g550/w_0 , 
    n_389, scr_out[24]);
  or \scr_ff_mux_state_427_13_g534/org (scr_out_p[8], 
    \scr_ff_mux_state_427_13_g534/w_0 , \scr_ff_mux_state_427_13_g534/w_1 , 
    \scr_ff_mux_state_427_13_g534/w_2 , \scr_ff_mux_state_427_13_g534/w_3 , 
    \scr_ff_mux_state_427_13_g534/w_4 );
  and \scr_ff_mux_state_427_13_g534/a_4 (\scr_ff_mux_state_427_13_g534/w_4 , set, 
    \scr_ff_mux_state_427_13_g534/data4 );
  and \scr_ff_mux_state_427_13_g534/a_3 (\scr_ff_mux_state_427_13_g534/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g534/data3 );
  and \scr_ff_mux_state_427_13_g534/a_2 (\scr_ff_mux_state_427_13_g534/w_2 , 
    n_391, scr_in[8]);
  and \scr_ff_mux_state_427_13_g534/a_1 (\scr_ff_mux_state_427_13_g534/w_1 , 
    n_390, n_171);
  and \scr_ff_mux_state_427_13_g534/a_0 (\scr_ff_mux_state_427_13_g534/w_0 , 
    n_389, scr_out[8]);
  or \scr_ff_mux_state_427_13_g522/org (scr_out_p[25], 
    \scr_ff_mux_state_427_13_g522/w_0 , \scr_ff_mux_state_427_13_g522/w_1 , 
    \scr_ff_mux_state_427_13_g522/w_2 , \scr_ff_mux_state_427_13_g522/w_3 , 
    \scr_ff_mux_state_427_13_g522/w_4 );
  and \scr_ff_mux_state_427_13_g522/a_4 (\scr_ff_mux_state_427_13_g522/w_4 , set, 
    \scr_ff_mux_state_427_13_g522/data4 );
  and \scr_ff_mux_state_427_13_g522/a_3 (\scr_ff_mux_state_427_13_g522/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g522/data3 );
  and \scr_ff_mux_state_427_13_g522/a_2 (\scr_ff_mux_state_427_13_g522/w_2 , 
    n_391, scr_in[25]);
  and \scr_ff_mux_state_427_13_g522/a_1 (\scr_ff_mux_state_427_13_g522/w_1 , 
    n_390, n_291);
  and \scr_ff_mux_state_427_13_g522/a_0 (\scr_ff_mux_state_427_13_g522/w_0 , 
    n_389, scr_out[25]);
  or \scr_ff_mux_state_427_13_g506/org (scr_out_p[7], 
    \scr_ff_mux_state_427_13_g506/w_0 , \scr_ff_mux_state_427_13_g506/w_1 , 
    \scr_ff_mux_state_427_13_g506/w_2 , \scr_ff_mux_state_427_13_g506/w_3 , 
    \scr_ff_mux_state_427_13_g506/w_4 );
  and \scr_ff_mux_state_427_13_g506/a_4 (\scr_ff_mux_state_427_13_g506/w_4 , set, 
    \scr_ff_mux_state_427_13_g506/data4 );
  and \scr_ff_mux_state_427_13_g506/a_3 (\scr_ff_mux_state_427_13_g506/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g506/data3 );
  and \scr_ff_mux_state_427_13_g506/a_2 (\scr_ff_mux_state_427_13_g506/w_2 , 
    n_391, scr_in[7]);
  and \scr_ff_mux_state_427_13_g506/a_1 (\scr_ff_mux_state_427_13_g506/w_1 , 
    n_390, n_178);
  and \scr_ff_mux_state_427_13_g506/a_0 (\scr_ff_mux_state_427_13_g506/w_0 , 
    n_389, scr_out[7]);
  or \scr_ff_mux_state_427_13_g494/org (scr_out_p[17], 
    \scr_ff_mux_state_427_13_g494/w_0 , \scr_ff_mux_state_427_13_g494/w_1 , 
    \scr_ff_mux_state_427_13_g494/w_2 , \scr_ff_mux_state_427_13_g494/w_3 , 
    \scr_ff_mux_state_427_13_g494/w_4 );
  and \scr_ff_mux_state_427_13_g494/a_4 (\scr_ff_mux_state_427_13_g494/w_4 , set, 
    \scr_ff_mux_state_427_13_g494/data4 );
  and \scr_ff_mux_state_427_13_g494/a_3 (\scr_ff_mux_state_427_13_g494/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g494/data3 );
  and \scr_ff_mux_state_427_13_g494/a_2 (\scr_ff_mux_state_427_13_g494/w_2 , 
    n_391, scr_in[17]);
  and \scr_ff_mux_state_427_13_g494/a_1 (\scr_ff_mux_state_427_13_g494/w_1 , 
    n_390, n_343);
  and \scr_ff_mux_state_427_13_g494/a_0 (\scr_ff_mux_state_427_13_g494/w_0 , 
    n_389, scr_out[17]);
  or \scr_ff_mux_state_427_13_g478/org (scr_out_p[18], 
    \scr_ff_mux_state_427_13_g478/w_0 , \scr_ff_mux_state_427_13_g478/w_1 , 
    \scr_ff_mux_state_427_13_g478/w_2 , \scr_ff_mux_state_427_13_g478/w_3 , 
    \scr_ff_mux_state_427_13_g478/w_4 );
  and \scr_ff_mux_state_427_13_g478/a_4 (\scr_ff_mux_state_427_13_g478/w_4 , set, 
    \scr_ff_mux_state_427_13_g478/data4 );
  and \scr_ff_mux_state_427_13_g478/a_3 (\scr_ff_mux_state_427_13_g478/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g478/data3 );
  and \scr_ff_mux_state_427_13_g478/a_2 (\scr_ff_mux_state_427_13_g478/w_2 , 
    n_391, scr_in[18]);
  and \scr_ff_mux_state_427_13_g478/a_1 (\scr_ff_mux_state_427_13_g478/w_1 , 
    n_390, n_336);
  and \scr_ff_mux_state_427_13_g478/a_0 (\scr_ff_mux_state_427_13_g478/w_0 , 
    n_389, scr_out[18]);
  or \scr_ff_mux_state_427_13_g466/org (scr_out_p[22], 
    \scr_ff_mux_state_427_13_g466/w_0 , \scr_ff_mux_state_427_13_g466/w_1 , 
    \scr_ff_mux_state_427_13_g466/w_2 , \scr_ff_mux_state_427_13_g466/w_3 , 
    \scr_ff_mux_state_427_13_g466/w_4 );
  and \scr_ff_mux_state_427_13_g466/a_4 (\scr_ff_mux_state_427_13_g466/w_4 , set, 
    \scr_ff_mux_state_427_13_g466/data4 );
  and \scr_ff_mux_state_427_13_g466/a_3 (\scr_ff_mux_state_427_13_g466/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g466/data3 );
  and \scr_ff_mux_state_427_13_g466/a_2 (\scr_ff_mux_state_427_13_g466/w_2 , 
    n_391, scr_in[22]);
  and \scr_ff_mux_state_427_13_g466/a_1 (\scr_ff_mux_state_427_13_g466/w_1 , 
    n_390, n_309);
  and \scr_ff_mux_state_427_13_g466/a_0 (\scr_ff_mux_state_427_13_g466/w_0 , 
    n_389, scr_out[22]);
  or \scr_ff_mux_state_427_13_g450/org (scr_out_p[4], 
    \scr_ff_mux_state_427_13_g450/w_0 , \scr_ff_mux_state_427_13_g450/w_1 , 
    \scr_ff_mux_state_427_13_g450/w_2 , \scr_ff_mux_state_427_13_g450/w_3 , 
    \scr_ff_mux_state_427_13_g450/w_4 );
  and \scr_ff_mux_state_427_13_g450/a_4 (\scr_ff_mux_state_427_13_g450/w_4 , set, 
    \scr_ff_mux_state_427_13_g450/data4 );
  and \scr_ff_mux_state_427_13_g450/a_3 (\scr_ff_mux_state_427_13_g450/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g450/data3 );
  and \scr_ff_mux_state_427_13_g450/a_2 (\scr_ff_mux_state_427_13_g450/w_2 , 
    n_391, scr_in[4]);
  and \scr_ff_mux_state_427_13_g450/a_1 (\scr_ff_mux_state_427_13_g450/w_1 , 
    n_390, n_199);
  and \scr_ff_mux_state_427_13_g450/a_0 (\scr_ff_mux_state_427_13_g450/w_0 , 
    n_389, scr_out[4]);
  or \scr_ff_mux_state_427_13_g438/org (scr_out_p[5], 
    \scr_ff_mux_state_427_13_g438/w_0 , \scr_ff_mux_state_427_13_g438/w_1 , 
    \scr_ff_mux_state_427_13_g438/w_2 , \scr_ff_mux_state_427_13_g438/w_3 , 
    \scr_ff_mux_state_427_13_g438/w_4 );
  and \scr_ff_mux_state_427_13_g438/a_4 (\scr_ff_mux_state_427_13_g438/w_4 , set, 
    \scr_ff_mux_state_427_13_g438/data4 );
  and \scr_ff_mux_state_427_13_g438/a_3 (\scr_ff_mux_state_427_13_g438/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g438/data3 );
  and \scr_ff_mux_state_427_13_g438/a_2 (\scr_ff_mux_state_427_13_g438/w_2 , 
    n_391, scr_in[5]);
  and \scr_ff_mux_state_427_13_g438/a_1 (\scr_ff_mux_state_427_13_g438/w_1 , 
    n_390, n_192);
  and \scr_ff_mux_state_427_13_g438/a_0 (\scr_ff_mux_state_427_13_g438/w_0 , 
    n_389, scr_out[5]);
  or \scr_ff_mux_state_427_13_g422/org (scr_out_p[6], 
    \scr_ff_mux_state_427_13_g422/w_0 , \scr_ff_mux_state_427_13_g422/w_1 , 
    \scr_ff_mux_state_427_13_g422/w_2 , \scr_ff_mux_state_427_13_g422/w_3 , 
    \scr_ff_mux_state_427_13_g422/w_4 );
  and \scr_ff_mux_state_427_13_g422/a_4 (\scr_ff_mux_state_427_13_g422/w_4 , set, 
    \scr_ff_mux_state_427_13_g422/data4 );
  and \scr_ff_mux_state_427_13_g422/a_3 (\scr_ff_mux_state_427_13_g422/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g422/data3 );
  and \scr_ff_mux_state_427_13_g422/a_2 (\scr_ff_mux_state_427_13_g422/w_2 , 
    n_391, scr_in[6]);
  and \scr_ff_mux_state_427_13_g422/a_1 (\scr_ff_mux_state_427_13_g422/w_1 , 
    n_390, n_185);
  and \scr_ff_mux_state_427_13_g422/a_0 (\scr_ff_mux_state_427_13_g422/w_0 , 
    n_389, scr_out[6]);
  or \scr_ff_mux_state_427_13_g410/org (scr_out_p[21], 
    \scr_ff_mux_state_427_13_g410/w_0 , \scr_ff_mux_state_427_13_g410/w_1 , 
    \scr_ff_mux_state_427_13_g410/w_2 , \scr_ff_mux_state_427_13_g410/w_3 , 
    \scr_ff_mux_state_427_13_g410/w_4 );
  and \scr_ff_mux_state_427_13_g410/a_4 (\scr_ff_mux_state_427_13_g410/w_4 , set, 
    \scr_ff_mux_state_427_13_g410/data4 );
  and \scr_ff_mux_state_427_13_g410/a_3 (\scr_ff_mux_state_427_13_g410/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g410/data3 );
  and \scr_ff_mux_state_427_13_g410/a_2 (\scr_ff_mux_state_427_13_g410/w_2 , 
    n_391, scr_in[21]);
  and \scr_ff_mux_state_427_13_g410/a_1 (\scr_ff_mux_state_427_13_g410/w_1 , 
    n_390, n_316);
  and \scr_ff_mux_state_427_13_g410/a_0 (\scr_ff_mux_state_427_13_g410/w_0 , 
    n_389, scr_out[21]);
  or \scr_ff_mux_state_427_13_g394/org (scr_out_p[3], 
    \scr_ff_mux_state_427_13_g394/w_0 , \scr_ff_mux_state_427_13_g394/w_1 , 
    \scr_ff_mux_state_427_13_g394/w_2 , \scr_ff_mux_state_427_13_g394/w_3 , 
    \scr_ff_mux_state_427_13_g394/w_4 );
  and \scr_ff_mux_state_427_13_g394/a_4 (\scr_ff_mux_state_427_13_g394/w_4 , set, 
    \scr_ff_mux_state_427_13_g394/data4 );
  and \scr_ff_mux_state_427_13_g394/a_3 (\scr_ff_mux_state_427_13_g394/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g394/data3 );
  and \scr_ff_mux_state_427_13_g394/a_2 (\scr_ff_mux_state_427_13_g394/w_2 , 
    n_391, scr_in[3]);
  and \scr_ff_mux_state_427_13_g394/a_1 (\scr_ff_mux_state_427_13_g394/w_1 , 
    n_390, n_81);
  and \scr_ff_mux_state_427_13_g394/a_0 (\scr_ff_mux_state_427_13_g394/w_0 , 
    n_389, scr_out[3]);
  or \scr_ff_mux_state_427_13_g382/org (scr_out_p[19], 
    \scr_ff_mux_state_427_13_g382/w_0 , \scr_ff_mux_state_427_13_g382/w_1 , 
    \scr_ff_mux_state_427_13_g382/w_2 , \scr_ff_mux_state_427_13_g382/w_3 , 
    \scr_ff_mux_state_427_13_g382/w_4 );
  and \scr_ff_mux_state_427_13_g382/a_4 (\scr_ff_mux_state_427_13_g382/w_4 , set, 
    \scr_ff_mux_state_427_13_g382/data4 );
  and \scr_ff_mux_state_427_13_g382/a_3 (\scr_ff_mux_state_427_13_g382/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g382/data3 );
  and \scr_ff_mux_state_427_13_g382/a_2 (\scr_ff_mux_state_427_13_g382/w_2 , 
    n_391, scr_in[19]);
  and \scr_ff_mux_state_427_13_g382/a_1 (\scr_ff_mux_state_427_13_g382/w_1 , 
    n_390, n_329);
  and \scr_ff_mux_state_427_13_g382/a_0 (\scr_ff_mux_state_427_13_g382/w_0 , 
    n_389, scr_out[19]);
  or \scr_ff_mux_state_427_13_g366/org (scr_out_p[20], 
    \scr_ff_mux_state_427_13_g366/w_0 , \scr_ff_mux_state_427_13_g366/w_1 , 
    \scr_ff_mux_state_427_13_g366/w_2 , \scr_ff_mux_state_427_13_g366/w_3 , 
    \scr_ff_mux_state_427_13_g366/w_4 );
  and \scr_ff_mux_state_427_13_g366/a_4 (\scr_ff_mux_state_427_13_g366/w_4 , set, 
    \scr_ff_mux_state_427_13_g366/data4 );
  and \scr_ff_mux_state_427_13_g366/a_3 (\scr_ff_mux_state_427_13_g366/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g366/data3 );
  and \scr_ff_mux_state_427_13_g366/a_2 (\scr_ff_mux_state_427_13_g366/w_2 , 
    n_391, scr_in[20]);
  and \scr_ff_mux_state_427_13_g366/a_1 (\scr_ff_mux_state_427_13_g366/w_1 , 
    n_390, n_322);
  and \scr_ff_mux_state_427_13_g366/a_0 (\scr_ff_mux_state_427_13_g366/w_0 , 
    n_389, scr_out[20]);
  or \scr_ff_mux_state_427_13_g354/org (scr_out_p[1], 
    \scr_ff_mux_state_427_13_g354/w_0 , \scr_ff_mux_state_427_13_g354/w_1 , 
    \scr_ff_mux_state_427_13_g354/w_2 , \scr_ff_mux_state_427_13_g354/w_3 , 
    \scr_ff_mux_state_427_13_g354/w_4 );
  and \scr_ff_mux_state_427_13_g354/a_4 (\scr_ff_mux_state_427_13_g354/w_4 , set, 
    \scr_ff_mux_state_427_13_g354/data4 );
  and \scr_ff_mux_state_427_13_g354/a_3 (\scr_ff_mux_state_427_13_g354/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g354/data3 );
  and \scr_ff_mux_state_427_13_g354/a_2 (\scr_ff_mux_state_427_13_g354/w_2 , 
    n_391, scr_in[1]);
  and \scr_ff_mux_state_427_13_g354/a_1 (\scr_ff_mux_state_427_13_g354/w_1 , 
    n_390, n_93);
  and \scr_ff_mux_state_427_13_g354/a_0 (\scr_ff_mux_state_427_13_g354/w_0 , 
    n_389, scr_out[1]);
  or \scr_ff_mux_state_427_13_g338/org (scr_out_p[2], 
    \scr_ff_mux_state_427_13_g338/w_0 , \scr_ff_mux_state_427_13_g338/w_1 , 
    \scr_ff_mux_state_427_13_g338/w_2 , \scr_ff_mux_state_427_13_g338/w_3 , 
    \scr_ff_mux_state_427_13_g338/w_4 );
  and \scr_ff_mux_state_427_13_g338/a_4 (\scr_ff_mux_state_427_13_g338/w_4 , set, 
    \scr_ff_mux_state_427_13_g338/data4 );
  and \scr_ff_mux_state_427_13_g338/a_3 (\scr_ff_mux_state_427_13_g338/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g338/data3 );
  and \scr_ff_mux_state_427_13_g338/a_2 (\scr_ff_mux_state_427_13_g338/w_2 , 
    n_391, scr_in[2]);
  and \scr_ff_mux_state_427_13_g338/a_1 (\scr_ff_mux_state_427_13_g338/w_1 , 
    n_390, n_87);
  and \scr_ff_mux_state_427_13_g338/a_0 (\scr_ff_mux_state_427_13_g338/w_0 , 
    n_389, scr_out[2]);
  or \scr_ff_mux_state_427_13_g326/org (scr_out_p[0], 
    \scr_ff_mux_state_427_13_g326/w_0 , \scr_ff_mux_state_427_13_g326/w_1 , 
    \scr_ff_mux_state_427_13_g326/w_2 , \scr_ff_mux_state_427_13_g326/w_3 , 
    \scr_ff_mux_state_427_13_g326/w_4 );
  and \scr_ff_mux_state_427_13_g326/a_4 (\scr_ff_mux_state_427_13_g326/w_4 , set, 
    \scr_ff_mux_state_427_13_g326/data4 );
  and \scr_ff_mux_state_427_13_g326/a_3 (\scr_ff_mux_state_427_13_g326/w_3 , 
    n_392, \scr_ff_mux_state_427_13_g326/data3 );
  and \scr_ff_mux_state_427_13_g326/a_2 (\scr_ff_mux_state_427_13_g326/w_2 , 
    n_391, scr_in[0]);
  and \scr_ff_mux_state_427_13_g326/a_1 (\scr_ff_mux_state_427_13_g326/w_1 , 
    n_390, a15);
  and \scr_ff_mux_state_427_13_g326/a_0 (\scr_ff_mux_state_427_13_g326/w_0 , 
    n_389, scr_out[0]);
  xor g10(\a10[0] , scr_out[25], scr_out[21]);
  xor g11(\a9[0] , scr_out[26], scr_out[22]);
  xor g12(\a8[0] , scr_out[27], scr_out[23]);
  xor g128(n_170, n_101, \a8[0] );
  xor g129(n_171, n_170, \a7[0] );
  xor g13(\a7[0] , scr_out[28], scr_out[24]);
  xor g136(n_177, n_75, \a9[0] );
  xor g137(n_178, n_177, \a8[0] );
  xor g14(\a6[0] , scr_out[29], scr_out[25]);
  xor g144(n_184, n_111, \a10[0] );
  xor g145(n_185, n_184, \a9[0] );
  xor g15(\a5[0] , scr_out[30], scr_out[26]);
  xor g152(n_191, n_87, \a11[0] );
  xor g153(n_192, n_191, \a10[0] );
  xor g16(\a4[0] , scr_out[31], scr_out[27]);
  xor g160(n_198, n_93, \a12[0] );
  xor g161(n_199, n_198, \a11[0] );
  xor g17(n_74, a15, \a12[0] );
  xor g172(n_209, n_84, \a5[0] );
  xor g173(scram[11], n_209, \a4[0] );
  xor g178(n_214, n_90, \a6[0] );
  xor g179(scram[10], n_214, \a5[0] );
  xor g18(n_75, n_74, \a11[0] );
  xor g184(n_219, n_96, \a7[0] );
  xor g185(scram[9], n_219, \a6[0] );
  xor g19(n_76, n_75, \a10[0] );
  xor g208(n_266, n_76, \a7[0] );
  xor g209(n_267, \a6[0] , \a5[0] );
  xor g210(n_268, scr_out[31], n_266);
  xor g211(n_269, n_267, n_268);
  xor g212(n_270, n_84, \a6[0] );
  xor g213(n_271, scr_out[30], scr_out[31]);
  xor g214(n_272, n_270, n_271);
  xor g215(n_273, n_90, \a7[0] );
  xor g216(n_274, scr_out[29], scr_out[30]);
  xor g217(n_275, n_273, n_274);
  xor g218(n_276, n_96, \a8[0] );
  xor g219(n_277, scr_out[28], scr_out[29]);
  xor g220(n_278, n_276, n_277);
  xor g221(n_279, n_101, \a9[0] );
  xor g222(n_280, \a4[0] , scr_out[28]);
  xor g223(n_281, scr_out[31], n_279);
  xor g224(n_282, n_280, n_281);
  xor g225(n_283, n_76, \a5[0] );
  xor g226(n_284, \a4[0] , scr_out[30]);
  xor g227(n_285, scr_out[31], n_283);
  xor g228(n_286, n_284, n_285);
  xor g229(n_287, n_111, \a11[0] );
  xor g232(n_290, n_287, n_267);
  xor g233(n_291, n_274, n_290);
  xor g234(n_292, n_88, \a7[0] );
  xor g235(n_293, \a6[0] , scr_out[28]);
  xor g236(n_294, scr_out[29], scr_out[31]);
  xor g237(n_295, n_292, n_293);
  xor g238(n_296, n_294, n_295);
  xor g239(n_297, n_94, \a8[0] );
  xor g24(n_80, a15, \a13[0] );
  xor g240(n_298, \a7[0] , \a4[0] );
  xor g241(n_299, scr_out[28], scr_out[30]);
  xor g242(n_300, scr_out[31], n_297);
  xor g243(n_301, n_298, n_299);
  xor g244(n_302, n_300, n_301);
  xor g245(n_303, n_93, \a9[0] );
  xor g246(n_304, \a8[0] , \a5[0] );
  xor g247(n_305, \a4[0] , scr_out[29]);
  xor g249(n_307, n_303, n_304);
  xor g25(n_81, n_80, \a12[0] );
  xor g250(n_308, n_305, n_271);
  xor g251(n_309, n_307, n_308);
  xor g252(n_310, a15, \a10[0] );
  xor g253(n_311, \a9[0] , \a6[0] );
  xor g254(n_312, \a5[0] , scr_out[28]);
  xor g256(n_314, n_310, n_311);
  xor g257(n_315, n_312, n_274);
  xor g258(n_316, n_314, n_315);
  xor g259(n_317, \a11[0] , \a10[0] );
  xor g260(n_318, \a7[0] , \a6[0] );
  xor g262(n_320, scr_out[29], n_317);
  xor g263(n_321, n_318, n_280);
  xor g264(n_322, n_320, n_321);
  xor g265(n_323, \a12[0] , \a11[0] );
  xor g266(n_324, \a8[0] , \a7[0] );
  xor g267(n_325, \a5[0] , \a4[0] );
  xor g268(n_326, scr_out[28], scr_out[31]);
  xor g269(n_327, n_323, n_324);
  xor g270(n_328, n_325, n_326);
  xor g271(n_329, n_327, n_328);
  xor g272(n_330, n_111, \a9[0] );
  xor g273(n_331, \a8[0] , \a6[0] );
  xor g276(n_334, n_330, n_331);
  xor g277(n_335, n_325, n_271);
  xor g278(n_336, n_334, n_335);
  xor g279(n_337, n_87, \a10[0] );
  xor g280(n_338, \a9[0] , \a7[0] );
  xor g283(n_341, n_337, n_338);
  xor g284(n_342, n_267, n_274);
  xor g285(n_343, n_341, n_342);
  xor g286(n_344, n_171, \a6[0] );
  xor g288(n_346, scr_out[31], n_344);
  xor g289(n_347, n_277, n_346);
  xor g290(n_348, n_178, \a7[0] );
  xor g293(n_351, n_348, n_280);
  xor g294(n_352, n_271, n_351);
  xor g295(n_353, n_185, \a8[0] );
  xor g298(n_356, n_353, n_325);
  xor g299(n_357, n_274, n_356);
  xor g300(n_358, n_192, \a9[0] );
  xor g303(n_361, n_358, n_267);
  xor g304(n_362, n_277, n_361);
  xor g305(n_363, n_199, \a10[0] );
  xor g308(n_366, n_363, n_318);
  xor g309(n_367, n_280, n_366);
  xor g311(n_369, scr_out[20], scr_out[16]);
  xor g312(a15, n_294, n_369);
  xor g313(n_370, n_81, \a11[0] );
  xor g315(n_84, n_370, n_324);
  xor g32(n_87, \a14[0] , \a13[0] );
  xor g33(n_88, n_87, \a12[0] );
  xor g34(n_89, n_88, \a9[0] );
  xor g35(n_90, n_89, \a8[0] );
  xor g39(n_93, a15, \a14[0] );
  xor g4(n_72, scr_out[30], scr_out[21]);
  xor g40(n_94, n_93, \a13[0] );
  xor g41(n_95, n_94, \a10[0] );
  xor g42(n_96, n_95, \a9[0] );
  xor g47(n_100, n_93, \a11[0] );
  xor g48(n_101, n_100, \a10[0] );
  xor g5(\a14[0] , n_72, scr_out[17]);
  xor g6(n_73, scr_out[31], scr_out[22]);
  xor g60(n_111, \a13[0] , \a12[0] );
  xor g7(\a13[0] , n_73, scr_out[18]);
  xor g8(\a12[0] , scr_out[23], scr_out[19]);
  xor g9(\a11[0] , scr_out[24], scr_out[20]);
  nor g22(n_389, scr_run, set, scr_init, reset);
  not g810(n_1118, reset);
  not g811(n_1119, scr_init);
  not g812(n_1120, scr_run);
  nor g813(n_390, scr_init, n_1120, reset, set);
  nor g814(n_391, n_1119, reset, set);
  nor g815(n_392, n_1118, set);
endmodule

