//
// Conformal-LEC: Version 11.10-d208 (10-Mar-2012) (64 bit executable)
//
module top(scr_out, scr_in, scr_init, scr_run, clk, reset, scr_out_p, set);
input  scr_init, scr_run, clk, reset, set;
input   [31:0] scr_out;
input   [31:0] scr_in;
output  [31:0] scr_out_p;
wire  \scr_ff_mux_state_427_13_g792/w_0 , \scr_ff_mux_state_427_13_g792/w_1 , 
    \scr_ff_mux_state_427_13_g792/w_2 , \scr_ff_mux_state_427_13_g792/w_3 , 
    \scr_ff_mux_state_427_13_g792/w_4 , \scr_ff_mux_state_427_13_g780/w_0 , 
    \scr_ff_mux_state_427_13_g780/w_1 , \scr_ff_mux_state_427_13_g780/w_2 , 
    \scr_ff_mux_state_427_13_g780/w_3 , \scr_ff_mux_state_427_13_g780/w_4 , 
    \scr_ff_mux_state_427_13_g764/w_0 , \scr_ff_mux_state_427_13_g764/w_1 , 
    \scr_ff_mux_state_427_13_g764/w_2 , \scr_ff_mux_state_427_13_g764/w_3 , 
    \scr_ff_mux_state_427_13_g764/w_4 , \scr_ff_mux_state_427_13_g752/w_0 , 
    \scr_ff_mux_state_427_13_g752/w_1 , \scr_ff_mux_state_427_13_g752/w_2 , 
    \scr_ff_mux_state_427_13_g752/w_3 , \scr_ff_mux_state_427_13_g752/w_4 , 
    \scr_ff_mux_state_427_13_g736/w_0 , \scr_ff_mux_state_427_13_g736/w_1 , 
    \scr_ff_mux_state_427_13_g736/w_2 , \scr_ff_mux_state_427_13_g736/w_3 , 
    \scr_ff_mux_state_427_13_g736/w_4 , \scr_ff_mux_state_427_13_g724/w_0 , 
    \scr_ff_mux_state_427_13_g724/w_1 , \scr_ff_mux_state_427_13_g724/w_2 , 
    \scr_ff_mux_state_427_13_g724/w_3 , \scr_ff_mux_state_427_13_g724/w_4 , 
    \scr_ff_mux_state_427_13_g708/w_0 , \scr_ff_mux_state_427_13_g708/w_1 , 
    \scr_ff_mux_state_427_13_g708/w_2 , \scr_ff_mux_state_427_13_g708/w_3 , 
    \scr_ff_mux_state_427_13_g708/w_4 , \scr_ff_mux_state_427_13_g696/w_0 , 
    \scr_ff_mux_state_427_13_g696/w_1 , \scr_ff_mux_state_427_13_g696/w_2 , 
    \scr_ff_mux_state_427_13_g696/w_3 , \scr_ff_mux_state_427_13_g696/w_4 , 
    \scr_ff_mux_state_427_13_g680/w_0 , \scr_ff_mux_state_427_13_g680/w_1 , 
    \scr_ff_mux_state_427_13_g680/w_2 , \scr_ff_mux_state_427_13_g680/w_3 , 
    \scr_ff_mux_state_427_13_g680/w_4 , \scr_ff_mux_state_427_13_g668/w_0 , 
    \scr_ff_mux_state_427_13_g668/w_1 , \scr_ff_mux_state_427_13_g668/w_2 , 
    \scr_ff_mux_state_427_13_g668/w_3 , \scr_ff_mux_state_427_13_g668/w_4 , 
    \scr_ff_mux_state_427_13_g652/w_0 , \scr_ff_mux_state_427_13_g652/w_1 , 
    \scr_ff_mux_state_427_13_g652/w_2 , \scr_ff_mux_state_427_13_g652/w_3 , 
    \scr_ff_mux_state_427_13_g652/w_4 , \scr_ff_mux_state_427_13_g640/w_0 , 
    \scr_ff_mux_state_427_13_g640/w_1 , \scr_ff_mux_state_427_13_g640/w_2 , 
    \scr_ff_mux_state_427_13_g640/w_3 , \scr_ff_mux_state_427_13_g640/w_4 , 
    \scr_ff_mux_state_427_13_g624/w_0 , \scr_ff_mux_state_427_13_g624/w_1 , 
    \scr_ff_mux_state_427_13_g624/w_2 , \scr_ff_mux_state_427_13_g624/w_3 , 
    \scr_ff_mux_state_427_13_g624/w_4 , \scr_ff_mux_state_427_13_g612/w_0 , 
    \scr_ff_mux_state_427_13_g612/w_1 , \scr_ff_mux_state_427_13_g612/w_2 , 
    \scr_ff_mux_state_427_13_g612/w_3 , \scr_ff_mux_state_427_13_g612/w_4 , 
    \scr_ff_mux_state_427_13_g596/w_0 , \scr_ff_mux_state_427_13_g596/w_1 , 
    \scr_ff_mux_state_427_13_g596/w_2 , \scr_ff_mux_state_427_13_g596/w_3 , 
    \scr_ff_mux_state_427_13_g596/w_4 , \scr_ff_mux_state_427_13_g584/w_0 , 
    \scr_ff_mux_state_427_13_g584/w_1 , \scr_ff_mux_state_427_13_g584/w_2 , 
    \scr_ff_mux_state_427_13_g584/w_3 , \scr_ff_mux_state_427_13_g584/w_4 , 
    \scr_ff_mux_state_427_13_g568/w_0 , \scr_ff_mux_state_427_13_g568/w_1 , 
    \scr_ff_mux_state_427_13_g568/w_2 , \scr_ff_mux_state_427_13_g568/w_3 , 
    \scr_ff_mux_state_427_13_g568/w_4 , \scr_ff_mux_state_427_13_g556/w_0 , 
    \scr_ff_mux_state_427_13_g556/w_1 , \scr_ff_mux_state_427_13_g556/w_2 , 
    \scr_ff_mux_state_427_13_g556/w_3 , \scr_ff_mux_state_427_13_g556/w_4 , 
    \scr_ff_mux_state_427_13_g540/w_0 , \scr_ff_mux_state_427_13_g540/w_1 , 
    \scr_ff_mux_state_427_13_g540/w_2 , \scr_ff_mux_state_427_13_g540/w_3 , 
    \scr_ff_mux_state_427_13_g540/w_4 , \scr_ff_mux_state_427_13_g528/w_0 , 
    \scr_ff_mux_state_427_13_g528/w_1 , \scr_ff_mux_state_427_13_g528/w_2 , 
    \scr_ff_mux_state_427_13_g528/w_3 , \scr_ff_mux_state_427_13_g528/w_4 , 
    \scr_ff_mux_state_427_13_g512/w_0 , \scr_ff_mux_state_427_13_g512/w_1 , 
    \scr_ff_mux_state_427_13_g512/w_2 , \scr_ff_mux_state_427_13_g512/w_3 , 
    \scr_ff_mux_state_427_13_g512/w_4 , \scr_ff_mux_state_427_13_g500/w_0 , 
    \scr_ff_mux_state_427_13_g500/w_1 , \scr_ff_mux_state_427_13_g500/w_2 , 
    \scr_ff_mux_state_427_13_g500/w_3 , \scr_ff_mux_state_427_13_g500/w_4 , 
    \scr_ff_mux_state_427_13_g484/w_0 , \scr_ff_mux_state_427_13_g484/w_1 , 
    \scr_ff_mux_state_427_13_g484/w_2 , \scr_ff_mux_state_427_13_g484/w_3 , 
    \scr_ff_mux_state_427_13_g484/w_4 , \scr_ff_mux_state_427_13_g472/w_0 , 
    \scr_ff_mux_state_427_13_g472/w_1 , \scr_ff_mux_state_427_13_g472/w_2 , 
    \scr_ff_mux_state_427_13_g472/w_3 , \scr_ff_mux_state_427_13_g472/w_4 , 
    \scr_ff_mux_state_427_13_g456/w_0 , \scr_ff_mux_state_427_13_g456/w_1 , 
    \scr_ff_mux_state_427_13_g456/w_2 , \scr_ff_mux_state_427_13_g456/w_3 , 
    \scr_ff_mux_state_427_13_g456/w_4 , \scr_ff_mux_state_427_13_g444/w_0 , 
    \scr_ff_mux_state_427_13_g444/w_1 , \scr_ff_mux_state_427_13_g444/w_2 , 
    \scr_ff_mux_state_427_13_g444/w_3 , \scr_ff_mux_state_427_13_g444/w_4 , 
    \scr_ff_mux_state_427_13_g428/w_0 , \scr_ff_mux_state_427_13_g428/w_1 , 
    \scr_ff_mux_state_427_13_g428/w_2 , \scr_ff_mux_state_427_13_g428/w_3 , 
    \scr_ff_mux_state_427_13_g428/w_4 , \scr_ff_mux_state_427_13_g416/w_0 , 
    \scr_ff_mux_state_427_13_g416/w_1 , \scr_ff_mux_state_427_13_g416/w_2 , 
    \scr_ff_mux_state_427_13_g416/w_3 , \scr_ff_mux_state_427_13_g416/w_4 , 
    \scr_ff_mux_state_427_13_g400/w_0 , \scr_ff_mux_state_427_13_g400/w_1 , 
    \scr_ff_mux_state_427_13_g400/w_2 , \scr_ff_mux_state_427_13_g400/w_3 , 
    \scr_ff_mux_state_427_13_g400/w_4 , \scr_ff_mux_state_427_13_g388/w_0 , 
    \scr_ff_mux_state_427_13_g388/w_1 , \scr_ff_mux_state_427_13_g388/w_2 , 
    \scr_ff_mux_state_427_13_g388/w_3 , \scr_ff_mux_state_427_13_g388/w_4 , 
    \scr_ff_mux_state_427_13_g372/w_0 , \scr_ff_mux_state_427_13_g372/w_1 , 
    \scr_ff_mux_state_427_13_g372/w_2 , \scr_ff_mux_state_427_13_g372/w_3 , 
    \scr_ff_mux_state_427_13_g372/w_4 , \scr_ff_mux_state_427_13_g360/w_0 , 
    \scr_ff_mux_state_427_13_g360/w_1 , \scr_ff_mux_state_427_13_g360/w_2 , 
    \scr_ff_mux_state_427_13_g360/w_3 , \scr_ff_mux_state_427_13_g360/w_4 , 
    n_1153, n_1152, n_1151, n_425, n_424, n_423, n_422, n_404, n_402, n_401, 
    n_398, n_397, n_395, n_394, n_392, n_391, n_389, n_388, n_386, n_385, 
    n_383, n_382, n_380, n_379, n_377, n_376, n_374, n_373, n_372, n_371, 
    n_370, n_369, n_368, n_367, n_366, n_364, n_361, n_360, n_359, n_357, 
    n_353, n_352, n_351, n_350, n_347, n_346, n_345, n_344, n_341, n_340, 
    n_339, n_338, n_337, n_335, n_334, n_333, n_332, n_331, n_330, n_328, 
    n_327, n_326, n_325, n_324, n_322, n_321, n_320, n_319, n_318, n_316, 
    n_315, n_314, n_313, n_312, n_311, n_309, n_308, n_307, n_306, n_305, 
    n_304, n_303, n_302, n_301, n_300, n_299, n_298, n_297, n_296, n_295, 
    n_294, n_293, n_292, n_291, n_290, n_289, n_288, n_287, n_286, n_285, 
    n_284, n_283, n_282, n_281, n_280, n_279, n_278, n_277, n_276, n_275, 
    n_274, n_273, n_272, n_271, n_270, n_269, n_268, n_267, n_112, n_107, 
    n_106, n_102, n_101, n_96, n_95, n_90, n_89, n_88, n_84, n_83, n_78, n_74, 
    n_73, n_72, a15, \a14[0] , \a13[0] , \a12[0] , \a11[0] , \a10[0] , \a9[0] , 
    \a8[0] , \a7[0] , \a6[0] , \a5[0] , \a4[0] , set, reset, clk, scr_run, 
    scr_init;
wire  \scr_ff_mux_state_427_13_g792/data3 , \scr_ff_mux_state_427_13_g792/data4 , 
    \scr_ff_mux_state_427_13_g780/data3 , \scr_ff_mux_state_427_13_g780/data4 , 
    \scr_ff_mux_state_427_13_g764/data3 , \scr_ff_mux_state_427_13_g764/data4 , 
    \scr_ff_mux_state_427_13_g752/data3 , \scr_ff_mux_state_427_13_g752/data4 , 
    \scr_ff_mux_state_427_13_g736/data3 , \scr_ff_mux_state_427_13_g736/data4 , 
    \scr_ff_mux_state_427_13_g724/data3 , \scr_ff_mux_state_427_13_g724/data4 , 
    \scr_ff_mux_state_427_13_g708/data3 , \scr_ff_mux_state_427_13_g708/data4 , 
    \scr_ff_mux_state_427_13_g696/data3 , \scr_ff_mux_state_427_13_g696/data4 , 
    \scr_ff_mux_state_427_13_g680/data3 , \scr_ff_mux_state_427_13_g680/data4 , 
    \scr_ff_mux_state_427_13_g668/data3 , \scr_ff_mux_state_427_13_g668/data4 , 
    \scr_ff_mux_state_427_13_g652/data3 , \scr_ff_mux_state_427_13_g652/data4 , 
    \scr_ff_mux_state_427_13_g640/data3 , \scr_ff_mux_state_427_13_g640/data4 , 
    \scr_ff_mux_state_427_13_g624/data3 , \scr_ff_mux_state_427_13_g624/data4 , 
    \scr_ff_mux_state_427_13_g612/data3 , \scr_ff_mux_state_427_13_g612/data4 , 
    \scr_ff_mux_state_427_13_g596/data3 , \scr_ff_mux_state_427_13_g596/data4 , 
    \scr_ff_mux_state_427_13_g584/data3 , \scr_ff_mux_state_427_13_g584/data4 , 
    \scr_ff_mux_state_427_13_g568/data3 , \scr_ff_mux_state_427_13_g568/data4 , 
    \scr_ff_mux_state_427_13_g556/data3 , \scr_ff_mux_state_427_13_g556/data4 , 
    \scr_ff_mux_state_427_13_g540/data3 , \scr_ff_mux_state_427_13_g540/data4 , 
    \scr_ff_mux_state_427_13_g528/data3 , \scr_ff_mux_state_427_13_g528/data4 , 
    \scr_ff_mux_state_427_13_g512/data3 , \scr_ff_mux_state_427_13_g512/data4 , 
    \scr_ff_mux_state_427_13_g500/data3 , \scr_ff_mux_state_427_13_g500/data4 , 
    \scr_ff_mux_state_427_13_g484/data3 , \scr_ff_mux_state_427_13_g484/data4 , 
    \scr_ff_mux_state_427_13_g472/data3 , \scr_ff_mux_state_427_13_g472/data4 , 
    \scr_ff_mux_state_427_13_g456/data3 , \scr_ff_mux_state_427_13_g456/data4 , 
    \scr_ff_mux_state_427_13_g444/data3 , \scr_ff_mux_state_427_13_g444/data4 , 
    \scr_ff_mux_state_427_13_g428/data3 , \scr_ff_mux_state_427_13_g428/data4 , 
    \scr_ff_mux_state_427_13_g416/data3 , \scr_ff_mux_state_427_13_g416/data4 , 
    \scr_ff_mux_state_427_13_g400/data3 , \scr_ff_mux_state_427_13_g400/data4 , 
    \scr_ff_mux_state_427_13_g388/data3 , \scr_ff_mux_state_427_13_g388/data4 , 
    \scr_ff_mux_state_427_13_g372/data3 , \scr_ff_mux_state_427_13_g372/data4 , 
    \scr_ff_mux_state_427_13_g360/data3 , \scr_ff_mux_state_427_13_g360/data4 ;
wire   [31:0] scr_out_p;
wire   [31:0] scr_in;
wire   [31:0] scr_out;
  assign \scr_ff_mux_state_427_13_g792/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g780/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g764/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g752/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g736/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g724/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g708/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g696/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g680/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g668/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g652/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g640/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g624/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g612/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g596/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g584/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g568/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g556/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g540/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g528/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g512/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g500/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g484/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g472/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g456/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g444/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g428/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g416/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g400/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g388/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g372/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g360/data4  = 1'b0;
  assign \scr_ff_mux_state_427_13_g792/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g780/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g764/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g752/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g736/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g724/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g708/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g696/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g680/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g668/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g652/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g640/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g624/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g612/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g596/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g584/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g568/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g556/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g540/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g528/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g512/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g500/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g484/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g472/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g456/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g444/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g428/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g416/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g400/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g388/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g372/data3  = 1'b1;
  assign \scr_ff_mux_state_427_13_g360/data3  = 1'b1;
  or \scr_ff_mux_state_427_13_g792/org (scr_out_p[27], 
    \scr_ff_mux_state_427_13_g792/w_0 , \scr_ff_mux_state_427_13_g792/w_1 , 
    \scr_ff_mux_state_427_13_g792/w_2 , \scr_ff_mux_state_427_13_g792/w_3 , 
    \scr_ff_mux_state_427_13_g792/w_4 );
  and \scr_ff_mux_state_427_13_g792/a_4 (\scr_ff_mux_state_427_13_g792/w_4 , set, 
    \scr_ff_mux_state_427_13_g792/data4 );
  and \scr_ff_mux_state_427_13_g792/a_3 (\scr_ff_mux_state_427_13_g792/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g792/data3 );
  and \scr_ff_mux_state_427_13_g792/a_2 (\scr_ff_mux_state_427_13_g792/w_2 , 
    n_424, scr_in[27]);
  and \scr_ff_mux_state_427_13_g792/a_1 (\scr_ff_mux_state_427_13_g792/w_1 , 
    n_423, n_285);
  and \scr_ff_mux_state_427_13_g792/a_0 (\scr_ff_mux_state_427_13_g792/w_0 , 
    n_422, scr_out[27]);
  or \scr_ff_mux_state_427_13_g780/org (scr_out_p[28], 
    \scr_ff_mux_state_427_13_g780/w_0 , \scr_ff_mux_state_427_13_g780/w_1 , 
    \scr_ff_mux_state_427_13_g780/w_2 , \scr_ff_mux_state_427_13_g780/w_3 , 
    \scr_ff_mux_state_427_13_g780/w_4 );
  and \scr_ff_mux_state_427_13_g780/a_4 (\scr_ff_mux_state_427_13_g780/w_4 , set, 
    \scr_ff_mux_state_427_13_g780/data4 );
  and \scr_ff_mux_state_427_13_g780/a_3 (\scr_ff_mux_state_427_13_g780/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g780/data3 );
  and \scr_ff_mux_state_427_13_g780/a_2 (\scr_ff_mux_state_427_13_g780/w_2 , 
    n_424, scr_in[28]);
  and \scr_ff_mux_state_427_13_g780/a_1 (\scr_ff_mux_state_427_13_g780/w_1 , 
    n_423, n_281);
  and \scr_ff_mux_state_427_13_g780/a_0 (\scr_ff_mux_state_427_13_g780/w_0 , 
    n_422, scr_out[28]);
  or \scr_ff_mux_state_427_13_g764/org (scr_out_p[29], 
    \scr_ff_mux_state_427_13_g764/w_0 , \scr_ff_mux_state_427_13_g764/w_1 , 
    \scr_ff_mux_state_427_13_g764/w_2 , \scr_ff_mux_state_427_13_g764/w_3 , 
    \scr_ff_mux_state_427_13_g764/w_4 );
  and \scr_ff_mux_state_427_13_g764/a_4 (\scr_ff_mux_state_427_13_g764/w_4 , set, 
    \scr_ff_mux_state_427_13_g764/data4 );
  and \scr_ff_mux_state_427_13_g764/a_3 (\scr_ff_mux_state_427_13_g764/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g764/data3 );
  and \scr_ff_mux_state_427_13_g764/a_2 (\scr_ff_mux_state_427_13_g764/w_2 , 
    n_424, scr_in[29]);
  and \scr_ff_mux_state_427_13_g764/a_1 (\scr_ff_mux_state_427_13_g764/w_1 , 
    n_423, n_277);
  and \scr_ff_mux_state_427_13_g764/a_0 (\scr_ff_mux_state_427_13_g764/w_0 , 
    n_422, scr_out[29]);
  or \scr_ff_mux_state_427_13_g752/org (scr_out_p[12], 
    \scr_ff_mux_state_427_13_g752/w_0 , \scr_ff_mux_state_427_13_g752/w_1 , 
    \scr_ff_mux_state_427_13_g752/w_2 , \scr_ff_mux_state_427_13_g752/w_3 , 
    \scr_ff_mux_state_427_13_g752/w_4 );
  and \scr_ff_mux_state_427_13_g752/a_4 (\scr_ff_mux_state_427_13_g752/w_4 , set, 
    \scr_ff_mux_state_427_13_g752/data4 );
  and \scr_ff_mux_state_427_13_g752/a_3 (\scr_ff_mux_state_427_13_g752/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g752/data3 );
  and \scr_ff_mux_state_427_13_g752/a_2 (\scr_ff_mux_state_427_13_g752/w_2 , 
    n_424, scr_in[12]);
  and \scr_ff_mux_state_427_13_g752/a_1 (\scr_ff_mux_state_427_13_g752/w_1 , 
    n_423, n_376);
  and \scr_ff_mux_state_427_13_g752/a_0 (\scr_ff_mux_state_427_13_g752/w_0 , 
    n_422, scr_out[12]);
  or \scr_ff_mux_state_427_13_g736/org (scr_out_p[30], 
    \scr_ff_mux_state_427_13_g736/w_0 , \scr_ff_mux_state_427_13_g736/w_1 , 
    \scr_ff_mux_state_427_13_g736/w_2 , \scr_ff_mux_state_427_13_g736/w_3 , 
    \scr_ff_mux_state_427_13_g736/w_4 );
  and \scr_ff_mux_state_427_13_g736/a_4 (\scr_ff_mux_state_427_13_g736/w_4 , set, 
    \scr_ff_mux_state_427_13_g736/data4 );
  and \scr_ff_mux_state_427_13_g736/a_3 (\scr_ff_mux_state_427_13_g736/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g736/data3 );
  and \scr_ff_mux_state_427_13_g736/a_2 (\scr_ff_mux_state_427_13_g736/w_2 , 
    n_424, scr_in[30]);
  and \scr_ff_mux_state_427_13_g736/a_1 (\scr_ff_mux_state_427_13_g736/w_1 , 
    n_423, n_273);
  and \scr_ff_mux_state_427_13_g736/a_0 (\scr_ff_mux_state_427_13_g736/w_0 , 
    n_422, scr_out[30]);
  or \scr_ff_mux_state_427_13_g724/org (scr_out_p[16], 
    \scr_ff_mux_state_427_13_g724/w_0 , \scr_ff_mux_state_427_13_g724/w_1 , 
    \scr_ff_mux_state_427_13_g724/w_2 , \scr_ff_mux_state_427_13_g724/w_3 , 
    \scr_ff_mux_state_427_13_g724/w_4 );
  and \scr_ff_mux_state_427_13_g724/a_4 (\scr_ff_mux_state_427_13_g724/w_4 , set, 
    \scr_ff_mux_state_427_13_g724/data4 );
  and \scr_ff_mux_state_427_13_g724/a_3 (\scr_ff_mux_state_427_13_g724/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g724/data3 );
  and \scr_ff_mux_state_427_13_g724/a_2 (\scr_ff_mux_state_427_13_g724/w_2 , 
    n_424, scr_in[16]);
  and \scr_ff_mux_state_427_13_g724/a_1 (\scr_ff_mux_state_427_13_g724/w_1 , 
    n_423, n_352);
  and \scr_ff_mux_state_427_13_g724/a_0 (\scr_ff_mux_state_427_13_g724/w_0 , 
    n_422, scr_out[16]);
  or \scr_ff_mux_state_427_13_g708/org (scr_out_p[31], 
    \scr_ff_mux_state_427_13_g708/w_0 , \scr_ff_mux_state_427_13_g708/w_1 , 
    \scr_ff_mux_state_427_13_g708/w_2 , \scr_ff_mux_state_427_13_g708/w_3 , 
    \scr_ff_mux_state_427_13_g708/w_4 );
  and \scr_ff_mux_state_427_13_g708/a_4 (\scr_ff_mux_state_427_13_g708/w_4 , set, 
    \scr_ff_mux_state_427_13_g708/data4 );
  and \scr_ff_mux_state_427_13_g708/a_3 (\scr_ff_mux_state_427_13_g708/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g708/data3 );
  and \scr_ff_mux_state_427_13_g708/a_2 (\scr_ff_mux_state_427_13_g708/w_2 , 
    n_424, scr_in[31]);
  and \scr_ff_mux_state_427_13_g708/a_1 (\scr_ff_mux_state_427_13_g708/w_1 , 
    n_423, n_269);
  and \scr_ff_mux_state_427_13_g708/a_0 (\scr_ff_mux_state_427_13_g708/w_0 , 
    n_422, scr_out[31]);
  or \scr_ff_mux_state_427_13_g696/org (scr_out_p[23], 
    \scr_ff_mux_state_427_13_g696/w_0 , \scr_ff_mux_state_427_13_g696/w_1 , 
    \scr_ff_mux_state_427_13_g696/w_2 , \scr_ff_mux_state_427_13_g696/w_3 , 
    \scr_ff_mux_state_427_13_g696/w_4 );
  and \scr_ff_mux_state_427_13_g696/a_4 (\scr_ff_mux_state_427_13_g696/w_4 , set, 
    \scr_ff_mux_state_427_13_g696/data4 );
  and \scr_ff_mux_state_427_13_g696/a_3 (\scr_ff_mux_state_427_13_g696/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g696/data3 );
  and \scr_ff_mux_state_427_13_g696/a_2 (\scr_ff_mux_state_427_13_g696/w_2 , 
    n_424, scr_in[23]);
  and \scr_ff_mux_state_427_13_g696/a_1 (\scr_ff_mux_state_427_13_g696/w_1 , 
    n_423, n_306);
  and \scr_ff_mux_state_427_13_g696/a_0 (\scr_ff_mux_state_427_13_g696/w_0 , 
    n_422, scr_out[23]);
  or \scr_ff_mux_state_427_13_g680/org (scr_out_p[24], 
    \scr_ff_mux_state_427_13_g680/w_0 , \scr_ff_mux_state_427_13_g680/w_1 , 
    \scr_ff_mux_state_427_13_g680/w_2 , \scr_ff_mux_state_427_13_g680/w_3 , 
    \scr_ff_mux_state_427_13_g680/w_4 );
  and \scr_ff_mux_state_427_13_g680/a_4 (\scr_ff_mux_state_427_13_g680/w_4 , set, 
    \scr_ff_mux_state_427_13_g680/data4 );
  and \scr_ff_mux_state_427_13_g680/a_3 (\scr_ff_mux_state_427_13_g680/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g680/data3 );
  and \scr_ff_mux_state_427_13_g680/a_2 (\scr_ff_mux_state_427_13_g680/w_2 , 
    n_424, scr_in[24]);
  and \scr_ff_mux_state_427_13_g680/a_1 (\scr_ff_mux_state_427_13_g680/w_1 , 
    n_423, n_300);
  and \scr_ff_mux_state_427_13_g680/a_0 (\scr_ff_mux_state_427_13_g680/w_0 , 
    n_422, scr_out[24]);
  or \scr_ff_mux_state_427_13_g668/org (scr_out_p[26], 
    \scr_ff_mux_state_427_13_g668/w_0 , \scr_ff_mux_state_427_13_g668/w_1 , 
    \scr_ff_mux_state_427_13_g668/w_2 , \scr_ff_mux_state_427_13_g668/w_3 , 
    \scr_ff_mux_state_427_13_g668/w_4 );
  and \scr_ff_mux_state_427_13_g668/a_4 (\scr_ff_mux_state_427_13_g668/w_4 , set, 
    \scr_ff_mux_state_427_13_g668/data4 );
  and \scr_ff_mux_state_427_13_g668/a_3 (\scr_ff_mux_state_427_13_g668/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g668/data3 );
  and \scr_ff_mux_state_427_13_g668/a_2 (\scr_ff_mux_state_427_13_g668/w_2 , 
    n_424, scr_in[26]);
  and \scr_ff_mux_state_427_13_g668/a_1 (\scr_ff_mux_state_427_13_g668/w_1 , 
    n_423, n_290);
  and \scr_ff_mux_state_427_13_g668/a_0 (\scr_ff_mux_state_427_13_g668/w_0 , 
    n_422, scr_out[26]);
  or \scr_ff_mux_state_427_13_g652/org (scr_out_p[9], 
    \scr_ff_mux_state_427_13_g652/w_0 , \scr_ff_mux_state_427_13_g652/w_1 , 
    \scr_ff_mux_state_427_13_g652/w_2 , \scr_ff_mux_state_427_13_g652/w_3 , 
    \scr_ff_mux_state_427_13_g652/w_4 );
  and \scr_ff_mux_state_427_13_g652/a_4 (\scr_ff_mux_state_427_13_g652/w_4 , set, 
    \scr_ff_mux_state_427_13_g652/data4 );
  and \scr_ff_mux_state_427_13_g652/a_3 (\scr_ff_mux_state_427_13_g652/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g652/data3 );
  and \scr_ff_mux_state_427_13_g652/a_2 (\scr_ff_mux_state_427_13_g652/w_2 , 
    n_424, scr_in[9]);
  and \scr_ff_mux_state_427_13_g652/a_1 (\scr_ff_mux_state_427_13_g652/w_1 , 
    n_423, n_385);
  and \scr_ff_mux_state_427_13_g652/a_0 (\scr_ff_mux_state_427_13_g652/w_0 , 
    n_422, scr_out[9]);
  or \scr_ff_mux_state_427_13_g640/org (scr_out_p[10], 
    \scr_ff_mux_state_427_13_g640/w_0 , \scr_ff_mux_state_427_13_g640/w_1 , 
    \scr_ff_mux_state_427_13_g640/w_2 , \scr_ff_mux_state_427_13_g640/w_3 , 
    \scr_ff_mux_state_427_13_g640/w_4 );
  and \scr_ff_mux_state_427_13_g640/a_4 (\scr_ff_mux_state_427_13_g640/w_4 , set, 
    \scr_ff_mux_state_427_13_g640/data4 );
  and \scr_ff_mux_state_427_13_g640/a_3 (\scr_ff_mux_state_427_13_g640/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g640/data3 );
  and \scr_ff_mux_state_427_13_g640/a_2 (\scr_ff_mux_state_427_13_g640/w_2 , 
    n_424, scr_in[10]);
  and \scr_ff_mux_state_427_13_g640/a_1 (\scr_ff_mux_state_427_13_g640/w_1 , 
    n_423, n_382);
  and \scr_ff_mux_state_427_13_g640/a_0 (\scr_ff_mux_state_427_13_g640/w_0 , 
    n_422, scr_out[10]);
  or \scr_ff_mux_state_427_13_g624/org (scr_out_p[11], 
    \scr_ff_mux_state_427_13_g624/w_0 , \scr_ff_mux_state_427_13_g624/w_1 , 
    \scr_ff_mux_state_427_13_g624/w_2 , \scr_ff_mux_state_427_13_g624/w_3 , 
    \scr_ff_mux_state_427_13_g624/w_4 );
  and \scr_ff_mux_state_427_13_g624/a_4 (\scr_ff_mux_state_427_13_g624/w_4 , set, 
    \scr_ff_mux_state_427_13_g624/data4 );
  and \scr_ff_mux_state_427_13_g624/a_3 (\scr_ff_mux_state_427_13_g624/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g624/data3 );
  and \scr_ff_mux_state_427_13_g624/a_2 (\scr_ff_mux_state_427_13_g624/w_2 , 
    n_424, scr_in[11]);
  and \scr_ff_mux_state_427_13_g624/a_1 (\scr_ff_mux_state_427_13_g624/w_1 , 
    n_423, n_379);
  and \scr_ff_mux_state_427_13_g624/a_0 (\scr_ff_mux_state_427_13_g624/w_0 , 
    n_422, scr_out[11]);
  or \scr_ff_mux_state_427_13_g612/org (scr_out_p[15], 
    \scr_ff_mux_state_427_13_g612/w_0 , \scr_ff_mux_state_427_13_g612/w_1 , 
    \scr_ff_mux_state_427_13_g612/w_2 , \scr_ff_mux_state_427_13_g612/w_3 , 
    \scr_ff_mux_state_427_13_g612/w_4 );
  and \scr_ff_mux_state_427_13_g612/a_4 (\scr_ff_mux_state_427_13_g612/w_4 , set, 
    \scr_ff_mux_state_427_13_g612/data4 );
  and \scr_ff_mux_state_427_13_g612/a_3 (\scr_ff_mux_state_427_13_g612/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g612/data3 );
  and \scr_ff_mux_state_427_13_g612/a_2 (\scr_ff_mux_state_427_13_g612/w_2 , 
    n_424, scr_in[15]);
  and \scr_ff_mux_state_427_13_g612/a_1 (\scr_ff_mux_state_427_13_g612/w_1 , 
    n_423, n_359);
  and \scr_ff_mux_state_427_13_g612/a_0 (\scr_ff_mux_state_427_13_g612/w_0 , 
    n_422, scr_out[15]);
  or \scr_ff_mux_state_427_13_g596/org (scr_out_p[25], 
    \scr_ff_mux_state_427_13_g596/w_0 , \scr_ff_mux_state_427_13_g596/w_1 , 
    \scr_ff_mux_state_427_13_g596/w_2 , \scr_ff_mux_state_427_13_g596/w_3 , 
    \scr_ff_mux_state_427_13_g596/w_4 );
  and \scr_ff_mux_state_427_13_g596/a_4 (\scr_ff_mux_state_427_13_g596/w_4 , set, 
    \scr_ff_mux_state_427_13_g596/data4 );
  and \scr_ff_mux_state_427_13_g596/a_3 (\scr_ff_mux_state_427_13_g596/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g596/data3 );
  and \scr_ff_mux_state_427_13_g596/a_2 (\scr_ff_mux_state_427_13_g596/w_2 , 
    n_424, scr_in[25]);
  and \scr_ff_mux_state_427_13_g596/a_1 (\scr_ff_mux_state_427_13_g596/w_1 , 
    n_423, n_295);
  and \scr_ff_mux_state_427_13_g596/a_0 (\scr_ff_mux_state_427_13_g596/w_0 , 
    n_422, scr_out[25]);
  or \scr_ff_mux_state_427_13_g584/org (scr_out_p[8], 
    \scr_ff_mux_state_427_13_g584/w_0 , \scr_ff_mux_state_427_13_g584/w_1 , 
    \scr_ff_mux_state_427_13_g584/w_2 , \scr_ff_mux_state_427_13_g584/w_3 , 
    \scr_ff_mux_state_427_13_g584/w_4 );
  and \scr_ff_mux_state_427_13_g584/a_4 (\scr_ff_mux_state_427_13_g584/w_4 , set, 
    \scr_ff_mux_state_427_13_g584/data4 );
  and \scr_ff_mux_state_427_13_g584/a_3 (\scr_ff_mux_state_427_13_g584/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g584/data3 );
  and \scr_ff_mux_state_427_13_g584/a_2 (\scr_ff_mux_state_427_13_g584/w_2 , 
    n_424, scr_in[8]);
  and \scr_ff_mux_state_427_13_g584/a_1 (\scr_ff_mux_state_427_13_g584/w_1 , 
    n_423, n_388);
  and \scr_ff_mux_state_427_13_g584/a_0 (\scr_ff_mux_state_427_13_g584/w_0 , 
    n_422, scr_out[8]);
  or \scr_ff_mux_state_427_13_g568/org (scr_out_p[13], 
    \scr_ff_mux_state_427_13_g568/w_0 , \scr_ff_mux_state_427_13_g568/w_1 , 
    \scr_ff_mux_state_427_13_g568/w_2 , \scr_ff_mux_state_427_13_g568/w_3 , 
    \scr_ff_mux_state_427_13_g568/w_4 );
  and \scr_ff_mux_state_427_13_g568/a_4 (\scr_ff_mux_state_427_13_g568/w_4 , set, 
    \scr_ff_mux_state_427_13_g568/data4 );
  and \scr_ff_mux_state_427_13_g568/a_3 (\scr_ff_mux_state_427_13_g568/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g568/data3 );
  and \scr_ff_mux_state_427_13_g568/a_2 (\scr_ff_mux_state_427_13_g568/w_2 , 
    n_424, scr_in[13]);
  and \scr_ff_mux_state_427_13_g568/a_1 (\scr_ff_mux_state_427_13_g568/w_1 , 
    n_423, n_373);
  and \scr_ff_mux_state_427_13_g568/a_0 (\scr_ff_mux_state_427_13_g568/w_0 , 
    n_422, scr_out[13]);
  or \scr_ff_mux_state_427_13_g556/org (scr_out_p[14], 
    \scr_ff_mux_state_427_13_g556/w_0 , \scr_ff_mux_state_427_13_g556/w_1 , 
    \scr_ff_mux_state_427_13_g556/w_2 , \scr_ff_mux_state_427_13_g556/w_3 , 
    \scr_ff_mux_state_427_13_g556/w_4 );
  and \scr_ff_mux_state_427_13_g556/a_4 (\scr_ff_mux_state_427_13_g556/w_4 , set, 
    \scr_ff_mux_state_427_13_g556/data4 );
  and \scr_ff_mux_state_427_13_g556/a_3 (\scr_ff_mux_state_427_13_g556/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g556/data3 );
  and \scr_ff_mux_state_427_13_g556/a_2 (\scr_ff_mux_state_427_13_g556/w_2 , 
    n_424, scr_in[14]);
  and \scr_ff_mux_state_427_13_g556/a_1 (\scr_ff_mux_state_427_13_g556/w_1 , 
    n_423, n_366);
  and \scr_ff_mux_state_427_13_g556/a_0 (\scr_ff_mux_state_427_13_g556/w_0 , 
    n_422, scr_out[14]);
  or \scr_ff_mux_state_427_13_g540/org (scr_out_p[17], 
    \scr_ff_mux_state_427_13_g540/w_0 , \scr_ff_mux_state_427_13_g540/w_1 , 
    \scr_ff_mux_state_427_13_g540/w_2 , \scr_ff_mux_state_427_13_g540/w_3 , 
    \scr_ff_mux_state_427_13_g540/w_4 );
  and \scr_ff_mux_state_427_13_g540/a_4 (\scr_ff_mux_state_427_13_g540/w_4 , set, 
    \scr_ff_mux_state_427_13_g540/data4 );
  and \scr_ff_mux_state_427_13_g540/a_3 (\scr_ff_mux_state_427_13_g540/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g540/data3 );
  and \scr_ff_mux_state_427_13_g540/a_2 (\scr_ff_mux_state_427_13_g540/w_2 , 
    n_424, scr_in[17]);
  and \scr_ff_mux_state_427_13_g540/a_1 (\scr_ff_mux_state_427_13_g540/w_1 , 
    n_423, n_346);
  and \scr_ff_mux_state_427_13_g540/a_0 (\scr_ff_mux_state_427_13_g540/w_0 , 
    n_422, scr_out[17]);
  or \scr_ff_mux_state_427_13_g528/org (scr_out_p[18], 
    \scr_ff_mux_state_427_13_g528/w_0 , \scr_ff_mux_state_427_13_g528/w_1 , 
    \scr_ff_mux_state_427_13_g528/w_2 , \scr_ff_mux_state_427_13_g528/w_3 , 
    \scr_ff_mux_state_427_13_g528/w_4 );
  and \scr_ff_mux_state_427_13_g528/a_4 (\scr_ff_mux_state_427_13_g528/w_4 , set, 
    \scr_ff_mux_state_427_13_g528/data4 );
  and \scr_ff_mux_state_427_13_g528/a_3 (\scr_ff_mux_state_427_13_g528/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g528/data3 );
  and \scr_ff_mux_state_427_13_g528/a_2 (\scr_ff_mux_state_427_13_g528/w_2 , 
    n_424, scr_in[18]);
  and \scr_ff_mux_state_427_13_g528/a_1 (\scr_ff_mux_state_427_13_g528/w_1 , 
    n_423, n_339);
  and \scr_ff_mux_state_427_13_g528/a_0 (\scr_ff_mux_state_427_13_g528/w_0 , 
    n_422, scr_out[18]);
  or \scr_ff_mux_state_427_13_g512/org (scr_out_p[22], 
    \scr_ff_mux_state_427_13_g512/w_0 , \scr_ff_mux_state_427_13_g512/w_1 , 
    \scr_ff_mux_state_427_13_g512/w_2 , \scr_ff_mux_state_427_13_g512/w_3 , 
    \scr_ff_mux_state_427_13_g512/w_4 );
  and \scr_ff_mux_state_427_13_g512/a_4 (\scr_ff_mux_state_427_13_g512/w_4 , set, 
    \scr_ff_mux_state_427_13_g512/data4 );
  and \scr_ff_mux_state_427_13_g512/a_3 (\scr_ff_mux_state_427_13_g512/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g512/data3 );
  and \scr_ff_mux_state_427_13_g512/a_2 (\scr_ff_mux_state_427_13_g512/w_2 , 
    n_424, scr_in[22]);
  and \scr_ff_mux_state_427_13_g512/a_1 (\scr_ff_mux_state_427_13_g512/w_1 , 
    n_423, n_313);
  and \scr_ff_mux_state_427_13_g512/a_0 (\scr_ff_mux_state_427_13_g512/w_0 , 
    n_422, scr_out[22]);
  or \scr_ff_mux_state_427_13_g500/org (scr_out_p[7], 
    \scr_ff_mux_state_427_13_g500/w_0 , \scr_ff_mux_state_427_13_g500/w_1 , 
    \scr_ff_mux_state_427_13_g500/w_2 , \scr_ff_mux_state_427_13_g500/w_3 , 
    \scr_ff_mux_state_427_13_g500/w_4 );
  and \scr_ff_mux_state_427_13_g500/a_4 (\scr_ff_mux_state_427_13_g500/w_4 , set, 
    \scr_ff_mux_state_427_13_g500/data4 );
  and \scr_ff_mux_state_427_13_g500/a_3 (\scr_ff_mux_state_427_13_g500/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g500/data3 );
  and \scr_ff_mux_state_427_13_g500/a_2 (\scr_ff_mux_state_427_13_g500/w_2 , 
    n_424, scr_in[7]);
  and \scr_ff_mux_state_427_13_g500/a_1 (\scr_ff_mux_state_427_13_g500/w_1 , 
    n_423, n_391);
  and \scr_ff_mux_state_427_13_g500/a_0 (\scr_ff_mux_state_427_13_g500/w_0 , 
    n_422, scr_out[7]);
  or \scr_ff_mux_state_427_13_g484/org (scr_out_p[21], 
    \scr_ff_mux_state_427_13_g484/w_0 , \scr_ff_mux_state_427_13_g484/w_1 , 
    \scr_ff_mux_state_427_13_g484/w_2 , \scr_ff_mux_state_427_13_g484/w_3 , 
    \scr_ff_mux_state_427_13_g484/w_4 );
  and \scr_ff_mux_state_427_13_g484/a_4 (\scr_ff_mux_state_427_13_g484/w_4 , set, 
    \scr_ff_mux_state_427_13_g484/data4 );
  and \scr_ff_mux_state_427_13_g484/a_3 (\scr_ff_mux_state_427_13_g484/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g484/data3 );
  and \scr_ff_mux_state_427_13_g484/a_2 (\scr_ff_mux_state_427_13_g484/w_2 , 
    n_424, scr_in[21]);
  and \scr_ff_mux_state_427_13_g484/a_1 (\scr_ff_mux_state_427_13_g484/w_1 , 
    n_423, n_320);
  and \scr_ff_mux_state_427_13_g484/a_0 (\scr_ff_mux_state_427_13_g484/w_0 , 
    n_422, scr_out[21]);
  or \scr_ff_mux_state_427_13_g472/org (scr_out_p[2], 
    \scr_ff_mux_state_427_13_g472/w_0 , \scr_ff_mux_state_427_13_g472/w_1 , 
    \scr_ff_mux_state_427_13_g472/w_2 , \scr_ff_mux_state_427_13_g472/w_3 , 
    \scr_ff_mux_state_427_13_g472/w_4 );
  and \scr_ff_mux_state_427_13_g472/a_4 (\scr_ff_mux_state_427_13_g472/w_4 , set, 
    \scr_ff_mux_state_427_13_g472/data4 );
  and \scr_ff_mux_state_427_13_g472/a_3 (\scr_ff_mux_state_427_13_g472/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g472/data3 );
  and \scr_ff_mux_state_427_13_g472/a_2 (\scr_ff_mux_state_427_13_g472/w_2 , 
    n_424, scr_in[2]);
  and \scr_ff_mux_state_427_13_g472/a_1 (\scr_ff_mux_state_427_13_g472/w_1 , 
    n_423, n_95);
  and \scr_ff_mux_state_427_13_g472/a_0 (\scr_ff_mux_state_427_13_g472/w_0 , 
    n_422, scr_out[2]);
  or \scr_ff_mux_state_427_13_g456/org (scr_out_p[3], 
    \scr_ff_mux_state_427_13_g456/w_0 , \scr_ff_mux_state_427_13_g456/w_1 , 
    \scr_ff_mux_state_427_13_g456/w_2 , \scr_ff_mux_state_427_13_g456/w_3 , 
    \scr_ff_mux_state_427_13_g456/w_4 );
  and \scr_ff_mux_state_427_13_g456/a_4 (\scr_ff_mux_state_427_13_g456/w_4 , set, 
    \scr_ff_mux_state_427_13_g456/data4 );
  and \scr_ff_mux_state_427_13_g456/a_3 (\scr_ff_mux_state_427_13_g456/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g456/data3 );
  and \scr_ff_mux_state_427_13_g456/a_2 (\scr_ff_mux_state_427_13_g456/w_2 , 
    n_424, scr_in[3]);
  and \scr_ff_mux_state_427_13_g456/a_1 (\scr_ff_mux_state_427_13_g456/w_1 , 
    n_423, n_89);
  and \scr_ff_mux_state_427_13_g456/a_0 (\scr_ff_mux_state_427_13_g456/w_0 , 
    n_422, scr_out[3]);
  or \scr_ff_mux_state_427_13_g444/org (scr_out_p[4], 
    \scr_ff_mux_state_427_13_g444/w_0 , \scr_ff_mux_state_427_13_g444/w_1 , 
    \scr_ff_mux_state_427_13_g444/w_2 , \scr_ff_mux_state_427_13_g444/w_3 , 
    \scr_ff_mux_state_427_13_g444/w_4 );
  and \scr_ff_mux_state_427_13_g444/a_4 (\scr_ff_mux_state_427_13_g444/w_4 , set, 
    \scr_ff_mux_state_427_13_g444/data4 );
  and \scr_ff_mux_state_427_13_g444/a_3 (\scr_ff_mux_state_427_13_g444/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g444/data3 );
  and \scr_ff_mux_state_427_13_g444/a_2 (\scr_ff_mux_state_427_13_g444/w_2 , 
    n_424, scr_in[4]);
  and \scr_ff_mux_state_427_13_g444/a_1 (\scr_ff_mux_state_427_13_g444/w_1 , 
    n_423, n_83);
  and \scr_ff_mux_state_427_13_g444/a_0 (\scr_ff_mux_state_427_13_g444/w_0 , 
    n_422, scr_out[4]);
  or \scr_ff_mux_state_427_13_g428/org (scr_out_p[5], 
    \scr_ff_mux_state_427_13_g428/w_0 , \scr_ff_mux_state_427_13_g428/w_1 , 
    \scr_ff_mux_state_427_13_g428/w_2 , \scr_ff_mux_state_427_13_g428/w_3 , 
    \scr_ff_mux_state_427_13_g428/w_4 );
  and \scr_ff_mux_state_427_13_g428/a_4 (\scr_ff_mux_state_427_13_g428/w_4 , set, 
    \scr_ff_mux_state_427_13_g428/data4 );
  and \scr_ff_mux_state_427_13_g428/a_3 (\scr_ff_mux_state_427_13_g428/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g428/data3 );
  and \scr_ff_mux_state_427_13_g428/a_2 (\scr_ff_mux_state_427_13_g428/w_2 , 
    n_424, scr_in[5]);
  and \scr_ff_mux_state_427_13_g428/a_1 (\scr_ff_mux_state_427_13_g428/w_1 , 
    n_423, n_397);
  and \scr_ff_mux_state_427_13_g428/a_0 (\scr_ff_mux_state_427_13_g428/w_0 , 
    n_422, scr_out[5]);
  or \scr_ff_mux_state_427_13_g416/org (scr_out_p[6], 
    \scr_ff_mux_state_427_13_g416/w_0 , \scr_ff_mux_state_427_13_g416/w_1 , 
    \scr_ff_mux_state_427_13_g416/w_2 , \scr_ff_mux_state_427_13_g416/w_3 , 
    \scr_ff_mux_state_427_13_g416/w_4 );
  and \scr_ff_mux_state_427_13_g416/a_4 (\scr_ff_mux_state_427_13_g416/w_4 , set, 
    \scr_ff_mux_state_427_13_g416/data4 );
  and \scr_ff_mux_state_427_13_g416/a_3 (\scr_ff_mux_state_427_13_g416/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g416/data3 );
  and \scr_ff_mux_state_427_13_g416/a_2 (\scr_ff_mux_state_427_13_g416/w_2 , 
    n_424, scr_in[6]);
  and \scr_ff_mux_state_427_13_g416/a_1 (\scr_ff_mux_state_427_13_g416/w_1 , 
    n_423, n_394);
  and \scr_ff_mux_state_427_13_g416/a_0 (\scr_ff_mux_state_427_13_g416/w_0 , 
    n_422, scr_out[6]);
  or \scr_ff_mux_state_427_13_g400/org (scr_out_p[19], 
    \scr_ff_mux_state_427_13_g400/w_0 , \scr_ff_mux_state_427_13_g400/w_1 , 
    \scr_ff_mux_state_427_13_g400/w_2 , \scr_ff_mux_state_427_13_g400/w_3 , 
    \scr_ff_mux_state_427_13_g400/w_4 );
  and \scr_ff_mux_state_427_13_g400/a_4 (\scr_ff_mux_state_427_13_g400/w_4 , set, 
    \scr_ff_mux_state_427_13_g400/data4 );
  and \scr_ff_mux_state_427_13_g400/a_3 (\scr_ff_mux_state_427_13_g400/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g400/data3 );
  and \scr_ff_mux_state_427_13_g400/a_2 (\scr_ff_mux_state_427_13_g400/w_2 , 
    n_424, scr_in[19]);
  and \scr_ff_mux_state_427_13_g400/a_1 (\scr_ff_mux_state_427_13_g400/w_1 , 
    n_423, n_333);
  and \scr_ff_mux_state_427_13_g400/a_0 (\scr_ff_mux_state_427_13_g400/w_0 , 
    n_422, scr_out[19]);
  or \scr_ff_mux_state_427_13_g388/org (scr_out_p[20], 
    \scr_ff_mux_state_427_13_g388/w_0 , \scr_ff_mux_state_427_13_g388/w_1 , 
    \scr_ff_mux_state_427_13_g388/w_2 , \scr_ff_mux_state_427_13_g388/w_3 , 
    \scr_ff_mux_state_427_13_g388/w_4 );
  and \scr_ff_mux_state_427_13_g388/a_4 (\scr_ff_mux_state_427_13_g388/w_4 , set, 
    \scr_ff_mux_state_427_13_g388/data4 );
  and \scr_ff_mux_state_427_13_g388/a_3 (\scr_ff_mux_state_427_13_g388/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g388/data3 );
  and \scr_ff_mux_state_427_13_g388/a_2 (\scr_ff_mux_state_427_13_g388/w_2 , 
    n_424, scr_in[20]);
  and \scr_ff_mux_state_427_13_g388/a_1 (\scr_ff_mux_state_427_13_g388/w_1 , 
    n_423, n_326);
  and \scr_ff_mux_state_427_13_g388/a_0 (\scr_ff_mux_state_427_13_g388/w_0 , 
    n_422, scr_out[20]);
  or \scr_ff_mux_state_427_13_g372/org (scr_out_p[1], 
    \scr_ff_mux_state_427_13_g372/w_0 , \scr_ff_mux_state_427_13_g372/w_1 , 
    \scr_ff_mux_state_427_13_g372/w_2 , \scr_ff_mux_state_427_13_g372/w_3 , 
    \scr_ff_mux_state_427_13_g372/w_4 );
  and \scr_ff_mux_state_427_13_g372/a_4 (\scr_ff_mux_state_427_13_g372/w_4 , set, 
    \scr_ff_mux_state_427_13_g372/data4 );
  and \scr_ff_mux_state_427_13_g372/a_3 (\scr_ff_mux_state_427_13_g372/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g372/data3 );
  and \scr_ff_mux_state_427_13_g372/a_2 (\scr_ff_mux_state_427_13_g372/w_2 , 
    n_424, scr_in[1]);
  and \scr_ff_mux_state_427_13_g372/a_1 (\scr_ff_mux_state_427_13_g372/w_1 , 
    n_423, n_74);
  and \scr_ff_mux_state_427_13_g372/a_0 (\scr_ff_mux_state_427_13_g372/w_0 , 
    n_422, scr_out[1]);
  or \scr_ff_mux_state_427_13_g360/org (scr_out_p[0], 
    \scr_ff_mux_state_427_13_g360/w_0 , \scr_ff_mux_state_427_13_g360/w_1 , 
    \scr_ff_mux_state_427_13_g360/w_2 , \scr_ff_mux_state_427_13_g360/w_3 , 
    \scr_ff_mux_state_427_13_g360/w_4 );
  and \scr_ff_mux_state_427_13_g360/a_4 (\scr_ff_mux_state_427_13_g360/w_4 , set, 
    \scr_ff_mux_state_427_13_g360/data4 );
  and \scr_ff_mux_state_427_13_g360/a_3 (\scr_ff_mux_state_427_13_g360/w_3 , 
    n_425, \scr_ff_mux_state_427_13_g360/data3 );
  and \scr_ff_mux_state_427_13_g360/a_2 (\scr_ff_mux_state_427_13_g360/w_2 , 
    n_424, scr_in[0]);
  and \scr_ff_mux_state_427_13_g360/a_1 (\scr_ff_mux_state_427_13_g360/w_1 , 
    n_423, a15);
  and \scr_ff_mux_state_427_13_g360/a_0 (\scr_ff_mux_state_427_13_g360/w_0 , 
    n_422, scr_out[0]);
  xor g10(\a10[0] , scr_out[25], scr_out[21]);
  xor g11(\a9[0] , scr_out[26], scr_out[22]);
  xor g12(\a8[0] , scr_out[27], scr_out[23]);
  xor g13(\a7[0] , scr_out[28], scr_out[24]);
  xor g14(\a6[0] , scr_out[29], scr_out[25]);
  xor g15(\a5[0] , scr_out[30], scr_out[26]);
  xor g16(\a4[0] , scr_out[31], scr_out[27]);
  xor g17(n_74, a15, \a14[0] );
  xor g209(n_267, n_78, \a6[0] );
  xor g210(n_268, \a5[0] , scr_out[31]);
  xor g211(n_269, n_267, n_268);
  xor g212(n_270, n_84, \a7[0] );
  xor g213(n_271, \a6[0] , scr_out[30]);
  xor g214(n_272, scr_out[31], n_270);
  xor g215(n_273, n_271, n_272);
  xor g216(n_274, n_90, \a8[0] );
  xor g217(n_275, \a7[0] , scr_out[29]);
  xor g218(n_276, scr_out[30], n_274);
  xor g219(n_277, n_275, n_276);
  xor g220(n_278, n_96, \a9[0] );
  xor g221(n_279, \a8[0] , scr_out[28]);
  xor g222(n_280, scr_out[29], n_278);
  xor g223(n_281, n_279, n_280);
  xor g224(n_282, n_102, \a9[0] );
  xor g225(n_283, \a4[0] , scr_out[28]);
  xor g226(n_284, scr_out[31], n_282);
  xor g227(n_285, n_283, n_284);
  xor g228(n_286, n_107, \a10[0] );
  xor g229(n_287, \a5[0] , \a4[0] );
  xor g230(n_288, scr_out[30], scr_out[31]);
  xor g231(n_289, n_286, n_287);
  xor g232(n_290, n_288, n_289);
  xor g233(n_291, n_112, \a11[0] );
  xor g234(n_292, \a6[0] , \a5[0] );
  xor g235(n_293, scr_out[29], scr_out[30]);
  xor g236(n_294, n_291, n_292);
  xor g237(n_295, n_293, n_294);
  xor g238(n_296, n_89, \a7[0] );
  xor g239(n_297, \a6[0] , scr_out[28]);
  xor g240(n_298, scr_out[29], scr_out[31]);
  xor g241(n_299, n_296, n_297);
  xor g242(n_300, n_298, n_299);
  xor g243(n_301, n_95, \a8[0] );
  xor g244(n_302, \a7[0] , \a4[0] );
  xor g245(n_303, scr_out[28], scr_out[30]);
  xor g246(n_304, scr_out[31], n_301);
  xor g247(n_305, n_302, n_303);
  xor g248(n_306, n_304, n_305);
  xor g249(n_307, n_74, \a9[0] );
  xor g250(n_308, \a8[0] , \a5[0] );
  xor g251(n_309, \a4[0] , scr_out[29]);
  xor g253(n_311, n_307, n_308);
  xor g254(n_312, n_309, n_288);
  xor g255(n_313, n_311, n_312);
  xor g256(n_314, a15, \a10[0] );
  xor g257(n_315, \a9[0] , \a6[0] );
  xor g258(n_316, \a5[0] , scr_out[28]);
  xor g260(n_318, n_314, n_315);
  xor g261(n_319, n_316, n_293);
  xor g262(n_320, n_318, n_319);
  xor g263(n_321, \a11[0] , \a10[0] );
  xor g264(n_322, \a7[0] , \a6[0] );
  xor g266(n_324, scr_out[29], n_321);
  xor g267(n_325, n_322, n_283);
  xor g268(n_326, n_324, n_325);
  xor g269(n_327, \a12[0] , \a11[0] );
  xor g270(n_328, \a8[0] , \a7[0] );
  xor g272(n_330, scr_out[28], scr_out[31]);
  xor g273(n_331, n_327, n_328);
  xor g274(n_332, n_287, n_330);
  xor g275(n_333, n_331, n_332);
  xor g276(n_334, n_112, \a9[0] );
  xor g277(n_335, \a8[0] , \a6[0] );
  xor g279(n_337, scr_out[30], n_334);
  xor g28(n_84, n_83, \a8[0] );
  xor g280(n_338, n_335, n_287);
  xor g281(n_339, n_337, n_338);
  xor g282(n_340, n_88, \a10[0] );
  xor g283(n_341, \a9[0] , \a7[0] );
  xor g286(n_344, n_340, n_341);
  xor g287(n_345, n_292, n_298);
  xor g288(n_346, n_344, n_345);
  xor g289(n_347, n_102, \a8[0] );
  xor g292(n_350, scr_out[31], n_347);
  xor g293(n_351, n_322, n_303);
  xor g294(n_352, n_350, n_351);
  xor g295(n_353, n_107, \a9[0] );
  xor g299(n_357, n_353, n_328);
  xor g301(n_359, n_357, n_312);
  xor g302(n_360, n_112, \a10[0] );
  xor g303(n_361, \a9[0] , \a8[0] );
  xor g306(n_364, n_360, n_361);
  xor g308(n_366, n_364, n_319);
  xor g309(n_367, n_88, \a11[0] );
  xor g310(n_368, \a10[0] , \a9[0] );
  xor g311(n_369, \a6[0] , \a4[0] );
  xor g312(n_370, scr_out[28], scr_out[29]);
  xor g313(n_371, n_367, n_368);
  xor g314(n_372, n_369, n_370);
  xor g315(n_373, n_371, n_372);
  xor g316(n_374, n_78, \a5[0] );
  xor g318(n_376, n_374, n_283);
  xor g319(n_377, n_84, \a6[0] );
  xor g321(n_379, n_377, n_287);
  xor g322(n_380, n_90, \a7[0] );
  xor g324(n_382, n_380, n_292);
  xor g325(n_383, n_96, \a8[0] );
  xor g327(n_385, n_383, n_322);
  xor g328(n_386, n_101, \a9[0] );
  xor g33(n_88, \a14[0] , \a13[0] );
  xor g330(n_388, n_386, n_328);
  xor g331(n_389, n_106, \a10[0] );
  xor g333(n_391, n_389, n_361);
  xor g334(n_392, \a13[0] , \a11[0] );
  xor g336(n_394, n_392, n_368);
  xor g337(n_395, \a14[0] , \a12[0] );
  xor g339(n_397, n_395, n_321);
  xor g34(n_89, n_88, \a12[0] );
  xor g340(n_398, a15, \a13[0] );
  xor g342(n_83, n_398, n_327);
  xor g344(n_401, scr_out[20], scr_out[16]);
  xor g345(a15, n_298, n_401);
  xor g346(n_402, n_74, \a12[0] );
  xor g348(n_404, \a7[0] , n_402);
  xor g349(n_78, n_321, n_404);
  xor g35(n_90, n_89, \a9[0] );
  xor g4(n_72, scr_out[30], scr_out[21]);
  xor g41(n_95, n_74, \a13[0] );
  xor g42(n_96, n_95, \a10[0] );
  xor g48(n_101, n_74, \a11[0] );
  xor g49(n_102, n_101, \a10[0] );
  xor g5(\a14[0] , n_72, scr_out[17]);
  xor g54(n_106, a15, \a12[0] );
  xor g55(n_107, n_106, \a11[0] );
  xor g6(n_73, scr_out[31], scr_out[22]);
  xor g61(n_112, \a13[0] , \a12[0] );
  xor g7(\a13[0] , n_73, scr_out[18]);
  xor g8(\a12[0] , scr_out[23], scr_out[19]);
  xor g9(\a11[0] , scr_out[24], scr_out[20]);
  nor g22(n_422, scr_run, set, scr_init, reset);
  not g843(n_1151, reset);
  not g844(n_1152, scr_init);
  not g845(n_1153, scr_run);
  nor g846(n_423, scr_init, n_1153, reset, set);
  nor g847(n_424, n_1152, reset, set);
  nor g848(n_425, n_1151, set);
endmodule

