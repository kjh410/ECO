module top(out,reg_0,reg_1,fib,State,clk,rst,enb,reg_0_p,reg_1_p,fib_p,State_p);
	input clk, rst, enb;
	input [16:0]reg_0_p, reg_1_p, fib_p;
	input [2:0]State_p;
	output [16:0]out, reg_0, reg_1, fib;
	output [2:0]State;
	wire \g318/inv_sel0, \g318/w_0, \g318/w_1, \g312/inv_sel0, \g312/w_0, \g312/w_1, \g306/inv_sel0, \g306/w_0, \g306/w_1, \g300/inv_sel0, \g300/w_0, \g300/w_1, \g294/inv_sel0, \g294/w_0, \g294/w_1, \g288/inv_sel0, \g288/w_0, \g288/w_1, \g282/inv_sel0, \g282/w_0, \g282/w_1, \g276/inv_sel0, \g276/w_0, \g276/w_1, \g270/inv_sel0, \g270/w_0, \g270/w_1, \g264/inv_sel0, \g264/w_0, \g264/w_1, \g258/inv_sel0, \g258/w_0, \g258/w_1, \g252/inv_sel0, \g252/w_0, \g252/w_1, \g246/inv_sel0, \g246/w_0, \g246/w_1, \g240/inv_sel0, \g240/w_0, \g240/w_1, \g234/inv_sel0, \g234/w_0, \g234/w_1, \g228/inv_sel0, \g228/w_0, \g228/w_1, \g222/inv_sel0, \g222/w_0, \g222/w_1, \g216/inv_sel0, \g216/w_0, \g216/w_1, \g215/inv_sel0, \g215/w_0, \g215/w_1, \g214/inv_sel0, \g214/w_0, \g214/w_1, \g209/inv_sel0, \g209/w_0, \g209/w_1, \g208/inv_sel0, \g208/w_0, \g208/w_1, \g207/inv_sel0, \g207/w_0, \g207/w_1, \g202/inv_sel0, \g202/w_0, \g202/w_1, \g201/inv_sel0, \g201/w_0, \g201/w_1, \g200/inv_sel0, \g200/w_0, \g200/w_1, \g195/inv_sel0, \g195/w_0, \g195/w_1, \g194/inv_sel0, \g194/w_0, \g194/w_1, \g193/inv_sel0, \g193/w_0, \g193/w_1, \g188/inv_sel0, \g188/w_0, \g188/w_1, \g187/inv_sel0, \g187/w_0, \g187/w_1, \g186/inv_sel0, \g186/w_0, \g186/w_1, \g181/inv_sel0, \g181/w_0, \g181/w_1, \g180/inv_sel0, \g180/w_0, \g180/w_1, \g179/inv_sel0, \g179/w_0, \g179/w_1, \g174/inv_sel0, \g174/w_0, \g174/w_1, \g173/inv_sel0, \g173/w_0, \g173/w_1, \g172/inv_sel0, \g172/w_0, \g172/w_1, \g167/inv_sel0, \g167/w_0, \g167/w_1, \g166/inv_sel0, \g166/w_0, \g166/w_1, \g165/inv_sel0, \g165/w_0, \g165/w_1, \g160/inv_sel0, \g160/w_0, \g160/w_1, \g159/inv_sel0, \g159/w_0, \g159/w_1, \g158/inv_sel0, \g158/w_0, \g158/w_1, \g153/inv_sel0, \g153/w_0, \g153/w_1, \g152/inv_sel0, \g152/w_0, \g152/w_1, \g151/inv_sel0, \g151/w_0, \g151/w_1, \g146/inv_sel0, \g146/w_0, \g146/w_1, \g145/inv_sel0, \g145/w_0, \g145/w_1, \g144/inv_sel0, \g144/w_0, \g144/w_1, \g139/inv_sel0, \g139/w_0, \g139/w_1, \g138/inv_sel0, \g138/w_0, \g138/w_1, \g137/inv_sel0, \g137/w_0, \g137/w_1, \g132/inv_sel0, \g132/w_0, \g132/w_1, \g131/inv_sel0, \g131/w_0, \g131/w_1, \g130/inv_sel0, \g130/w_0, \g130/w_1, \g125/inv_sel0, \g125/w_0, \g125/w_1, \g124/inv_sel0, \g124/w_0, \g124/w_1, \g123/inv_sel0, \g123/w_0, \g123/w_1, \g118/inv_sel0, \g118/w_0, \g118/w_1, \g117/inv_sel0, \g117/w_0, \g117/w_1, \g116/inv_sel0, \g116/w_0, \g116/w_1, \g111/inv_sel0, \g111/w_0, \g111/w_1, \g110/inv_sel0, \g110/w_0, \g110/w_1, \g109/inv_sel0, \g109/w_0, \g109/w_1, \g104/inv_sel0, \g104/w_0, \g104/w_1, \g103/inv_sel0, \g103/w_0, \g103/w_1, \g102/inv_sel0, \g102/w_0, \g102/w_1, \g97/inv_sel0, \g97/w_0, \g97/w_1, \g91/inv_sel0, \g91/w_0, \g91/w_1, \g85/inv_sel0, \g85/w_0, \g85/w_1, \g79/inv_sel0, \g79/w_0, \g79/w_1, \g73/inv_sel0, \g73/w_0, \g73/w_1, \g67/inv_sel0, \g67/w_0, \g67/w_1, \g61/inv_sel0, \g61/w_0, \g61/w_1, \g55/inv_sel0, \g55/w_0, \g55/w_1, \g49/inv_sel0, \g49/w_0, \g49/w_1, \g43/inv_sel0, \g43/w_0, \g43/w_1, \g37/inv_sel0, \g37/w_0, \g37/w_1, \g31/inv_sel0, \g31/w_0, \g31/w_1, \g25/inv_sel0, \g25/w_0, \g25/w_1, \g1008/inv_sel0, \g1008/w_0, \g1008/w_1, \g13/inv_sel0, \g13/w_0, \g13/w_1, \g9/inv_sel0, \g9/w_0, \g9/w_1, \g3/inv_sel0, \g3/w_0, \g3/w_1, n_1708, n_1707, n_1706, n_1705, n_1704, n_1703, n_1702, n_1701, n_1700, n_1699, n_1698, n_1697, n_1422, n_1421, n_1420, n_1419, n_1418, n_1417, n_1416, n_1415, n_1414, n_1413, n_1412, n_1411, n_1410, n_1409, n_1408, n_1407, n_1406, n_1405, n_1404, n_1403, n_1402, n_1401, n_1400, n_1399, n_1398, n_1397, n_1396, n_1395, n_1394, n_1393, n_1392, n_1391, n_1390, n_1389, n_1388, n_1387, n_1220, n_1219, n_1218, n_1217, n_1216, n_1215, n_1214, n_1213, n_1212, n_1211, n_1210, n_1209, n_1208, n_1207, n_1206, n_1205, n_1203, n_1202, n_1201, n_1200, n_1199, n_1198, n_1197, n_1196, n_1195, n_1194, n_1193, n_1192, n_1191, n_1190, n_1189, n_1188, n_1187, n_1186, n_1185, n_1184, n_1183, n_1182, n_1181, n_1180, n_1179, n_1178, n_1177, n_1176, n_1175, n_1174, n_1173, n_1172, n_1171, n_1170, n_1169, n_1168, n_1167, n_1166, n_1165, n_1164, n_1163, n_1162, n_1161, n_1160, n_1159, n_1158, n_1157, n_1156, n_1155, n_1154, n_1153, n_1152, n_1151, n_1150, n_1149, n_1148, n_1147, n_1146, n_1145, n_1144, n_1143, n_1142, n_1141, n_1140, n_1139, n_1138, n_1137, n_1136, n_1135, n_1134, n_1133, n_1132, n_1131, n_1130, n_1129, n_1128, n_1127, n_1126, n_1125, n_1124, n_1123, n_1122, n_1121, n_1120, n_1119, n_1116, n_1115, n_881, n_598, n_595, n_594, n_395, n_393, n_392, n_391, n_390, n_387, n_386, n_385, n_384, n_381, n_380, n_379, n_378, n_375, n_374, n_373, n_372, n_369, n_368, n_367, n_366, n_363, n_362, n_361, n_360, n_357, n_356, n_355, n_354, n_351, n_350, n_349, n_348, n_345, n_344, n_343, n_342, n_339, n_338, n_337, n_336, n_333, n_332, n_331, n_330, n_327, n_326, n_325, n_324, n_321, n_320, n_319, n_318, n_315, n_314, n_313, n_312, n_309, n_308, n_307, n_306, n_303, n_302, n_301, n_300, n_297, n_296, n_295, n_294, n_291, n_290, n_289, n_288, n_287, n_286, n_282, n_281, n_280, n_279, n_278, n_277, n_273, n_272, n_271, n_270, n_269, n_268, n_264, n_263, n_262, n_261, n_260, n_259, n_255, n_254, n_253, n_252, n_251, n_250, n_246, n_245, n_244, n_243, n_242, n_241, n_237, n_236, n_235, n_234, n_233, n_232, n_228, n_227, n_226, n_208, n_207, n_206, n_205, n_201, n_200, n_199, n_198, n_197, n_196, n_192, n_191, n_190, n_189, n_188, n_187, n_183, n_182, n_181, n_180, n_179, n_178, n_174, n_173, n_172, n_171, n_170, n_169, n_165, n_164, n_163, n_162, n_161, n_160, n_156, n_155, n_154, n_153, n_152, n_151, n_147, n_146, n_145, n_144, n_143, n_142, n_138, n_137, n_136, n_135, n_130, n_129, n_128, n_127, n_122, n_121, n_120, n_119, n_114, n_113, n_112, n_111, n_106, n_105, n_104, n_103, n_98, n_97, n_96, n_95, n_90, n_89, n_88, n_87, n_81, n_77, n_73, n_69, n_65, n_61, n_57, n_53, n_49, n_45, n_41, n_37, n_33, n_29, n_25, n_21, n_17, n_14, n_12, n_10, n_8, add_107_31_n_225, add_107_31_n_222, add_107_31_n_220, add_107_31_n_217, add_107_31_n_214, add_107_31_n_211, add_107_31_n_209, add_107_31_n_205, add_107_31_n_202, add_107_31_n_200, add_107_31_n_196, add_107_31_n_191, add_107_31_n_189, add_107_31_n_188, add_107_31_n_187, add_107_31_n_185, add_107_31_n_184, add_107_31_n_182, add_107_31_n_181, add_107_31_n_178, add_107_31_n_176, add_107_31_n_169, add_107_31_n_166, add_107_31_n_164, add_107_31_n_162, add_107_31_n_160, add_107_31_n_158, add_107_31_n_154, add_107_31_n_152, add_107_31_n_151, add_107_31_n_147, add_107_31_n_142, add_107_31_n_139, add_107_31_n_134, add_107_31_n_132, add_107_31_n_130, add_107_31_n_129, add_107_31_n_124, add_107_31_n_122, add_107_31_n_120, add_107_31_n_119, add_107_31_n_114, add_107_31_n_112, add_107_31_n_110, add_107_31_n_109, add_107_31_n_108, add_107_31_n_106, add_107_31_n_103, add_107_31_n_102, add_107_31_n_100, add_107_31_n_99, add_107_31_n_98, add_107_31_n_97, add_107_31_n_96, add_107_31_n_94, add_107_31_n_93, add_107_31_n_92, add_107_31_n_91, add_107_31_n_90, add_107_31_n_88, add_107_31_n_87, add_107_31_n_86, add_107_31_n_85, add_107_31_n_84, add_107_31_n_82, add_107_31_n_81, add_107_31_n_80, add_107_31_n_79, add_107_31_n_78, add_107_31_n_76, add_107_31_n_75, add_107_31_n_74, add_107_31_n_73, add_107_31_n_72, add_107_31_n_70, add_107_31_n_69, add_107_31_n_68, add_107_31_n_67, add_107_31_n_66, add_107_31_n_64, add_107_31_n_63, add_107_31_n_62, add_107_31_n_61, add_107_31_n_59, add_107_31_n_56, add_107_31_n_53, enb, rst, clk;
	wire [2:0]State;
	wire [16:0]fib, reg_1, reg_0, out;
	wire [2:0]State_p;
	wire [16:0]fib_p, reg_1_p, reg_0_p;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, sub_wire1, w_eco5, sub_wire2, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, sub_wire3, w_eco15, w_eco16, w_eco17, w_eco18, sub_wire4, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, sub_wire5, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, sub_wire6, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, sub_wire7, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, sub_wire8, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, sub_wire9, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, sub_wire10, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, sub_wire11, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634, w_eco1635, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914, w_eco1915, w_eco1916, w_eco1917, w_eco1918, w_eco1919, w_eco1920, w_eco1921, w_eco1922, w_eco1923, w_eco1924, w_eco1925, w_eco1926, w_eco1927, w_eco1928, w_eco1929, w_eco1930, w_eco1931, w_eco1932, w_eco1933, w_eco1934, w_eco1935, w_eco1936, w_eco1937, w_eco1938, w_eco1939, w_eco1940, w_eco1941, w_eco1942, w_eco1943, w_eco1944, w_eco1945, w_eco1946, w_eco1947, w_eco1948, w_eco1949, w_eco1950, w_eco1951, w_eco1952, w_eco1953, w_eco1954, w_eco1955, w_eco1956, w_eco1957, w_eco1958, w_eco1959, w_eco1960, w_eco1961, w_eco1962, w_eco1963, w_eco1964, w_eco1965, w_eco1966, w_eco1967, w_eco1968, w_eco1969, w_eco1970, w_eco1971, w_eco1972, w_eco1973, w_eco1974, w_eco1975, w_eco1976, w_eco1977, w_eco1978, w_eco1979, w_eco1980, w_eco1981, w_eco1982, w_eco1983, w_eco1984, w_eco1985, w_eco1986, w_eco1987, w_eco1988, w_eco1989, w_eco1990, w_eco1991, w_eco1992, w_eco1993, w_eco1994, w_eco1995, w_eco1996, w_eco1997, w_eco1998, w_eco1999, w_eco2000, w_eco2001, w_eco2002, w_eco2003, w_eco2004, w_eco2005, w_eco2006, w_eco2007, w_eco2008, w_eco2009, w_eco2010, w_eco2011, w_eco2012, w_eco2013, w_eco2014, w_eco2015, w_eco2016, w_eco2017, w_eco2018, w_eco2019, w_eco2020, w_eco2021, w_eco2022, w_eco2023, w_eco2024, w_eco2025, w_eco2026, w_eco2027, w_eco2028, w_eco2029, w_eco2030, w_eco2031, w_eco2032, w_eco2033, w_eco2034, w_eco2035, w_eco2036, w_eco2037, w_eco2038, w_eco2039, w_eco2040, w_eco2041, w_eco2042, w_eco2043, w_eco2044, w_eco2045, w_eco2046, w_eco2047, w_eco2048, w_eco2049, w_eco2050, w_eco2051, w_eco2052, w_eco2053, w_eco2054, w_eco2055, w_eco2056, w_eco2057, w_eco2058, w_eco2059, w_eco2060, w_eco2061, w_eco2062, w_eco2063, w_eco2064, w_eco2065, w_eco2066, w_eco2067, w_eco2068, w_eco2069, w_eco2070, w_eco2071, w_eco2072, w_eco2073, w_eco2074, w_eco2075, w_eco2076, w_eco2077, w_eco2078, w_eco2079, w_eco2080, w_eco2081, w_eco2082, w_eco2083, w_eco2084, w_eco2085, w_eco2086, w_eco2087, w_eco2088, w_eco2089, w_eco2090, w_eco2091, w_eco2092, w_eco2093, w_eco2094, w_eco2095, w_eco2096, w_eco2097, w_eco2098, w_eco2099, w_eco2100, w_eco2101, w_eco2102, w_eco2103, w_eco2104, w_eco2105, w_eco2106, w_eco2107, w_eco2108, w_eco2109, w_eco2110, w_eco2111, w_eco2112, w_eco2113, w_eco2114, w_eco2115, w_eco2116, w_eco2117, w_eco2118, w_eco2119, w_eco2120, w_eco2121, w_eco2122, w_eco2123, w_eco2124, w_eco2125, w_eco2126, w_eco2127, w_eco2128, w_eco2129, w_eco2130, w_eco2131, w_eco2132, w_eco2133, w_eco2134, w_eco2135, w_eco2136, w_eco2137, w_eco2138, w_eco2139, w_eco2140, w_eco2141, w_eco2142, w_eco2143, w_eco2144, w_eco2145, w_eco2146, w_eco2147, w_eco2148, w_eco2149, w_eco2150, w_eco2151, w_eco2152, w_eco2153, w_eco2154, w_eco2155, w_eco2156, w_eco2157, w_eco2158, w_eco2159, w_eco2160, w_eco2161, w_eco2162, w_eco2163, w_eco2164, w_eco2165, w_eco2166, w_eco2167, w_eco2168, w_eco2169, w_eco2170, w_eco2171, w_eco2172, w_eco2173, w_eco2174, w_eco2175, w_eco2176, w_eco2177, w_eco2178, w_eco2179, w_eco2180, w_eco2181, w_eco2182, w_eco2183, w_eco2184, w_eco2185, w_eco2186, w_eco2187, w_eco2188, w_eco2189, w_eco2190, w_eco2191, w_eco2192, w_eco2193, w_eco2194, w_eco2195, w_eco2196, w_eco2197, w_eco2198, w_eco2199, w_eco2200, w_eco2201, w_eco2202, w_eco2203, w_eco2204, w_eco2205, w_eco2206, w_eco2207, w_eco2208, w_eco2209, w_eco2210, w_eco2211, w_eco2212, w_eco2213, w_eco2214, w_eco2215, w_eco2216, w_eco2217, w_eco2218, w_eco2219, w_eco2220, w_eco2221, w_eco2222, w_eco2223, w_eco2224, w_eco2225, w_eco2226, w_eco2227, w_eco2228, w_eco2229, w_eco2230, w_eco2231, w_eco2232, w_eco2233, w_eco2234, w_eco2235, w_eco2236, w_eco2237, w_eco2238, w_eco2239, w_eco2240, w_eco2241, w_eco2242, w_eco2243, w_eco2244, w_eco2245, w_eco2246, w_eco2247, w_eco2248, w_eco2249, w_eco2250, w_eco2251, w_eco2252, w_eco2253, w_eco2254, w_eco2255, w_eco2256, w_eco2257, w_eco2258, w_eco2259, w_eco2260, w_eco2261, w_eco2262, w_eco2263, w_eco2264, w_eco2265, w_eco2266, w_eco2267, w_eco2268, w_eco2269, w_eco2270, w_eco2271, w_eco2272, w_eco2273, w_eco2274, w_eco2275, w_eco2276, w_eco2277, w_eco2278, w_eco2279, w_eco2280, w_eco2281, w_eco2282, w_eco2283, w_eco2284, w_eco2285, w_eco2286, w_eco2287, w_eco2288, w_eco2289, w_eco2290, w_eco2291, w_eco2292, w_eco2293, w_eco2294, w_eco2295, w_eco2296, w_eco2297, w_eco2298, w_eco2299, w_eco2300, w_eco2301, w_eco2302, w_eco2303, w_eco2304, w_eco2305, w_eco2306, w_eco2307, w_eco2308, w_eco2309, w_eco2310, w_eco2311, w_eco2312, w_eco2313, w_eco2314, w_eco2315, w_eco2316, w_eco2317, w_eco2318, w_eco2319, w_eco2320, w_eco2321, w_eco2322, w_eco2323, w_eco2324, w_eco2325, w_eco2326, w_eco2327, w_eco2328, w_eco2329, w_eco2330, w_eco2331, w_eco2332, w_eco2333, w_eco2334, w_eco2335, w_eco2336, w_eco2337, w_eco2338, w_eco2339, w_eco2340, w_eco2341, w_eco2342, w_eco2343, w_eco2344, w_eco2345, w_eco2346, w_eco2347, w_eco2348, w_eco2349, w_eco2350, w_eco2351, w_eco2352, w_eco2353, w_eco2354, w_eco2355, w_eco2356, w_eco2357, w_eco2358, w_eco2359, w_eco2360, w_eco2361, w_eco2362, w_eco2363, w_eco2364, w_eco2365, w_eco2366, w_eco2367, w_eco2368, w_eco2369, w_eco2370, w_eco2371, w_eco2372, w_eco2373, w_eco2374, w_eco2375, w_eco2376, w_eco2377, w_eco2378, w_eco2379, w_eco2380, w_eco2381, w_eco2382, w_eco2383, w_eco2384, w_eco2385, w_eco2386, w_eco2387, w_eco2388, w_eco2389, w_eco2390, w_eco2391, w_eco2392, w_eco2393, w_eco2394, w_eco2395, w_eco2396, w_eco2397, w_eco2398, w_eco2399, w_eco2400, w_eco2401, w_eco2402, w_eco2403, w_eco2404, w_eco2405, w_eco2406, w_eco2407, w_eco2408, w_eco2409, w_eco2410, w_eco2411, w_eco2412, w_eco2413, w_eco2414, w_eco2415, w_eco2416, w_eco2417, w_eco2418, w_eco2419, w_eco2420, w_eco2421, w_eco2422, w_eco2423, w_eco2424, w_eco2425, w_eco2426, w_eco2427, w_eco2428, w_eco2429, w_eco2430, w_eco2431, w_eco2432, w_eco2433, w_eco2434, w_eco2435, w_eco2436, w_eco2437, w_eco2438, w_eco2439, w_eco2440, w_eco2441, w_eco2442, w_eco2443, w_eco2444, w_eco2445, w_eco2446, w_eco2447, w_eco2448, w_eco2449, w_eco2450, w_eco2451, w_eco2452, w_eco2453, w_eco2454, w_eco2455, w_eco2456, w_eco2457, w_eco2458, w_eco2459, w_eco2460, w_eco2461, w_eco2462, w_eco2463, w_eco2464, w_eco2465, w_eco2466, w_eco2467, w_eco2468, w_eco2469, w_eco2470, w_eco2471, w_eco2472, w_eco2473, w_eco2474, w_eco2475, w_eco2476, w_eco2477, w_eco2478, w_eco2479, w_eco2480, w_eco2481, w_eco2482, w_eco2483, w_eco2484, w_eco2485, w_eco2486, w_eco2487, w_eco2488, w_eco2489, w_eco2490, w_eco2491, w_eco2492, w_eco2493, w_eco2494, w_eco2495, w_eco2496, w_eco2497, w_eco2498, w_eco2499, w_eco2500, w_eco2501, w_eco2502, w_eco2503, w_eco2504, w_eco2505, w_eco2506, w_eco2507, w_eco2508, w_eco2509, w_eco2510, w_eco2511, w_eco2512, w_eco2513, w_eco2514, w_eco2515, w_eco2516, w_eco2517, w_eco2518, w_eco2519, w_eco2520, w_eco2521, w_eco2522, w_eco2523, w_eco2524, w_eco2525, w_eco2526, w_eco2527, w_eco2528, w_eco2529, w_eco2530, w_eco2531, w_eco2532, w_eco2533, w_eco2534, w_eco2535, w_eco2536, w_eco2537, w_eco2538, w_eco2539, w_eco2540, w_eco2541, w_eco2542, w_eco2543, w_eco2544, w_eco2545, w_eco2546, w_eco2547, w_eco2548, w_eco2549, w_eco2550, w_eco2551, w_eco2552, w_eco2553, w_eco2554, w_eco2555, w_eco2556, w_eco2557, w_eco2558, w_eco2559, w_eco2560, w_eco2561, w_eco2562, w_eco2563, w_eco2564, w_eco2565, w_eco2566, w_eco2567, w_eco2568, w_eco2569, w_eco2570, w_eco2571, w_eco2572, w_eco2573, w_eco2574, w_eco2575, w_eco2576, w_eco2577, w_eco2578, w_eco2579, w_eco2580, w_eco2581, w_eco2582, w_eco2583, w_eco2584, w_eco2585, w_eco2586, w_eco2587, w_eco2588, w_eco2589, w_eco2590, w_eco2591, w_eco2592, w_eco2593, w_eco2594, w_eco2595, w_eco2596, w_eco2597, w_eco2598, w_eco2599, w_eco2600, w_eco2601, w_eco2602, w_eco2603, w_eco2604, w_eco2605, w_eco2606, w_eco2607, w_eco2608, w_eco2609, w_eco2610, w_eco2611, w_eco2612, w_eco2613, w_eco2614, w_eco2615, w_eco2616, w_eco2617, w_eco2618, w_eco2619, w_eco2620, w_eco2621, w_eco2622, w_eco2623, w_eco2624, w_eco2625, w_eco2626, w_eco2627, w_eco2628, w_eco2629, w_eco2630, w_eco2631, w_eco2632, w_eco2633, w_eco2634, w_eco2635, w_eco2636, w_eco2637, w_eco2638, w_eco2639, w_eco2640, w_eco2641, w_eco2642, w_eco2643, w_eco2644, w_eco2645, w_eco2646, w_eco2647, w_eco2648, w_eco2649, w_eco2650, w_eco2651, w_eco2652, w_eco2653, w_eco2654, w_eco2655, w_eco2656, w_eco2657, w_eco2658, w_eco2659, w_eco2660, w_eco2661, w_eco2662, w_eco2663, w_eco2664, w_eco2665, w_eco2666, w_eco2667, w_eco2668, w_eco2669, w_eco2670, w_eco2671, w_eco2672, w_eco2673, w_eco2674, w_eco2675, w_eco2676, w_eco2677, w_eco2678, w_eco2679, w_eco2680, w_eco2681, w_eco2682, w_eco2683, w_eco2684, w_eco2685, w_eco2686, w_eco2687, w_eco2688, w_eco2689, w_eco2690, w_eco2691, w_eco2692, w_eco2693, w_eco2694, w_eco2695, w_eco2696, w_eco2697, w_eco2698, w_eco2699, w_eco2700, w_eco2701, w_eco2702, w_eco2703, w_eco2704, w_eco2705, w_eco2706, w_eco2707, w_eco2708, w_eco2709, w_eco2710, w_eco2711, w_eco2712, w_eco2713, w_eco2714, w_eco2715, w_eco2716, w_eco2717, w_eco2718, w_eco2719, w_eco2720, w_eco2721, w_eco2722, w_eco2723, w_eco2724, w_eco2725, w_eco2726, w_eco2727, w_eco2728, w_eco2729, w_eco2730, w_eco2731, w_eco2732, w_eco2733, w_eco2734, w_eco2735, w_eco2736, w_eco2737, w_eco2738, w_eco2739, w_eco2740, w_eco2741, w_eco2742, w_eco2743, w_eco2744, w_eco2745, w_eco2746, w_eco2747, w_eco2748, w_eco2749, w_eco2750, w_eco2751, w_eco2752, w_eco2753, w_eco2754, w_eco2755, w_eco2756, w_eco2757, w_eco2758, w_eco2759, w_eco2760, w_eco2761, w_eco2762, w_eco2763, w_eco2764, w_eco2765, w_eco2766, w_eco2767, w_eco2768, w_eco2769, w_eco2770, w_eco2771, w_eco2772, w_eco2773, w_eco2774, w_eco2775, w_eco2776, w_eco2777, w_eco2778, w_eco2779, w_eco2780, w_eco2781, w_eco2782, w_eco2783, w_eco2784, w_eco2785, w_eco2786, w_eco2787, w_eco2788, w_eco2789, w_eco2790, w_eco2791, w_eco2792, w_eco2793, w_eco2794, w_eco2795, w_eco2796, w_eco2797, w_eco2798, w_eco2799, w_eco2800, w_eco2801, w_eco2802, w_eco2803, w_eco2804, w_eco2805, w_eco2806, w_eco2807, w_eco2808, w_eco2809, w_eco2810, w_eco2811, w_eco2812, w_eco2813, w_eco2814, w_eco2815, w_eco2816, w_eco2817, w_eco2818, w_eco2819, w_eco2820, w_eco2821, w_eco2822, w_eco2823, w_eco2824, w_eco2825, w_eco2826, w_eco2827, w_eco2828, w_eco2829, w_eco2830, w_eco2831, w_eco2832, w_eco2833, w_eco2834, w_eco2835, w_eco2836, w_eco2837, w_eco2838, w_eco2839, w_eco2840, w_eco2841, w_eco2842, w_eco2843, w_eco2844, w_eco2845, w_eco2846, w_eco2847, w_eco2848, w_eco2849, w_eco2850, w_eco2851, w_eco2852, w_eco2853, w_eco2854, w_eco2855, w_eco2856, w_eco2857, w_eco2858, w_eco2859, w_eco2860, w_eco2861, w_eco2862, w_eco2863, w_eco2864, w_eco2865, w_eco2866, w_eco2867, w_eco2868, w_eco2869, w_eco2870, w_eco2871, w_eco2872, w_eco2873, w_eco2874, w_eco2875, w_eco2876, w_eco2877, w_eco2878, w_eco2879, w_eco2880, w_eco2881, w_eco2882, w_eco2883, w_eco2884, w_eco2885, w_eco2886, w_eco2887, w_eco2888, w_eco2889, w_eco2890, w_eco2891, w_eco2892, w_eco2893, w_eco2894, w_eco2895, w_eco2896, w_eco2897, w_eco2898, w_eco2899, w_eco2900, w_eco2901, w_eco2902, w_eco2903, w_eco2904, w_eco2905, w_eco2906, w_eco2907, w_eco2908, w_eco2909, w_eco2910, w_eco2911, w_eco2912, w_eco2913, w_eco2914, w_eco2915, w_eco2916, w_eco2917, w_eco2918, w_eco2919, w_eco2920, w_eco2921, w_eco2922, w_eco2923, w_eco2924, w_eco2925, w_eco2926, w_eco2927, w_eco2928, w_eco2929, w_eco2930, w_eco2931, w_eco2932, w_eco2933, w_eco2934, w_eco2935, w_eco2936, w_eco2937, w_eco2938, w_eco2939, w_eco2940, w_eco2941, w_eco2942, w_eco2943, w_eco2944, w_eco2945, w_eco2946, w_eco2947, w_eco2948, w_eco2949, w_eco2950, w_eco2951, w_eco2952, w_eco2953, w_eco2954, w_eco2955, w_eco2956, w_eco2957, w_eco2958, w_eco2959, w_eco2960, w_eco2961, w_eco2962, w_eco2963, w_eco2964, w_eco2965, w_eco2966, w_eco2967, w_eco2968, w_eco2969, w_eco2970, w_eco2971, w_eco2972, w_eco2973, w_eco2974, w_eco2975, w_eco2976, w_eco2977, w_eco2978, w_eco2979, w_eco2980, w_eco2981, w_eco2982, w_eco2983, w_eco2984, w_eco2985, w_eco2986, w_eco2987, w_eco2988, w_eco2989, w_eco2990, w_eco2991, w_eco2992, w_eco2993, w_eco2994, w_eco2995, w_eco2996, w_eco2997, w_eco2998, w_eco2999, w_eco3000, w_eco3001, w_eco3002, w_eco3003, w_eco3004, w_eco3005, w_eco3006, w_eco3007, w_eco3008, w_eco3009, w_eco3010, w_eco3011, w_eco3012, w_eco3013, w_eco3014, w_eco3015, w_eco3016, w_eco3017, w_eco3018, w_eco3019, w_eco3020, w_eco3021, w_eco3022, w_eco3023, w_eco3024, w_eco3025, w_eco3026, w_eco3027, w_eco3028, w_eco3029, w_eco3030, w_eco3031, w_eco3032, w_eco3033, w_eco3034, w_eco3035, w_eco3036, w_eco3037, w_eco3038, w_eco3039, w_eco3040, w_eco3041, w_eco3042, w_eco3043, w_eco3044, w_eco3045, w_eco3046, w_eco3047, w_eco3048, w_eco3049, w_eco3050, w_eco3051, w_eco3052, w_eco3053, w_eco3054, w_eco3055, w_eco3056, w_eco3057, w_eco3058, w_eco3059, w_eco3060, w_eco3061, w_eco3062, w_eco3063, w_eco3064, w_eco3065, w_eco3066, w_eco3067, w_eco3068, w_eco3069, w_eco3070, w_eco3071, w_eco3072, w_eco3073, w_eco3074, w_eco3075, w_eco3076, w_eco3077, w_eco3078, w_eco3079, w_eco3080, w_eco3081, w_eco3082, w_eco3083, w_eco3084, w_eco3085, w_eco3086, w_eco3087, w_eco3088, w_eco3089, w_eco3090, w_eco3091, w_eco3092, w_eco3093, w_eco3094, w_eco3095, w_eco3096, w_eco3097, w_eco3098, w_eco3099, w_eco3100, w_eco3101, w_eco3102, w_eco3103, w_eco3104, w_eco3105, w_eco3106, w_eco3107, w_eco3108, w_eco3109, w_eco3110, w_eco3111, w_eco3112, w_eco3113, w_eco3114, w_eco3115, w_eco3116, w_eco3117, w_eco3118, w_eco3119, w_eco3120, w_eco3121, w_eco3122, w_eco3123, w_eco3124, w_eco3125, w_eco3126, w_eco3127, w_eco3128, w_eco3129, w_eco3130, w_eco3131, w_eco3132, w_eco3133, w_eco3134, w_eco3135, w_eco3136, w_eco3137, w_eco3138, w_eco3139, w_eco3140, w_eco3141, w_eco3142, w_eco3143, w_eco3144, w_eco3145, w_eco3146, w_eco3147, w_eco3148, w_eco3149, w_eco3150, w_eco3151, w_eco3152, w_eco3153, w_eco3154, w_eco3155, w_eco3156, w_eco3157, w_eco3158, w_eco3159, w_eco3160, w_eco3161, w_eco3162, w_eco3163, w_eco3164, w_eco3165, w_eco3166, w_eco3167, w_eco3168, w_eco3169, w_eco3170, w_eco3171, w_eco3172, w_eco3173, w_eco3174, w_eco3175, w_eco3176, w_eco3177, w_eco3178, w_eco3179, w_eco3180, w_eco3181, w_eco3182, w_eco3183, w_eco3184, w_eco3185, w_eco3186, w_eco3187, w_eco3188, w_eco3189, w_eco3190, w_eco3191, w_eco3192, w_eco3193, w_eco3194, w_eco3195, w_eco3196, w_eco3197, w_eco3198, w_eco3199, w_eco3200, w_eco3201, w_eco3202, w_eco3203, w_eco3204, w_eco3205, w_eco3206, w_eco3207, w_eco3208, w_eco3209, w_eco3210, w_eco3211, w_eco3212, w_eco3213, w_eco3214, w_eco3215, w_eco3216, w_eco3217, w_eco3218, w_eco3219, w_eco3220, w_eco3221, w_eco3222, w_eco3223, w_eco3224, w_eco3225, w_eco3226, w_eco3227, w_eco3228, w_eco3229, w_eco3230, w_eco3231, w_eco3232, w_eco3233, w_eco3234, w_eco3235, w_eco3236, w_eco3237, w_eco3238, w_eco3239, w_eco3240, w_eco3241, w_eco3242, w_eco3243, w_eco3244, w_eco3245, w_eco3246, w_eco3247, w_eco3248, w_eco3249, w_eco3250, w_eco3251, w_eco3252, w_eco3253, w_eco3254, w_eco3255, w_eco3256, w_eco3257, w_eco3258, w_eco3259, w_eco3260, w_eco3261, w_eco3262, w_eco3263, w_eco3264, w_eco3265, w_eco3266, w_eco3267, w_eco3268, w_eco3269, w_eco3270, w_eco3271, w_eco3272, w_eco3273, w_eco3274, w_eco3275, w_eco3276, w_eco3277, w_eco3278, w_eco3279, w_eco3280, w_eco3281, w_eco3282, w_eco3283, w_eco3284, w_eco3285, w_eco3286, w_eco3287, w_eco3288, w_eco3289, w_eco3290, w_eco3291, w_eco3292, w_eco3293, w_eco3294, w_eco3295, w_eco3296, w_eco3297, w_eco3298, w_eco3299, w_eco3300, w_eco3301, w_eco3302, w_eco3303, w_eco3304, w_eco3305, w_eco3306, w_eco3307, w_eco3308, w_eco3309, w_eco3310, w_eco3311, w_eco3312, w_eco3313, w_eco3314, w_eco3315, w_eco3316, w_eco3317, w_eco3318, w_eco3319, w_eco3320, w_eco3321, w_eco3322, w_eco3323, w_eco3324, w_eco3325, w_eco3326, w_eco3327, w_eco3328, w_eco3329, w_eco3330, w_eco3331, w_eco3332, w_eco3333, w_eco3334, w_eco3335, w_eco3336, w_eco3337, w_eco3338, w_eco3339, w_eco3340, w_eco3341, w_eco3342, w_eco3343, w_eco3344, w_eco3345, w_eco3346, w_eco3347, w_eco3348, w_eco3349, w_eco3350, w_eco3351, w_eco3352, w_eco3353, w_eco3354, w_eco3355, w_eco3356, w_eco3357, w_eco3358, w_eco3359, w_eco3360, w_eco3361, w_eco3362, w_eco3363, w_eco3364, w_eco3365, w_eco3366, w_eco3367, w_eco3368, w_eco3369, w_eco3370, w_eco3371, w_eco3372, w_eco3373, w_eco3374, w_eco3375, w_eco3376, w_eco3377, w_eco3378, w_eco3379, w_eco3380, w_eco3381, w_eco3382, w_eco3383, w_eco3384, w_eco3385, w_eco3386, w_eco3387, w_eco3388, w_eco3389, w_eco3390, w_eco3391, w_eco3392, w_eco3393, w_eco3394, w_eco3395, w_eco3396, w_eco3397, w_eco3398, w_eco3399, w_eco3400, w_eco3401, w_eco3402, w_eco3403, w_eco3404, w_eco3405, w_eco3406, w_eco3407, w_eco3408, w_eco3409, w_eco3410, w_eco3411, w_eco3412, w_eco3413, w_eco3414, w_eco3415, w_eco3416, w_eco3417, w_eco3418, w_eco3419, w_eco3420, w_eco3421, w_eco3422, w_eco3423, w_eco3424, w_eco3425, w_eco3426, w_eco3427, w_eco3428, w_eco3429, w_eco3430, w_eco3431, w_eco3432, w_eco3433, w_eco3434, w_eco3435, w_eco3436, w_eco3437, w_eco3438, w_eco3439, w_eco3440, w_eco3441, w_eco3442, w_eco3443, w_eco3444, w_eco3445, w_eco3446, w_eco3447, w_eco3448, w_eco3449, w_eco3450, w_eco3451, w_eco3452, w_eco3453, w_eco3454, w_eco3455, w_eco3456, w_eco3457, w_eco3458, w_eco3459, w_eco3460, w_eco3461, w_eco3462, w_eco3463, w_eco3464, w_eco3465, w_eco3466, w_eco3467, w_eco3468, w_eco3469, w_eco3470, w_eco3471, w_eco3472, w_eco3473, w_eco3474, w_eco3475, w_eco3476, w_eco3477, w_eco3478, w_eco3479, w_eco3480, w_eco3481, w_eco3482, w_eco3483, w_eco3484, w_eco3485, w_eco3486, w_eco3487, w_eco3488, w_eco3489, w_eco3490, w_eco3491, w_eco3492, w_eco3493, w_eco3494, w_eco3495, w_eco3496, w_eco3497, w_eco3498, w_eco3499, w_eco3500, w_eco3501, w_eco3502, w_eco3503, w_eco3504, w_eco3505, w_eco3506, w_eco3507, w_eco3508, w_eco3509, w_eco3510, w_eco3511, w_eco3512, w_eco3513, w_eco3514, w_eco3515, w_eco3516, w_eco3517, w_eco3518, w_eco3519, w_eco3520, w_eco3521, w_eco3522, w_eco3523, w_eco3524, w_eco3525, w_eco3526, w_eco3527, w_eco3528, w_eco3529, w_eco3530, w_eco3531, w_eco3532, w_eco3533, w_eco3534, w_eco3535, w_eco3536, w_eco3537, w_eco3538, w_eco3539, w_eco3540, w_eco3541, w_eco3542, w_eco3543, w_eco3544, w_eco3545, w_eco3546, w_eco3547, w_eco3548, w_eco3549, w_eco3550, w_eco3551, w_eco3552, w_eco3553, w_eco3554, w_eco3555, w_eco3556, w_eco3557, w_eco3558, w_eco3559, w_eco3560, w_eco3561, w_eco3562, w_eco3563, w_eco3564, w_eco3565, w_eco3566, w_eco3567, w_eco3568, w_eco3569, w_eco3570, w_eco3571, w_eco3572, w_eco3573, w_eco3574, w_eco3575, w_eco3576, w_eco3577, w_eco3578, w_eco3579, w_eco3580, w_eco3581, w_eco3582, w_eco3583, w_eco3584, w_eco3585, w_eco3586, w_eco3587, w_eco3588, w_eco3589, w_eco3590, w_eco3591, w_eco3592, w_eco3593, w_eco3594, w_eco3595, w_eco3596, w_eco3597, w_eco3598, w_eco3599, w_eco3600, w_eco3601, w_eco3602, w_eco3603, w_eco3604, w_eco3605, w_eco3606, w_eco3607, w_eco3608, w_eco3609, w_eco3610, w_eco3611, w_eco3612, w_eco3613, w_eco3614, w_eco3615, w_eco3616, w_eco3617, w_eco3618, w_eco3619, w_eco3620, w_eco3621, w_eco3622, w_eco3623, w_eco3624, w_eco3625, w_eco3626, w_eco3627, w_eco3628, w_eco3629, w_eco3630, w_eco3631, w_eco3632, w_eco3633, w_eco3634, w_eco3635, w_eco3636, w_eco3637, w_eco3638, w_eco3639, w_eco3640, w_eco3641, w_eco3642, w_eco3643, w_eco3644, w_eco3645, w_eco3646, w_eco3647, w_eco3648, w_eco3649, w_eco3650, w_eco3651, w_eco3652, w_eco3653, w_eco3654, w_eco3655, w_eco3656, w_eco3657, w_eco3658, w_eco3659, w_eco3660, w_eco3661, w_eco3662, w_eco3663, w_eco3664, w_eco3665, w_eco3666, w_eco3667, w_eco3668, w_eco3669, w_eco3670, w_eco3671, w_eco3672, w_eco3673, w_eco3674, w_eco3675, w_eco3676, w_eco3677, w_eco3678, w_eco3679, w_eco3680, w_eco3681, w_eco3682, w_eco3683, w_eco3684, w_eco3685, w_eco3686, w_eco3687, w_eco3688, w_eco3689, w_eco3690, w_eco3691, w_eco3692, w_eco3693, w_eco3694, w_eco3695, w_eco3696, w_eco3697, w_eco3698, w_eco3699, w_eco3700, w_eco3701, w_eco3702, w_eco3703, w_eco3704, w_eco3705, w_eco3706, w_eco3707, w_eco3708, w_eco3709, w_eco3710, w_eco3711, w_eco3712, w_eco3713, w_eco3714, w_eco3715, w_eco3716, w_eco3717, w_eco3718, w_eco3719, w_eco3720, w_eco3721, w_eco3722, w_eco3723, w_eco3724, w_eco3725, w_eco3726, w_eco3727, w_eco3728, w_eco3729, w_eco3730, w_eco3731, w_eco3732, w_eco3733, w_eco3734, w_eco3735, w_eco3736, w_eco3737, w_eco3738, w_eco3739, w_eco3740, w_eco3741, w_eco3742, w_eco3743, w_eco3744, w_eco3745, w_eco3746, w_eco3747, w_eco3748, w_eco3749, w_eco3750, w_eco3751, w_eco3752, w_eco3753, w_eco3754, w_eco3755, w_eco3756, w_eco3757, w_eco3758, w_eco3759, w_eco3760, w_eco3761, w_eco3762, w_eco3763, w_eco3764, w_eco3765, w_eco3766, w_eco3767, w_eco3768, w_eco3769, w_eco3770, w_eco3771, w_eco3772, w_eco3773, w_eco3774, w_eco3775, w_eco3776, w_eco3777, w_eco3778, w_eco3779, w_eco3780, w_eco3781, w_eco3782, w_eco3783, w_eco3784, w_eco3785, w_eco3786, w_eco3787, w_eco3788, w_eco3789, w_eco3790, w_eco3791, w_eco3792, w_eco3793, w_eco3794, w_eco3795, w_eco3796, w_eco3797, w_eco3798, w_eco3799, w_eco3800, w_eco3801, w_eco3802, w_eco3803, w_eco3804, w_eco3805, w_eco3806, w_eco3807, w_eco3808, w_eco3809, w_eco3810, w_eco3811, w_eco3812, w_eco3813, w_eco3814, w_eco3815, w_eco3816, w_eco3817, w_eco3818, w_eco3819, w_eco3820, w_eco3821, w_eco3822, w_eco3823, w_eco3824, w_eco3825, w_eco3826, w_eco3827, w_eco3828, w_eco3829, w_eco3830, w_eco3831, w_eco3832, w_eco3833, w_eco3834, w_eco3835, w_eco3836, w_eco3837, w_eco3838, w_eco3839, w_eco3840, w_eco3841, w_eco3842, w_eco3843, w_eco3844, w_eco3845, w_eco3846, w_eco3847, w_eco3848, w_eco3849, w_eco3850, w_eco3851, w_eco3852, w_eco3853, w_eco3854, w_eco3855, w_eco3856, w_eco3857, w_eco3858, w_eco3859, w_eco3860, w_eco3861, w_eco3862, w_eco3863, w_eco3864, w_eco3865, w_eco3866, w_eco3867, w_eco3868, w_eco3869, w_eco3870, w_eco3871, w_eco3872, w_eco3873, w_eco3874, w_eco3875, w_eco3876, w_eco3877, w_eco3878, w_eco3879, w_eco3880, w_eco3881, w_eco3882, w_eco3883, w_eco3884, w_eco3885, w_eco3886, w_eco3887, w_eco3888, w_eco3889, w_eco3890, w_eco3891, w_eco3892, w_eco3893, w_eco3894, w_eco3895, w_eco3896, w_eco3897, w_eco3898, w_eco3899, w_eco3900, w_eco3901, w_eco3902, w_eco3903, w_eco3904, w_eco3905, w_eco3906, w_eco3907, w_eco3908, w_eco3909, w_eco3910, w_eco3911, w_eco3912, w_eco3913, w_eco3914, w_eco3915, w_eco3916, w_eco3917, w_eco3918, w_eco3919, w_eco3920, w_eco3921, w_eco3922, w_eco3923, w_eco3924, w_eco3925, w_eco3926, w_eco3927, w_eco3928, w_eco3929, w_eco3930, w_eco3931, w_eco3932, w_eco3933, w_eco3934, w_eco3935, w_eco3936, w_eco3937, w_eco3938, w_eco3939, w_eco3940, w_eco3941, w_eco3942, w_eco3943, w_eco3944, w_eco3945, w_eco3946, w_eco3947, w_eco3948, w_eco3949, w_eco3950, w_eco3951, w_eco3952, w_eco3953, w_eco3954, w_eco3955, w_eco3956, w_eco3957, w_eco3958, w_eco3959, w_eco3960, w_eco3961, w_eco3962, w_eco3963, w_eco3964, w_eco3965, w_eco3966, w_eco3967, w_eco3968, w_eco3969, w_eco3970, w_eco3971, w_eco3972, w_eco3973, w_eco3974, w_eco3975, w_eco3976, w_eco3977, w_eco3978, w_eco3979, w_eco3980, w_eco3981, w_eco3982, w_eco3983, w_eco3984, w_eco3985, w_eco3986, w_eco3987, w_eco3988, w_eco3989, w_eco3990, w_eco3991, w_eco3992, w_eco3993, w_eco3994, w_eco3995, w_eco3996, w_eco3997, w_eco3998, w_eco3999, w_eco4000, w_eco4001, w_eco4002, w_eco4003, w_eco4004, w_eco4005, w_eco4006, w_eco4007, w_eco4008, w_eco4009, w_eco4010, w_eco4011, w_eco4012, w_eco4013, w_eco4014, w_eco4015, w_eco4016, w_eco4017, w_eco4018, w_eco4019, w_eco4020, w_eco4021, w_eco4022, w_eco4023, w_eco4024, w_eco4025, w_eco4026, w_eco4027, w_eco4028, w_eco4029, w_eco4030, w_eco4031, w_eco4032, w_eco4033, w_eco4034, w_eco4035, w_eco4036, w_eco4037, w_eco4038, w_eco4039, w_eco4040, w_eco4041, w_eco4042, w_eco4043, w_eco4044, w_eco4045, w_eco4046, w_eco4047, w_eco4048, w_eco4049, w_eco4050, w_eco4051, w_eco4052, w_eco4053, w_eco4054, w_eco4055, w_eco4056, w_eco4057, w_eco4058, w_eco4059, w_eco4060, w_eco4061, w_eco4062, w_eco4063, w_eco4064, w_eco4065, w_eco4066, w_eco4067, w_eco4068, w_eco4069, w_eco4070, w_eco4071, w_eco4072, w_eco4073, w_eco4074, w_eco4075, w_eco4076, w_eco4077, w_eco4078, w_eco4079, w_eco4080, w_eco4081, w_eco4082, w_eco4083, w_eco4084, w_eco4085, w_eco4086, w_eco4087, w_eco4088, w_eco4089, w_eco4090, w_eco4091, w_eco4092, w_eco4093, w_eco4094, w_eco4095, w_eco4096, w_eco4097, w_eco4098, w_eco4099, w_eco4100, w_eco4101, w_eco4102, w_eco4103, w_eco4104, w_eco4105, w_eco4106, w_eco4107, w_eco4108, w_eco4109, w_eco4110, w_eco4111, w_eco4112, w_eco4113, w_eco4114, w_eco4115, w_eco4116, w_eco4117, w_eco4118, w_eco4119, w_eco4120, w_eco4121, w_eco4122, w_eco4123, w_eco4124, w_eco4125, w_eco4126, w_eco4127, w_eco4128, w_eco4129, w_eco4130, w_eco4131, w_eco4132, w_eco4133, w_eco4134, w_eco4135, w_eco4136, w_eco4137, w_eco4138, w_eco4139, w_eco4140, w_eco4141, w_eco4142, w_eco4143, w_eco4144, w_eco4145, w_eco4146, w_eco4147, w_eco4148, w_eco4149, w_eco4150, w_eco4151, w_eco4152, w_eco4153, w_eco4154, w_eco4155, w_eco4156, w_eco4157, w_eco4158, w_eco4159, w_eco4160, w_eco4161, w_eco4162, w_eco4163, w_eco4164, w_eco4165, w_eco4166, w_eco4167, w_eco4168, w_eco4169, w_eco4170, w_eco4171, w_eco4172, w_eco4173, w_eco4174, w_eco4175, w_eco4176, w_eco4177, w_eco4178, w_eco4179, w_eco4180, w_eco4181, w_eco4182, w_eco4183, w_eco4184, w_eco4185, w_eco4186, w_eco4187, w_eco4188, w_eco4189, w_eco4190, w_eco4191, w_eco4192, w_eco4193, w_eco4194, w_eco4195, w_eco4196, w_eco4197, w_eco4198, w_eco4199, w_eco4200, w_eco4201, w_eco4202, w_eco4203, w_eco4204, w_eco4205, w_eco4206, w_eco4207, w_eco4208, w_eco4209, w_eco4210, w_eco4211, w_eco4212, w_eco4213, w_eco4214, w_eco4215, w_eco4216, w_eco4217, w_eco4218, w_eco4219, w_eco4220, w_eco4221, w_eco4222, w_eco4223, w_eco4224, w_eco4225, w_eco4226, w_eco4227, w_eco4228, w_eco4229, w_eco4230, w_eco4231, w_eco4232, w_eco4233, w_eco4234, w_eco4235, w_eco4236, w_eco4237, w_eco4238, w_eco4239, w_eco4240, w_eco4241, w_eco4242, w_eco4243, w_eco4244, w_eco4245, w_eco4246, w_eco4247, w_eco4248, w_eco4249, w_eco4250, w_eco4251, w_eco4252, w_eco4253, w_eco4254, w_eco4255, w_eco4256, w_eco4257, w_eco4258, w_eco4259, w_eco4260, w_eco4261, w_eco4262, w_eco4263, w_eco4264, w_eco4265, w_eco4266, w_eco4267, w_eco4268, w_eco4269, w_eco4270, w_eco4271, w_eco4272, w_eco4273, w_eco4274, w_eco4275, w_eco4276, w_eco4277, w_eco4278, w_eco4279, w_eco4280, w_eco4281, w_eco4282, w_eco4283, w_eco4284, w_eco4285, w_eco4286, w_eco4287, w_eco4288, w_eco4289, w_eco4290, w_eco4291, w_eco4292, w_eco4293, w_eco4294, w_eco4295, w_eco4296, w_eco4297, w_eco4298, w_eco4299, w_eco4300, w_eco4301, w_eco4302, w_eco4303, w_eco4304, w_eco4305, w_eco4306, w_eco4307, w_eco4308, w_eco4309, w_eco4310, w_eco4311, w_eco4312, w_eco4313, w_eco4314, w_eco4315, w_eco4316, w_eco4317, w_eco4318, w_eco4319, w_eco4320, w_eco4321, w_eco4322, w_eco4323, w_eco4324, w_eco4325, w_eco4326, w_eco4327, w_eco4328, w_eco4329, w_eco4330, w_eco4331, w_eco4332, w_eco4333, w_eco4334, w_eco4335, w_eco4336, w_eco4337, w_eco4338, w_eco4339, w_eco4340, w_eco4341, w_eco4342, w_eco4343, w_eco4344, w_eco4345, w_eco4346, w_eco4347, w_eco4348, w_eco4349, w_eco4350, w_eco4351, w_eco4352, w_eco4353, w_eco4354, w_eco4355, w_eco4356, w_eco4357, w_eco4358, w_eco4359, w_eco4360, w_eco4361, w_eco4362, w_eco4363, w_eco4364, w_eco4365, w_eco4366, w_eco4367, w_eco4368, w_eco4369, w_eco4370, w_eco4371, w_eco4372, w_eco4373, w_eco4374, w_eco4375, w_eco4376, w_eco4377, w_eco4378, w_eco4379, w_eco4380, w_eco4381, w_eco4382, w_eco4383, w_eco4384, w_eco4385, w_eco4386, w_eco4387, w_eco4388, w_eco4389, w_eco4390, w_eco4391, w_eco4392, w_eco4393, w_eco4394, w_eco4395, w_eco4396, w_eco4397, w_eco4398, w_eco4399, w_eco4400, w_eco4401, w_eco4402, w_eco4403, w_eco4404, w_eco4405, w_eco4406, w_eco4407, w_eco4408, w_eco4409, w_eco4410, w_eco4411, w_eco4412, w_eco4413, w_eco4414, w_eco4415, w_eco4416, w_eco4417, w_eco4418, w_eco4419, w_eco4420, w_eco4421, w_eco4422, w_eco4423, w_eco4424, w_eco4425, w_eco4426, w_eco4427, w_eco4428, w_eco4429, w_eco4430, w_eco4431, w_eco4432, w_eco4433, w_eco4434, w_eco4435, w_eco4436, w_eco4437, w_eco4438, w_eco4439, w_eco4440, w_eco4441, w_eco4442, w_eco4443, w_eco4444, w_eco4445, w_eco4446, w_eco4447, w_eco4448, w_eco4449, w_eco4450, w_eco4451, w_eco4452, w_eco4453, w_eco4454, w_eco4455, w_eco4456, w_eco4457, w_eco4458, w_eco4459, w_eco4460, w_eco4461, w_eco4462, w_eco4463, w_eco4464, w_eco4465, w_eco4466, w_eco4467, w_eco4468, w_eco4469, w_eco4470, w_eco4471, w_eco4472, w_eco4473, w_eco4474, w_eco4475, w_eco4476, w_eco4477, w_eco4478, w_eco4479, w_eco4480, w_eco4481, w_eco4482, w_eco4483, w_eco4484, w_eco4485, w_eco4486, w_eco4487, w_eco4488, w_eco4489, w_eco4490, w_eco4491, w_eco4492, w_eco4493, w_eco4494, w_eco4495, w_eco4496, w_eco4497, w_eco4498, w_eco4499, w_eco4500, w_eco4501, w_eco4502, w_eco4503, w_eco4504, w_eco4505, w_eco4506, w_eco4507, w_eco4508, w_eco4509, w_eco4510, w_eco4511, w_eco4512, w_eco4513, w_eco4514, w_eco4515, w_eco4516, w_eco4517, w_eco4518, w_eco4519, w_eco4520, w_eco4521, w_eco4522, w_eco4523, w_eco4524, w_eco4525, w_eco4526, w_eco4527, w_eco4528, w_eco4529, w_eco4530, w_eco4531, w_eco4532, w_eco4533, w_eco4534, w_eco4535, w_eco4536, w_eco4537, w_eco4538, w_eco4539, w_eco4540, w_eco4541, w_eco4542, w_eco4543, w_eco4544, w_eco4545, w_eco4546, w_eco4547, w_eco4548, w_eco4549, w_eco4550, w_eco4551, w_eco4552, w_eco4553, w_eco4554, w_eco4555, w_eco4556, w_eco4557, w_eco4558, w_eco4559, w_eco4560, w_eco4561, w_eco4562, w_eco4563, w_eco4564, w_eco4565, w_eco4566, w_eco4567, w_eco4568, w_eco4569, w_eco4570, w_eco4571, w_eco4572, w_eco4573, w_eco4574, w_eco4575, w_eco4576, w_eco4577, w_eco4578, w_eco4579, w_eco4580, w_eco4581, w_eco4582, w_eco4583, w_eco4584, w_eco4585, w_eco4586, w_eco4587, w_eco4588, w_eco4589, w_eco4590, w_eco4591, w_eco4592, w_eco4593, w_eco4594, w_eco4595, w_eco4596, w_eco4597, w_eco4598, w_eco4599, w_eco4600, w_eco4601, w_eco4602, w_eco4603, w_eco4604, w_eco4605, w_eco4606, w_eco4607, w_eco4608, w_eco4609, w_eco4610, w_eco4611, w_eco4612, w_eco4613, w_eco4614, w_eco4615, w_eco4616, w_eco4617, w_eco4618, w_eco4619, w_eco4620, w_eco4621, w_eco4622, w_eco4623, w_eco4624, w_eco4625, w_eco4626, w_eco4627, w_eco4628, w_eco4629, w_eco4630, w_eco4631, w_eco4632, w_eco4633, w_eco4634, w_eco4635, w_eco4636, w_eco4637, w_eco4638, w_eco4639, w_eco4640, w_eco4641, w_eco4642, w_eco4643, w_eco4644, w_eco4645, w_eco4646, w_eco4647, w_eco4648, w_eco4649, w_eco4650, w_eco4651, w_eco4652, w_eco4653, w_eco4654, w_eco4655, w_eco4656, w_eco4657, w_eco4658, w_eco4659, w_eco4660, w_eco4661, w_eco4662, w_eco4663, w_eco4664, w_eco4665, w_eco4666, w_eco4667, w_eco4668, w_eco4669, w_eco4670, w_eco4671, w_eco4672, w_eco4673, w_eco4674, w_eco4675, w_eco4676, w_eco4677, w_eco4678, w_eco4679, w_eco4680, w_eco4681, w_eco4682, w_eco4683, w_eco4684, w_eco4685, w_eco4686, w_eco4687, w_eco4688, w_eco4689, w_eco4690, w_eco4691, w_eco4692, w_eco4693, w_eco4694, w_eco4695, w_eco4696, w_eco4697, w_eco4698, w_eco4699, w_eco4700, w_eco4701, w_eco4702, w_eco4703, w_eco4704, w_eco4705, w_eco4706, w_eco4707, w_eco4708, w_eco4709, w_eco4710, w_eco4711, w_eco4712, w_eco4713, w_eco4714, w_eco4715, w_eco4716, w_eco4717, w_eco4718, w_eco4719, w_eco4720, w_eco4721, w_eco4722, w_eco4723, w_eco4724, w_eco4725, w_eco4726, w_eco4727, w_eco4728, w_eco4729, w_eco4730, w_eco4731, w_eco4732, w_eco4733, w_eco4734, w_eco4735, w_eco4736, w_eco4737, w_eco4738, w_eco4739, w_eco4740, w_eco4741, w_eco4742, w_eco4743, w_eco4744, w_eco4745, w_eco4746, w_eco4747, w_eco4748, w_eco4749, w_eco4750, w_eco4751, w_eco4752, w_eco4753, w_eco4754, w_eco4755, w_eco4756, w_eco4757, w_eco4758, w_eco4759, w_eco4760, w_eco4761, w_eco4762, w_eco4763, w_eco4764, w_eco4765, w_eco4766, w_eco4767, w_eco4768, w_eco4769, w_eco4770, w_eco4771, w_eco4772, w_eco4773, w_eco4774, w_eco4775, w_eco4776, w_eco4777, w_eco4778, w_eco4779, w_eco4780, w_eco4781, w_eco4782, w_eco4783, w_eco4784, w_eco4785, w_eco4786, w_eco4787, w_eco4788, w_eco4789, w_eco4790, w_eco4791, w_eco4792, w_eco4793, w_eco4794, w_eco4795, w_eco4796, w_eco4797, w_eco4798, w_eco4799, w_eco4800, w_eco4801, w_eco4802, w_eco4803, w_eco4804, w_eco4805, w_eco4806, w_eco4807, w_eco4808, w_eco4809, w_eco4810, w_eco4811, w_eco4812, w_eco4813, w_eco4814, w_eco4815, w_eco4816, w_eco4817, w_eco4818, w_eco4819, w_eco4820, w_eco4821, w_eco4822, w_eco4823, w_eco4824, w_eco4825, w_eco4826, w_eco4827, w_eco4828, w_eco4829, w_eco4830, w_eco4831, w_eco4832, w_eco4833, w_eco4834, w_eco4835, w_eco4836, w_eco4837, w_eco4838, w_eco4839, w_eco4840, w_eco4841, w_eco4842, w_eco4843, w_eco4844, w_eco4845, w_eco4846, w_eco4847, w_eco4848, w_eco4849, w_eco4850, w_eco4851, w_eco4852, w_eco4853, w_eco4854, w_eco4855, w_eco4856, w_eco4857, w_eco4858, w_eco4859, w_eco4860, w_eco4861, w_eco4862, w_eco4863, w_eco4864, w_eco4865, w_eco4866, w_eco4867, w_eco4868, w_eco4869, w_eco4870, w_eco4871, w_eco4872, w_eco4873, w_eco4874, w_eco4875, w_eco4876, w_eco4877, w_eco4878, w_eco4879, w_eco4880, w_eco4881, w_eco4882, w_eco4883, w_eco4884, w_eco4885, w_eco4886, w_eco4887, w_eco4888, w_eco4889, w_eco4890, w_eco4891, w_eco4892, w_eco4893, w_eco4894, w_eco4895, w_eco4896, w_eco4897, w_eco4898, w_eco4899, w_eco4900, w_eco4901, w_eco4902, w_eco4903, w_eco4904, w_eco4905, w_eco4906, w_eco4907, w_eco4908, w_eco4909, w_eco4910, w_eco4911, w_eco4912, w_eco4913, w_eco4914, w_eco4915, w_eco4916, w_eco4917, w_eco4918, w_eco4919, w_eco4920, w_eco4921, w_eco4922, w_eco4923, w_eco4924, w_eco4925, w_eco4926, w_eco4927, w_eco4928, w_eco4929, w_eco4930, w_eco4931, w_eco4932, w_eco4933, w_eco4934, w_eco4935, w_eco4936, w_eco4937, w_eco4938, w_eco4939, w_eco4940, w_eco4941, w_eco4942, w_eco4943, w_eco4944, w_eco4945, w_eco4946, w_eco4947, w_eco4948, w_eco4949, w_eco4950, w_eco4951, w_eco4952, w_eco4953, w_eco4954, w_eco4955, w_eco4956, w_eco4957, w_eco4958, w_eco4959, w_eco4960, w_eco4961, w_eco4962, w_eco4963, w_eco4964, w_eco4965, w_eco4966, w_eco4967, w_eco4968, w_eco4969, w_eco4970, w_eco4971, w_eco4972, w_eco4973, w_eco4974, w_eco4975, w_eco4976, w_eco4977, w_eco4978, w_eco4979, w_eco4980, w_eco4981, w_eco4982, w_eco4983, w_eco4984, w_eco4985, w_eco4986, w_eco4987, w_eco4988, w_eco4989, w_eco4990, w_eco4991, w_eco4992, w_eco4993, w_eco4994, w_eco4995, w_eco4996, w_eco4997, w_eco4998, w_eco4999, w_eco5000, w_eco5001, w_eco5002, w_eco5003, w_eco5004, w_eco5005, w_eco5006, w_eco5007, w_eco5008, w_eco5009, w_eco5010, w_eco5011, w_eco5012, w_eco5013, w_eco5014, w_eco5015, w_eco5016, w_eco5017, w_eco5018, w_eco5019, w_eco5020, w_eco5021, w_eco5022, w_eco5023, w_eco5024, w_eco5025, w_eco5026, w_eco5027, w_eco5028, w_eco5029, w_eco5030, w_eco5031, w_eco5032, w_eco5033, w_eco5034, w_eco5035, w_eco5036, w_eco5037, w_eco5038, w_eco5039, w_eco5040, w_eco5041, w_eco5042, w_eco5043, w_eco5044, w_eco5045, w_eco5046, w_eco5047, w_eco5048, w_eco5049, w_eco5050, w_eco5051, w_eco5052, w_eco5053, w_eco5054, w_eco5055, w_eco5056, w_eco5057, w_eco5058, w_eco5059, w_eco5060, w_eco5061, w_eco5062, w_eco5063, w_eco5064, w_eco5065, w_eco5066, w_eco5067, w_eco5068, w_eco5069, w_eco5070, w_eco5071, w_eco5072, w_eco5073, w_eco5074, w_eco5075, w_eco5076, w_eco5077, w_eco5078, w_eco5079, w_eco5080, w_eco5081, w_eco5082, w_eco5083, w_eco5084, w_eco5085, w_eco5086, w_eco5087, w_eco5088, w_eco5089, w_eco5090, w_eco5091, w_eco5092, w_eco5093, w_eco5094, w_eco5095, w_eco5096, w_eco5097, w_eco5098, w_eco5099, w_eco5100, w_eco5101, w_eco5102, w_eco5103, w_eco5104, w_eco5105, w_eco5106, w_eco5107, w_eco5108, w_eco5109, w_eco5110, w_eco5111, w_eco5112, w_eco5113, w_eco5114, w_eco5115, w_eco5116, w_eco5117, w_eco5118, w_eco5119, w_eco5120, w_eco5121, w_eco5122, w_eco5123, w_eco5124, w_eco5125, w_eco5126, w_eco5127, w_eco5128, w_eco5129, w_eco5130, w_eco5131, w_eco5132, w_eco5133, w_eco5134, w_eco5135, w_eco5136, w_eco5137, w_eco5138, w_eco5139, w_eco5140, w_eco5141, w_eco5142, w_eco5143, w_eco5144, w_eco5145, w_eco5146, w_eco5147, w_eco5148, w_eco5149, w_eco5150, w_eco5151, w_eco5152, w_eco5153, w_eco5154, w_eco5155, w_eco5156, w_eco5157, w_eco5158, w_eco5159, w_eco5160, w_eco5161, w_eco5162, w_eco5163, w_eco5164, w_eco5165, w_eco5166, w_eco5167, w_eco5168, w_eco5169, w_eco5170, w_eco5171, w_eco5172, w_eco5173, w_eco5174, w_eco5175, w_eco5176, w_eco5177, w_eco5178, w_eco5179, w_eco5180, w_eco5181, w_eco5182, w_eco5183, w_eco5184, w_eco5185, w_eco5186, w_eco5187, w_eco5188, w_eco5189, w_eco5190, w_eco5191, w_eco5192, w_eco5193, w_eco5194, w_eco5195, w_eco5196, w_eco5197, w_eco5198, w_eco5199, w_eco5200, w_eco5201, w_eco5202, w_eco5203, w_eco5204, w_eco5205, w_eco5206, w_eco5207, w_eco5208, w_eco5209, w_eco5210, w_eco5211, w_eco5212, w_eco5213, w_eco5214, w_eco5215, w_eco5216, w_eco5217, w_eco5218, w_eco5219, w_eco5220, w_eco5221, w_eco5222, w_eco5223, w_eco5224, w_eco5225, w_eco5226, w_eco5227, w_eco5228, w_eco5229, w_eco5230, w_eco5231, w_eco5232, w_eco5233, w_eco5234, w_eco5235, w_eco5236, w_eco5237, w_eco5238, w_eco5239, w_eco5240, w_eco5241, w_eco5242, w_eco5243, w_eco5244, w_eco5245, w_eco5246, w_eco5247, w_eco5248, w_eco5249, w_eco5250, w_eco5251, w_eco5252, w_eco5253, w_eco5254, w_eco5255, w_eco5256, w_eco5257, w_eco5258, w_eco5259, w_eco5260, w_eco5261, w_eco5262, w_eco5263, w_eco5264, w_eco5265, w_eco5266, w_eco5267, w_eco5268, w_eco5269, w_eco5270, w_eco5271, w_eco5272, w_eco5273, w_eco5274, w_eco5275, w_eco5276, w_eco5277, w_eco5278, w_eco5279, w_eco5280, w_eco5281, w_eco5282, w_eco5283, w_eco5284, w_eco5285, w_eco5286, w_eco5287, w_eco5288, w_eco5289, w_eco5290, w_eco5291, w_eco5292, w_eco5293, w_eco5294, w_eco5295, w_eco5296, w_eco5297, w_eco5298, w_eco5299, w_eco5300, w_eco5301, w_eco5302, w_eco5303, w_eco5304, w_eco5305, w_eco5306, w_eco5307, w_eco5308, w_eco5309, w_eco5310, w_eco5311, w_eco5312, w_eco5313, w_eco5314, w_eco5315, w_eco5316, w_eco5317, w_eco5318, w_eco5319, w_eco5320, w_eco5321, w_eco5322, w_eco5323, w_eco5324, w_eco5325, w_eco5326, w_eco5327, w_eco5328, w_eco5329, w_eco5330, w_eco5331, w_eco5332, w_eco5333, w_eco5334, w_eco5335, w_eco5336, w_eco5337, w_eco5338, w_eco5339, w_eco5340, w_eco5341, w_eco5342, w_eco5343, w_eco5344, w_eco5345, w_eco5346, w_eco5347, w_eco5348, w_eco5349, w_eco5350, w_eco5351, w_eco5352, w_eco5353, w_eco5354, w_eco5355, w_eco5356, w_eco5357, w_eco5358, w_eco5359, w_eco5360, w_eco5361, w_eco5362, w_eco5363, w_eco5364, w_eco5365, w_eco5366, w_eco5367, w_eco5368, w_eco5369, w_eco5370, w_eco5371, w_eco5372, w_eco5373, w_eco5374, w_eco5375, w_eco5376, w_eco5377, w_eco5378, w_eco5379, w_eco5380, w_eco5381, w_eco5382, w_eco5383, w_eco5384, w_eco5385, w_eco5386, w_eco5387, w_eco5388, w_eco5389, w_eco5390, w_eco5391, w_eco5392, w_eco5393, w_eco5394, w_eco5395, w_eco5396, w_eco5397, w_eco5398, w_eco5399, w_eco5400, w_eco5401, w_eco5402, w_eco5403, w_eco5404, w_eco5405, w_eco5406, w_eco5407, w_eco5408, w_eco5409, w_eco5410, w_eco5411, w_eco5412, w_eco5413, w_eco5414, w_eco5415, w_eco5416, w_eco5417, w_eco5418, w_eco5419, w_eco5420, w_eco5421, w_eco5422, w_eco5423, w_eco5424, w_eco5425, w_eco5426, w_eco5427, w_eco5428, w_eco5429, w_eco5430, w_eco5431, w_eco5432, w_eco5433, w_eco5434, w_eco5435, w_eco5436, w_eco5437, w_eco5438, w_eco5439, w_eco5440, w_eco5441, w_eco5442, w_eco5443, w_eco5444, w_eco5445, w_eco5446, w_eco5447, w_eco5448, w_eco5449, w_eco5450, w_eco5451, w_eco5452, w_eco5453, w_eco5454, w_eco5455, w_eco5456, w_eco5457, w_eco5458, w_eco5459, w_eco5460, w_eco5461, w_eco5462, w_eco5463, w_eco5464, w_eco5465, w_eco5466, w_eco5467, w_eco5468, w_eco5469, w_eco5470, w_eco5471, w_eco5472, w_eco5473, w_eco5474, w_eco5475, w_eco5476, w_eco5477, w_eco5478, w_eco5479, w_eco5480, w_eco5481, w_eco5482, w_eco5483, w_eco5484, w_eco5485, w_eco5486, w_eco5487, w_eco5488, w_eco5489, w_eco5490, w_eco5491, w_eco5492, w_eco5493, w_eco5494, w_eco5495, w_eco5496, w_eco5497, w_eco5498, w_eco5499, w_eco5500, w_eco5501, w_eco5502, w_eco5503, w_eco5504, w_eco5505, w_eco5506, w_eco5507, w_eco5508, w_eco5509, w_eco5510, w_eco5511, w_eco5512, w_eco5513, w_eco5514, w_eco5515, w_eco5516, w_eco5517, w_eco5518, w_eco5519, w_eco5520, w_eco5521, w_eco5522, w_eco5523, w_eco5524, w_eco5525, w_eco5526, w_eco5527, w_eco5528, w_eco5529, w_eco5530, w_eco5531, w_eco5532, w_eco5533, w_eco5534, w_eco5535, w_eco5536, w_eco5537, w_eco5538, w_eco5539, w_eco5540, w_eco5541, w_eco5542, w_eco5543, w_eco5544, w_eco5545, w_eco5546, w_eco5547, w_eco5548, w_eco5549, w_eco5550, w_eco5551, w_eco5552, w_eco5553, w_eco5554, w_eco5555, w_eco5556, w_eco5557, w_eco5558, w_eco5559, w_eco5560, w_eco5561, w_eco5562, w_eco5563, w_eco5564, w_eco5565, w_eco5566, w_eco5567, w_eco5568, w_eco5569, w_eco5570, w_eco5571, w_eco5572, w_eco5573, w_eco5574, w_eco5575, w_eco5576, w_eco5577, w_eco5578, w_eco5579, w_eco5580, w_eco5581, w_eco5582, w_eco5583, w_eco5584, w_eco5585, w_eco5586, w_eco5587, w_eco5588, w_eco5589, w_eco5590, w_eco5591, w_eco5592, w_eco5593, w_eco5594, w_eco5595, w_eco5596, w_eco5597, w_eco5598, w_eco5599, w_eco5600, w_eco5601, w_eco5602, w_eco5603, w_eco5604, w_eco5605, w_eco5606, w_eco5607, w_eco5608, w_eco5609, w_eco5610, w_eco5611, w_eco5612, w_eco5613, w_eco5614, w_eco5615, w_eco5616, w_eco5617, w_eco5618, w_eco5619, w_eco5620, w_eco5621, w_eco5622, w_eco5623, w_eco5624, w_eco5625, w_eco5626, w_eco5627, w_eco5628, w_eco5629, w_eco5630, w_eco5631, w_eco5632, w_eco5633, w_eco5634, w_eco5635, w_eco5636, w_eco5637, w_eco5638, w_eco5639, w_eco5640, w_eco5641, w_eco5642, w_eco5643, w_eco5644, w_eco5645, w_eco5646, w_eco5647, w_eco5648, w_eco5649, w_eco5650, w_eco5651, w_eco5652, w_eco5653, w_eco5654, w_eco5655, w_eco5656, w_eco5657, w_eco5658, w_eco5659, w_eco5660, w_eco5661, w_eco5662, w_eco5663, w_eco5664, w_eco5665, w_eco5666, w_eco5667, w_eco5668, w_eco5669, w_eco5670, w_eco5671, w_eco5672, w_eco5673, w_eco5674, w_eco5675, w_eco5676, w_eco5677, w_eco5678, w_eco5679, w_eco5680, w_eco5681, w_eco5682, w_eco5683, w_eco5684, w_eco5685, w_eco5686, w_eco5687, w_eco5688, w_eco5689, w_eco5690, w_eco5691, w_eco5692, w_eco5693, w_eco5694, w_eco5695, w_eco5696, w_eco5697, w_eco5698, w_eco5699, w_eco5700, w_eco5701, w_eco5702, w_eco5703, w_eco5704, w_eco5705, w_eco5706, w_eco5707, w_eco5708, w_eco5709, w_eco5710, w_eco5711, w_eco5712, w_eco5713, w_eco5714, w_eco5715, w_eco5716, w_eco5717, w_eco5718, w_eco5719, w_eco5720, w_eco5721, w_eco5722, w_eco5723, w_eco5724, w_eco5725, w_eco5726, w_eco5727, w_eco5728, w_eco5729, w_eco5730, w_eco5731, w_eco5732, w_eco5733, w_eco5734, w_eco5735, w_eco5736, w_eco5737, w_eco5738, w_eco5739, w_eco5740, w_eco5741, w_eco5742, w_eco5743, w_eco5744, w_eco5745, w_eco5746, w_eco5747, w_eco5748, w_eco5749, w_eco5750, w_eco5751, w_eco5752, w_eco5753, w_eco5754, w_eco5755, w_eco5756, w_eco5757, w_eco5758, w_eco5759, w_eco5760, w_eco5761, w_eco5762, w_eco5763, w_eco5764, w_eco5765, w_eco5766, w_eco5767, w_eco5768, w_eco5769, w_eco5770, w_eco5771, w_eco5772, w_eco5773, w_eco5774, w_eco5775, w_eco5776, w_eco5777, w_eco5778, w_eco5779, w_eco5780, w_eco5781, w_eco5782, w_eco5783, w_eco5784, w_eco5785, w_eco5786, w_eco5787, w_eco5788, w_eco5789, w_eco5790, w_eco5791, w_eco5792, w_eco5793, w_eco5794, w_eco5795, w_eco5796, w_eco5797, w_eco5798, w_eco5799, w_eco5800, w_eco5801, w_eco5802, w_eco5803, w_eco5804, w_eco5805, w_eco5806, w_eco5807, w_eco5808, w_eco5809, w_eco5810, w_eco5811, w_eco5812, w_eco5813, w_eco5814, w_eco5815, w_eco5816, w_eco5817, w_eco5818, w_eco5819, w_eco5820, w_eco5821, w_eco5822, w_eco5823, w_eco5824, w_eco5825, w_eco5826, w_eco5827, w_eco5828, w_eco5829, w_eco5830, w_eco5831, w_eco5832, w_eco5833, w_eco5834, w_eco5835, w_eco5836, w_eco5837, w_eco5838, w_eco5839, w_eco5840, w_eco5841, w_eco5842, w_eco5843, w_eco5844, w_eco5845, w_eco5846, w_eco5847, w_eco5848, w_eco5849, w_eco5850, w_eco5851, w_eco5852, w_eco5853, w_eco5854, w_eco5855, w_eco5856, w_eco5857, w_eco5858, w_eco5859, w_eco5860, w_eco5861, w_eco5862, w_eco5863, w_eco5864, w_eco5865, w_eco5866, w_eco5867, w_eco5868, w_eco5869, w_eco5870, w_eco5871, w_eco5872, w_eco5873, w_eco5874, w_eco5875, w_eco5876, w_eco5877, w_eco5878, w_eco5879, w_eco5880, w_eco5881, w_eco5882, w_eco5883, w_eco5884, w_eco5885, w_eco5886, w_eco5887, w_eco5888, w_eco5889, w_eco5890, w_eco5891, w_eco5892, w_eco5893, w_eco5894, w_eco5895, w_eco5896, w_eco5897, w_eco5898, w_eco5899, w_eco5900, w_eco5901, w_eco5902, w_eco5903, w_eco5904, w_eco5905, w_eco5906, w_eco5907, w_eco5908, w_eco5909, w_eco5910, w_eco5911, w_eco5912, w_eco5913, w_eco5914, w_eco5915, w_eco5916, w_eco5917, w_eco5918, w_eco5919, w_eco5920, w_eco5921, w_eco5922, w_eco5923, w_eco5924, w_eco5925, w_eco5926, w_eco5927, w_eco5928, w_eco5929, w_eco5930, w_eco5931, w_eco5932, w_eco5933, w_eco5934, w_eco5935, w_eco5936, w_eco5937, w_eco5938, w_eco5939, w_eco5940, w_eco5941, w_eco5942, w_eco5943, w_eco5944, w_eco5945, w_eco5946, w_eco5947, w_eco5948, w_eco5949, w_eco5950, w_eco5951, w_eco5952, w_eco5953, w_eco5954, w_eco5955, w_eco5956, w_eco5957, w_eco5958, w_eco5959, w_eco5960, w_eco5961, w_eco5962, w_eco5963, w_eco5964, w_eco5965, w_eco5966, w_eco5967, w_eco5968, w_eco5969, w_eco5970, w_eco5971, w_eco5972, w_eco5973, w_eco5974, w_eco5975, w_eco5976, w_eco5977, w_eco5978, w_eco5979, w_eco5980, w_eco5981, w_eco5982, w_eco5983, w_eco5984, w_eco5985, w_eco5986, w_eco5987, w_eco5988, w_eco5989, w_eco5990, w_eco5991, w_eco5992, w_eco5993, w_eco5994, w_eco5995, w_eco5996, w_eco5997, w_eco5998, w_eco5999, w_eco6000, w_eco6001, w_eco6002, w_eco6003, w_eco6004, w_eco6005, w_eco6006, w_eco6007, w_eco6008, w_eco6009, w_eco6010, w_eco6011, w_eco6012, w_eco6013, w_eco6014, w_eco6015, w_eco6016, w_eco6017, w_eco6018, w_eco6019, w_eco6020, w_eco6021, w_eco6022, w_eco6023, w_eco6024, w_eco6025, w_eco6026, w_eco6027, w_eco6028, w_eco6029, w_eco6030, w_eco6031, w_eco6032, w_eco6033, w_eco6034, w_eco6035, w_eco6036, w_eco6037, w_eco6038, w_eco6039, w_eco6040, w_eco6041, w_eco6042, w_eco6043, w_eco6044, w_eco6045, w_eco6046, w_eco6047, w_eco6048, w_eco6049, w_eco6050, w_eco6051, w_eco6052, w_eco6053, w_eco6054, w_eco6055, w_eco6056, w_eco6057, w_eco6058, w_eco6059, w_eco6060, w_eco6061, w_eco6062, w_eco6063, w_eco6064, w_eco6065, w_eco6066, w_eco6067, w_eco6068, w_eco6069, w_eco6070, w_eco6071, w_eco6072, w_eco6073, w_eco6074, w_eco6075, w_eco6076, w_eco6077, w_eco6078, w_eco6079, w_eco6080, w_eco6081, w_eco6082, w_eco6083, w_eco6084, w_eco6085, w_eco6086, w_eco6087, w_eco6088, w_eco6089, w_eco6090, w_eco6091, w_eco6092, w_eco6093, w_eco6094, w_eco6095, w_eco6096, w_eco6097, w_eco6098, w_eco6099, w_eco6100, w_eco6101, w_eco6102, w_eco6103, w_eco6104, w_eco6105, w_eco6106, w_eco6107, w_eco6108, w_eco6109, w_eco6110, w_eco6111, w_eco6112, w_eco6113, w_eco6114, w_eco6115, w_eco6116, w_eco6117, w_eco6118, w_eco6119, w_eco6120, w_eco6121, w_eco6122, w_eco6123, w_eco6124, w_eco6125, w_eco6126, w_eco6127, w_eco6128, w_eco6129, w_eco6130, w_eco6131, w_eco6132, w_eco6133, w_eco6134, w_eco6135, w_eco6136, w_eco6137, w_eco6138, w_eco6139, w_eco6140, w_eco6141, w_eco6142, w_eco6143, w_eco6144, w_eco6145, w_eco6146, w_eco6147, w_eco6148, w_eco6149, w_eco6150, w_eco6151, w_eco6152, w_eco6153, w_eco6154, w_eco6155, w_eco6156, w_eco6157, w_eco6158, w_eco6159, w_eco6160, w_eco6161, w_eco6162, w_eco6163, w_eco6164, w_eco6165, w_eco6166, w_eco6167, w_eco6168, w_eco6169, w_eco6170, w_eco6171, w_eco6172, w_eco6173, w_eco6174, w_eco6175, w_eco6176, w_eco6177, w_eco6178, w_eco6179, w_eco6180, w_eco6181, w_eco6182, w_eco6183, w_eco6184, w_eco6185, w_eco6186, w_eco6187, w_eco6188, w_eco6189, w_eco6190, w_eco6191, w_eco6192, w_eco6193, w_eco6194, w_eco6195, w_eco6196, w_eco6197, w_eco6198, w_eco6199, w_eco6200, w_eco6201, w_eco6202, w_eco6203, w_eco6204, w_eco6205, w_eco6206, w_eco6207, w_eco6208, w_eco6209, w_eco6210, w_eco6211, w_eco6212, w_eco6213, w_eco6214, w_eco6215, w_eco6216, w_eco6217, w_eco6218, w_eco6219, w_eco6220, w_eco6221, w_eco6222, w_eco6223, w_eco6224, w_eco6225, w_eco6226, w_eco6227, w_eco6228, w_eco6229, w_eco6230, w_eco6231, w_eco6232, w_eco6233, w_eco6234, w_eco6235, w_eco6236, w_eco6237, w_eco6238, w_eco6239, w_eco6240, w_eco6241, w_eco6242, w_eco6243, w_eco6244, w_eco6245, w_eco6246, w_eco6247, w_eco6248, w_eco6249, w_eco6250, w_eco6251, w_eco6252, w_eco6253, w_eco6254, w_eco6255, w_eco6256, w_eco6257, w_eco6258, w_eco6259, w_eco6260, w_eco6261, w_eco6262, w_eco6263, w_eco6264, w_eco6265, w_eco6266, w_eco6267, w_eco6268, w_eco6269, w_eco6270, w_eco6271, w_eco6272, w_eco6273, w_eco6274, w_eco6275, w_eco6276, w_eco6277, w_eco6278, w_eco6279, w_eco6280, w_eco6281, w_eco6282, w_eco6283, w_eco6284, w_eco6285, w_eco6286, w_eco6287, w_eco6288, w_eco6289, w_eco6290, w_eco6291, w_eco6292, w_eco6293, w_eco6294, w_eco6295, w_eco6296, w_eco6297, w_eco6298, w_eco6299, w_eco6300, w_eco6301, w_eco6302, w_eco6303, w_eco6304, w_eco6305, w_eco6306, w_eco6307, w_eco6308, w_eco6309, w_eco6310, w_eco6311, w_eco6312, w_eco6313, w_eco6314, w_eco6315, w_eco6316, w_eco6317, w_eco6318, w_eco6319, w_eco6320, w_eco6321, w_eco6322, w_eco6323, w_eco6324, w_eco6325, w_eco6326, w_eco6327, w_eco6328, w_eco6329, w_eco6330, w_eco6331, w_eco6332, w_eco6333, w_eco6334, w_eco6335, w_eco6336, w_eco6337, w_eco6338, w_eco6339, w_eco6340, w_eco6341, w_eco6342, w_eco6343, w_eco6344, w_eco6345, w_eco6346, w_eco6347, w_eco6348, w_eco6349, w_eco6350, w_eco6351, w_eco6352, w_eco6353, w_eco6354, w_eco6355, w_eco6356, w_eco6357, w_eco6358, w_eco6359, w_eco6360, w_eco6361, w_eco6362, w_eco6363, w_eco6364, w_eco6365, w_eco6366, w_eco6367, w_eco6368, w_eco6369, w_eco6370, w_eco6371, w_eco6372, w_eco6373, w_eco6374, w_eco6375, w_eco6376, w_eco6377, w_eco6378, w_eco6379, w_eco6380, w_eco6381, w_eco6382, w_eco6383, w_eco6384, w_eco6385, w_eco6386, w_eco6387, w_eco6388, w_eco6389, w_eco6390, w_eco6391, w_eco6392, w_eco6393, w_eco6394, w_eco6395, w_eco6396, w_eco6397, w_eco6398, w_eco6399, w_eco6400, w_eco6401, w_eco6402, w_eco6403, w_eco6404, w_eco6405, w_eco6406, w_eco6407, w_eco6408, w_eco6409, w_eco6410, w_eco6411, w_eco6412, w_eco6413, w_eco6414, w_eco6415, w_eco6416, w_eco6417, w_eco6418, w_eco6419, w_eco6420, w_eco6421, w_eco6422, w_eco6423, w_eco6424, w_eco6425, w_eco6426, w_eco6427, w_eco6428, w_eco6429, w_eco6430, w_eco6431, w_eco6432, w_eco6433, w_eco6434, w_eco6435, w_eco6436, w_eco6437, w_eco6438, w_eco6439, w_eco6440, w_eco6441, w_eco6442, w_eco6443, w_eco6444, w_eco6445, w_eco6446, w_eco6447, w_eco6448, w_eco6449, w_eco6450, w_eco6451, w_eco6452, w_eco6453, w_eco6454, w_eco6455, w_eco6456, w_eco6457, w_eco6458, w_eco6459, w_eco6460, w_eco6461, w_eco6462, w_eco6463, w_eco6464, w_eco6465, w_eco6466, w_eco6467, w_eco6468, w_eco6469, w_eco6470, w_eco6471, w_eco6472, w_eco6473, w_eco6474, w_eco6475, w_eco6476, w_eco6477, w_eco6478, w_eco6479, w_eco6480, w_eco6481, w_eco6482, w_eco6483, w_eco6484, w_eco6485, w_eco6486, w_eco6487, w_eco6488, w_eco6489, w_eco6490, w_eco6491, w_eco6492, w_eco6493, w_eco6494, w_eco6495, w_eco6496, w_eco6497, w_eco6498, w_eco6499, w_eco6500, w_eco6501, w_eco6502, w_eco6503, w_eco6504, w_eco6505, w_eco6506, w_eco6507, w_eco6508, w_eco6509, w_eco6510, w_eco6511, w_eco6512, w_eco6513, w_eco6514, w_eco6515, w_eco6516, w_eco6517, w_eco6518, w_eco6519, w_eco6520, w_eco6521, w_eco6522, w_eco6523, w_eco6524, w_eco6525, w_eco6526, w_eco6527, w_eco6528, w_eco6529, w_eco6530, w_eco6531, w_eco6532, w_eco6533, w_eco6534, w_eco6535, w_eco6536, w_eco6537, w_eco6538, w_eco6539, w_eco6540, w_eco6541, w_eco6542, w_eco6543, w_eco6544, w_eco6545, w_eco6546, w_eco6547, w_eco6548, w_eco6549, w_eco6550, w_eco6551, w_eco6552, w_eco6553, w_eco6554, w_eco6555, w_eco6556, w_eco6557, w_eco6558, w_eco6559, w_eco6560, w_eco6561, w_eco6562, w_eco6563, w_eco6564, w_eco6565, w_eco6566, w_eco6567, w_eco6568, w_eco6569, w_eco6570, w_eco6571, w_eco6572, w_eco6573, w_eco6574, w_eco6575, w_eco6576, w_eco6577, w_eco6578, w_eco6579, w_eco6580, w_eco6581, w_eco6582, w_eco6583, w_eco6584, w_eco6585, w_eco6586, w_eco6587, w_eco6588, w_eco6589, w_eco6590, w_eco6591, w_eco6592, w_eco6593, w_eco6594, w_eco6595, w_eco6596, w_eco6597, w_eco6598, w_eco6599, w_eco6600, w_eco6601, w_eco6602, w_eco6603, w_eco6604, w_eco6605, w_eco6606, w_eco6607, w_eco6608, w_eco6609, w_eco6610, w_eco6611, w_eco6612, w_eco6613, w_eco6614, w_eco6615, w_eco6616, w_eco6617, w_eco6618, w_eco6619, w_eco6620, w_eco6621, w_eco6622, w_eco6623, w_eco6624, w_eco6625, w_eco6626, w_eco6627, w_eco6628, w_eco6629, w_eco6630, w_eco6631, w_eco6632, w_eco6633, w_eco6634, w_eco6635, w_eco6636, w_eco6637, w_eco6638, w_eco6639, w_eco6640, w_eco6641, w_eco6642, w_eco6643, w_eco6644, w_eco6645, w_eco6646, w_eco6647, w_eco6648, w_eco6649, w_eco6650, w_eco6651, w_eco6652, w_eco6653, w_eco6654, w_eco6655, w_eco6656, w_eco6657, w_eco6658, w_eco6659, w_eco6660, w_eco6661, w_eco6662, w_eco6663, w_eco6664, w_eco6665, w_eco6666, w_eco6667, w_eco6668, w_eco6669, w_eco6670, w_eco6671, w_eco6672, w_eco6673, w_eco6674, w_eco6675, w_eco6676, w_eco6677, w_eco6678, w_eco6679, w_eco6680, w_eco6681, w_eco6682, w_eco6683, w_eco6684, w_eco6685, w_eco6686, w_eco6687, w_eco6688, w_eco6689, w_eco6690, w_eco6691, w_eco6692, w_eco6693, w_eco6694, w_eco6695, w_eco6696, w_eco6697, w_eco6698, w_eco6699, w_eco6700, w_eco6701, w_eco6702, w_eco6703, w_eco6704, w_eco6705, w_eco6706, w_eco6707, w_eco6708, w_eco6709, w_eco6710, w_eco6711, w_eco6712, w_eco6713, w_eco6714, w_eco6715, w_eco6716, w_eco6717, w_eco6718, w_eco6719, w_eco6720, w_eco6721, w_eco6722, w_eco6723, w_eco6724, w_eco6725, w_eco6726, w_eco6727, w_eco6728, w_eco6729, w_eco6730, w_eco6731, w_eco6732, w_eco6733, w_eco6734, w_eco6735, w_eco6736, w_eco6737, w_eco6738, w_eco6739, w_eco6740, w_eco6741, w_eco6742, w_eco6743, w_eco6744, w_eco6745, w_eco6746, w_eco6747, w_eco6748, w_eco6749, w_eco6750, w_eco6751, w_eco6752, w_eco6753, w_eco6754, w_eco6755, w_eco6756, w_eco6757, w_eco6758, w_eco6759, w_eco6760, w_eco6761, w_eco6762, w_eco6763, w_eco6764, w_eco6765, w_eco6766, w_eco6767, w_eco6768, w_eco6769, w_eco6770, w_eco6771, w_eco6772, w_eco6773, w_eco6774, w_eco6775, w_eco6776, w_eco6777, w_eco6778, w_eco6779, w_eco6780, w_eco6781, w_eco6782, w_eco6783, w_eco6784, w_eco6785, w_eco6786, w_eco6787, w_eco6788, w_eco6789, w_eco6790, w_eco6791, w_eco6792, w_eco6793, w_eco6794, w_eco6795, w_eco6796, w_eco6797, w_eco6798, w_eco6799, w_eco6800, w_eco6801, w_eco6802, w_eco6803, w_eco6804, w_eco6805, w_eco6806, w_eco6807, w_eco6808, w_eco6809, w_eco6810, w_eco6811, w_eco6812, w_eco6813, w_eco6814, w_eco6815, w_eco6816, w_eco6817, w_eco6818, w_eco6819, w_eco6820, w_eco6821, w_eco6822, w_eco6823, w_eco6824, w_eco6825, w_eco6826, w_eco6827, w_eco6828, w_eco6829, w_eco6830, w_eco6831, w_eco6832, w_eco6833, w_eco6834, w_eco6835, w_eco6836, w_eco6837, w_eco6838, w_eco6839, w_eco6840, w_eco6841, w_eco6842, w_eco6843, w_eco6844, w_eco6845, w_eco6846, w_eco6847, w_eco6848, w_eco6849, w_eco6850, w_eco6851, w_eco6852, w_eco6853, w_eco6854, w_eco6855, w_eco6856, w_eco6857, w_eco6858, w_eco6859, w_eco6860, w_eco6861, w_eco6862, w_eco6863, w_eco6864, w_eco6865, w_eco6866, w_eco6867, w_eco6868, w_eco6869, w_eco6870, w_eco6871, w_eco6872, w_eco6873, w_eco6874, w_eco6875, w_eco6876, w_eco6877, w_eco6878, w_eco6879, w_eco6880, w_eco6881, w_eco6882, w_eco6883, w_eco6884, w_eco6885, w_eco6886, w_eco6887, w_eco6888, w_eco6889, w_eco6890, w_eco6891, w_eco6892, w_eco6893, w_eco6894, w_eco6895, w_eco6896, w_eco6897, w_eco6898, w_eco6899, w_eco6900, w_eco6901, w_eco6902, w_eco6903, w_eco6904, w_eco6905, w_eco6906, w_eco6907, w_eco6908, w_eco6909, w_eco6910, w_eco6911, w_eco6912, w_eco6913, w_eco6914, w_eco6915, w_eco6916, w_eco6917, w_eco6918, w_eco6919, w_eco6920, w_eco6921, w_eco6922, w_eco6923, w_eco6924, w_eco6925, w_eco6926, w_eco6927, w_eco6928, w_eco6929, w_eco6930, w_eco6931, w_eco6932, w_eco6933, w_eco6934, w_eco6935, w_eco6936, w_eco6937, w_eco6938, w_eco6939, w_eco6940, w_eco6941, w_eco6942, w_eco6943, w_eco6944, w_eco6945, w_eco6946, w_eco6947, w_eco6948, w_eco6949, w_eco6950, w_eco6951, w_eco6952, w_eco6953, w_eco6954, w_eco6955, w_eco6956, w_eco6957, w_eco6958, w_eco6959, w_eco6960, w_eco6961, w_eco6962, w_eco6963, w_eco6964, w_eco6965, w_eco6966, w_eco6967, w_eco6968, w_eco6969, w_eco6970, w_eco6971, w_eco6972, w_eco6973, w_eco6974, w_eco6975, w_eco6976, w_eco6977, w_eco6978, w_eco6979, w_eco6980, w_eco6981, w_eco6982, w_eco6983, w_eco6984, w_eco6985, w_eco6986, w_eco6987, w_eco6988, w_eco6989, w_eco6990, w_eco6991, w_eco6992, w_eco6993, w_eco6994, w_eco6995, w_eco6996, w_eco6997, w_eco6998, w_eco6999, w_eco7000, w_eco7001, w_eco7002, w_eco7003, w_eco7004, w_eco7005, w_eco7006, w_eco7007, w_eco7008, w_eco7009, w_eco7010, w_eco7011, w_eco7012, w_eco7013, w_eco7014, w_eco7015, w_eco7016, w_eco7017, w_eco7018, w_eco7019, w_eco7020, w_eco7021, w_eco7022, w_eco7023, w_eco7024, w_eco7025, w_eco7026, w_eco7027, w_eco7028, w_eco7029, w_eco7030, w_eco7031, w_eco7032, w_eco7033, w_eco7034, w_eco7035, w_eco7036, w_eco7037, w_eco7038, w_eco7039, w_eco7040, w_eco7041, w_eco7042, w_eco7043, w_eco7044, w_eco7045, w_eco7046, w_eco7047, w_eco7048, w_eco7049, w_eco7050, w_eco7051, w_eco7052, w_eco7053, w_eco7054, w_eco7055, w_eco7056, w_eco7057, w_eco7058, w_eco7059, w_eco7060, w_eco7061, w_eco7062, w_eco7063, w_eco7064, w_eco7065, w_eco7066, w_eco7067, w_eco7068, w_eco7069, w_eco7070, w_eco7071, w_eco7072, w_eco7073, w_eco7074, w_eco7075, w_eco7076, w_eco7077, w_eco7078, w_eco7079, w_eco7080, w_eco7081, w_eco7082, w_eco7083, w_eco7084, w_eco7085, w_eco7086, w_eco7087, w_eco7088, w_eco7089, w_eco7090, w_eco7091, w_eco7092, w_eco7093, w_eco7094, w_eco7095, w_eco7096, w_eco7097, w_eco7098, w_eco7099, w_eco7100, w_eco7101, w_eco7102, w_eco7103, w_eco7104, w_eco7105, w_eco7106, w_eco7107, w_eco7108, w_eco7109, w_eco7110, w_eco7111, w_eco7112, w_eco7113, w_eco7114, w_eco7115, w_eco7116, w_eco7117, w_eco7118, w_eco7119, w_eco7120, w_eco7121, w_eco7122, w_eco7123, w_eco7124, w_eco7125, w_eco7126, w_eco7127, w_eco7128, w_eco7129, w_eco7130, w_eco7131, w_eco7132, w_eco7133, w_eco7134, w_eco7135, w_eco7136, w_eco7137, w_eco7138, w_eco7139, w_eco7140, w_eco7141, w_eco7142, w_eco7143, w_eco7144, w_eco7145, w_eco7146, w_eco7147, w_eco7148, w_eco7149, w_eco7150, w_eco7151, w_eco7152, w_eco7153, w_eco7154, w_eco7155, w_eco7156, w_eco7157, w_eco7158, w_eco7159, w_eco7160, w_eco7161, w_eco7162, w_eco7163, w_eco7164, w_eco7165, w_eco7166, w_eco7167, w_eco7168, w_eco7169, w_eco7170, w_eco7171, w_eco7172, w_eco7173, w_eco7174, w_eco7175, w_eco7176, w_eco7177, w_eco7178, w_eco7179, w_eco7180, w_eco7181, w_eco7182, w_eco7183, w_eco7184, w_eco7185, w_eco7186, w_eco7187, w_eco7188, w_eco7189, w_eco7190, w_eco7191, w_eco7192, w_eco7193, w_eco7194, w_eco7195, w_eco7196, w_eco7197, w_eco7198, w_eco7199, w_eco7200, w_eco7201, w_eco7202, w_eco7203, w_eco7204, w_eco7205, w_eco7206, w_eco7207, w_eco7208, w_eco7209, w_eco7210, w_eco7211, w_eco7212, w_eco7213, w_eco7214, w_eco7215, w_eco7216, w_eco7217, w_eco7218, w_eco7219, w_eco7220, w_eco7221, w_eco7222, w_eco7223, w_eco7224, w_eco7225, w_eco7226, w_eco7227, w_eco7228, w_eco7229, w_eco7230, w_eco7231, w_eco7232, w_eco7233, w_eco7234, w_eco7235, w_eco7236, w_eco7237, w_eco7238, w_eco7239, w_eco7240, w_eco7241, w_eco7242, w_eco7243, w_eco7244, w_eco7245, w_eco7246, w_eco7247, w_eco7248, w_eco7249, w_eco7250, w_eco7251, w_eco7252, w_eco7253, w_eco7254, w_eco7255, w_eco7256, w_eco7257, w_eco7258, w_eco7259, w_eco7260, w_eco7261, w_eco7262, w_eco7263, w_eco7264, w_eco7265, w_eco7266, w_eco7267, w_eco7268, w_eco7269, w_eco7270, w_eco7271, w_eco7272, w_eco7273, w_eco7274, w_eco7275, w_eco7276, w_eco7277, w_eco7278, w_eco7279, w_eco7280, w_eco7281, w_eco7282, w_eco7283, w_eco7284, w_eco7285, w_eco7286, w_eco7287, w_eco7288, w_eco7289, w_eco7290, w_eco7291, w_eco7292, w_eco7293, w_eco7294, w_eco7295, w_eco7296, w_eco7297, w_eco7298, w_eco7299, w_eco7300, w_eco7301, w_eco7302, w_eco7303, w_eco7304, w_eco7305, w_eco7306, w_eco7307, w_eco7308, w_eco7309, w_eco7310, w_eco7311, w_eco7312, w_eco7313, w_eco7314, w_eco7315, w_eco7316, w_eco7317, w_eco7318, w_eco7319, w_eco7320, w_eco7321, w_eco7322, w_eco7323, w_eco7324, w_eco7325, w_eco7326, w_eco7327, w_eco7328, w_eco7329, w_eco7330, w_eco7331, w_eco7332, w_eco7333, w_eco7334, w_eco7335, w_eco7336, w_eco7337, w_eco7338, w_eco7339, w_eco7340, w_eco7341, w_eco7342, w_eco7343, w_eco7344, w_eco7345, w_eco7346, w_eco7347, w_eco7348, w_eco7349, w_eco7350, w_eco7351, w_eco7352, w_eco7353, w_eco7354, w_eco7355, w_eco7356, w_eco7357, w_eco7358, w_eco7359, w_eco7360, w_eco7361, w_eco7362, w_eco7363, w_eco7364, w_eco7365, w_eco7366, w_eco7367, w_eco7368, w_eco7369, w_eco7370, w_eco7371, w_eco7372, w_eco7373, w_eco7374, w_eco7375, w_eco7376, w_eco7377, w_eco7378, w_eco7379, w_eco7380, w_eco7381, w_eco7382, w_eco7383, w_eco7384, w_eco7385, w_eco7386, w_eco7387, w_eco7388, w_eco7389, w_eco7390, w_eco7391, w_eco7392, w_eco7393, w_eco7394, w_eco7395, w_eco7396, w_eco7397, w_eco7398, w_eco7399, w_eco7400, w_eco7401, w_eco7402, w_eco7403, w_eco7404, w_eco7405, w_eco7406, w_eco7407, w_eco7408, w_eco7409, w_eco7410, w_eco7411, w_eco7412, w_eco7413, w_eco7414, w_eco7415, w_eco7416, w_eco7417, w_eco7418, w_eco7419, w_eco7420, w_eco7421, w_eco7422, w_eco7423, w_eco7424, w_eco7425, w_eco7426, w_eco7427, w_eco7428, w_eco7429, w_eco7430, w_eco7431, w_eco7432, w_eco7433, w_eco7434, w_eco7435, w_eco7436, w_eco7437, w_eco7438, w_eco7439, w_eco7440, w_eco7441, w_eco7442, w_eco7443, w_eco7444, w_eco7445, w_eco7446, w_eco7447, w_eco7448, w_eco7449, w_eco7450, w_eco7451, w_eco7452, w_eco7453, w_eco7454, w_eco7455, w_eco7456, w_eco7457, w_eco7458, w_eco7459, w_eco7460, w_eco7461, w_eco7462, w_eco7463, w_eco7464, w_eco7465, w_eco7466, w_eco7467, w_eco7468, w_eco7469, w_eco7470, w_eco7471, w_eco7472, w_eco7473, w_eco7474, w_eco7475, w_eco7476, w_eco7477, w_eco7478, w_eco7479, w_eco7480, w_eco7481, w_eco7482, w_eco7483, w_eco7484, w_eco7485, w_eco7486, w_eco7487, w_eco7488, w_eco7489, w_eco7490, w_eco7491, w_eco7492, w_eco7493, w_eco7494, w_eco7495, w_eco7496, w_eco7497, w_eco7498, w_eco7499, w_eco7500, w_eco7501, w_eco7502, w_eco7503, w_eco7504, w_eco7505, w_eco7506, w_eco7507, w_eco7508, w_eco7509, w_eco7510, w_eco7511, w_eco7512, w_eco7513, w_eco7514, w_eco7515, w_eco7516, w_eco7517, w_eco7518, w_eco7519, w_eco7520, w_eco7521, w_eco7522, w_eco7523, w_eco7524, w_eco7525, w_eco7526, w_eco7527, w_eco7528, w_eco7529, w_eco7530, w_eco7531, w_eco7532, w_eco7533, w_eco7534, w_eco7535, w_eco7536, w_eco7537, w_eco7538, w_eco7539, w_eco7540, w_eco7541, w_eco7542, w_eco7543, w_eco7544, w_eco7545, w_eco7546, w_eco7547, w_eco7548, w_eco7549, w_eco7550, w_eco7551, w_eco7552, w_eco7553, w_eco7554, w_eco7555, w_eco7556, w_eco7557, w_eco7558, w_eco7559, w_eco7560, w_eco7561, w_eco7562, w_eco7563, w_eco7564, w_eco7565, w_eco7566, w_eco7567, w_eco7568, w_eco7569, w_eco7570, w_eco7571, w_eco7572, w_eco7573, w_eco7574, w_eco7575, w_eco7576, w_eco7577, w_eco7578, w_eco7579, w_eco7580, w_eco7581, w_eco7582, w_eco7583, w_eco7584, w_eco7585, w_eco7586, w_eco7587, w_eco7588, w_eco7589, w_eco7590, w_eco7591, w_eco7592, w_eco7593, w_eco7594, w_eco7595, w_eco7596, w_eco7597, w_eco7598, w_eco7599, w_eco7600, w_eco7601, w_eco7602, w_eco7603, w_eco7604, w_eco7605, w_eco7606, w_eco7607, w_eco7608, w_eco7609, w_eco7610, w_eco7611, w_eco7612, w_eco7613, w_eco7614, w_eco7615, w_eco7616, w_eco7617, w_eco7618, w_eco7619, w_eco7620, w_eco7621, w_eco7622, w_eco7623, w_eco7624, w_eco7625, w_eco7626, w_eco7627, w_eco7628, w_eco7629, w_eco7630, w_eco7631, w_eco7632, w_eco7633, w_eco7634, w_eco7635, w_eco7636, w_eco7637, w_eco7638, w_eco7639, w_eco7640, w_eco7641, w_eco7642, w_eco7643, w_eco7644, w_eco7645, w_eco7646, w_eco7647, w_eco7648, w_eco7649, w_eco7650, w_eco7651, w_eco7652, w_eco7653, w_eco7654, w_eco7655, w_eco7656, w_eco7657, w_eco7658, w_eco7659, w_eco7660, w_eco7661, w_eco7662, w_eco7663, w_eco7664, w_eco7665, w_eco7666, w_eco7667, w_eco7668, w_eco7669, w_eco7670, w_eco7671, w_eco7672, w_eco7673, w_eco7674, w_eco7675, w_eco7676, w_eco7677, w_eco7678, w_eco7679, w_eco7680, w_eco7681, w_eco7682, w_eco7683, w_eco7684, w_eco7685, w_eco7686, w_eco7687, w_eco7688, w_eco7689, w_eco7690, w_eco7691, w_eco7692, w_eco7693, w_eco7694, w_eco7695, w_eco7696, w_eco7697, w_eco7698, w_eco7699, w_eco7700, w_eco7701, w_eco7702, w_eco7703, w_eco7704, w_eco7705, w_eco7706, w_eco7707, w_eco7708, w_eco7709, w_eco7710, w_eco7711, w_eco7712, w_eco7713, w_eco7714, w_eco7715, w_eco7716, w_eco7717, w_eco7718, w_eco7719, w_eco7720, w_eco7721, w_eco7722, w_eco7723, w_eco7724, w_eco7725, w_eco7726, w_eco7727, w_eco7728, w_eco7729, w_eco7730, w_eco7731, w_eco7732, w_eco7733, w_eco7734, w_eco7735, w_eco7736, w_eco7737, w_eco7738, w_eco7739, w_eco7740, w_eco7741, w_eco7742, w_eco7743, w_eco7744, w_eco7745, w_eco7746, w_eco7747, w_eco7748, w_eco7749, w_eco7750, w_eco7751, w_eco7752, w_eco7753, w_eco7754, w_eco7755, w_eco7756, w_eco7757, w_eco7758, w_eco7759, w_eco7760, w_eco7761, w_eco7762, w_eco7763, w_eco7764, w_eco7765, w_eco7766, w_eco7767, w_eco7768, w_eco7769, w_eco7770, w_eco7771, w_eco7772, w_eco7773, w_eco7774, w_eco7775, w_eco7776, w_eco7777, w_eco7778, w_eco7779, w_eco7780, w_eco7781, w_eco7782, w_eco7783, w_eco7784, w_eco7785, w_eco7786, w_eco7787, w_eco7788, w_eco7789, w_eco7790, w_eco7791, w_eco7792, w_eco7793, w_eco7794, w_eco7795, w_eco7796, w_eco7797, w_eco7798, w_eco7799, w_eco7800, w_eco7801, w_eco7802, w_eco7803, w_eco7804, w_eco7805, w_eco7806, w_eco7807, w_eco7808, w_eco7809, w_eco7810, w_eco7811, w_eco7812, w_eco7813, w_eco7814, w_eco7815, w_eco7816, w_eco7817, w_eco7818, w_eco7819, w_eco7820, w_eco7821, w_eco7822, w_eco7823, w_eco7824, w_eco7825, w_eco7826, w_eco7827, w_eco7828, w_eco7829, w_eco7830, w_eco7831, w_eco7832, w_eco7833, w_eco7834, w_eco7835, w_eco7836, w_eco7837, w_eco7838, w_eco7839, w_eco7840, w_eco7841, w_eco7842, w_eco7843, w_eco7844, w_eco7845, w_eco7846, w_eco7847, w_eco7848, w_eco7849, w_eco7850, w_eco7851, w_eco7852, w_eco7853, w_eco7854, w_eco7855, w_eco7856, w_eco7857, w_eco7858, w_eco7859, w_eco7860, w_eco7861, w_eco7862, w_eco7863, w_eco7864, w_eco7865, w_eco7866, w_eco7867, w_eco7868, w_eco7869, w_eco7870, w_eco7871, w_eco7872, w_eco7873, w_eco7874, w_eco7875, w_eco7876, w_eco7877, w_eco7878, w_eco7879, w_eco7880, w_eco7881, w_eco7882, w_eco7883, w_eco7884, w_eco7885, w_eco7886, w_eco7887, w_eco7888, w_eco7889, w_eco7890, w_eco7891, w_eco7892, w_eco7893, w_eco7894, w_eco7895, w_eco7896, w_eco7897, w_eco7898, w_eco7899, w_eco7900, w_eco7901, w_eco7902, w_eco7903, w_eco7904, w_eco7905, w_eco7906, w_eco7907, w_eco7908, w_eco7909, w_eco7910, w_eco7911, w_eco7912, w_eco7913, w_eco7914, w_eco7915, w_eco7916, w_eco7917, w_eco7918, w_eco7919, w_eco7920, w_eco7921, w_eco7922, w_eco7923, w_eco7924, w_eco7925, w_eco7926, w_eco7927, w_eco7928, w_eco7929, w_eco7930, w_eco7931, w_eco7932, w_eco7933, w_eco7934, w_eco7935, w_eco7936, w_eco7937, w_eco7938, w_eco7939, w_eco7940, w_eco7941, w_eco7942, w_eco7943, w_eco7944, w_eco7945, w_eco7946, w_eco7947, w_eco7948, w_eco7949, w_eco7950, w_eco7951, w_eco7952, w_eco7953, w_eco7954, w_eco7955, w_eco7956, w_eco7957, w_eco7958, w_eco7959, w_eco7960, w_eco7961, w_eco7962, w_eco7963, w_eco7964, w_eco7965, w_eco7966, w_eco7967, w_eco7968, w_eco7969, w_eco7970, w_eco7971, w_eco7972, w_eco7973, w_eco7974, w_eco7975, w_eco7976, w_eco7977, w_eco7978, w_eco7979, w_eco7980, w_eco7981, w_eco7982, w_eco7983, w_eco7984, w_eco7985, w_eco7986, w_eco7987, w_eco7988, w_eco7989, w_eco7990, w_eco7991, w_eco7992, w_eco7993, w_eco7994, w_eco7995, w_eco7996, w_eco7997, w_eco7998, w_eco7999, w_eco8000, w_eco8001, w_eco8002, w_eco8003, w_eco8004, w_eco8005, w_eco8006, w_eco8007, w_eco8008, w_eco8009, w_eco8010, w_eco8011, w_eco8012, w_eco8013, w_eco8014, w_eco8015, w_eco8016, w_eco8017, w_eco8018, w_eco8019, w_eco8020, w_eco8021, w_eco8022, w_eco8023, w_eco8024, w_eco8025, w_eco8026, w_eco8027, w_eco8028, w_eco8029, w_eco8030, w_eco8031, w_eco8032, w_eco8033, w_eco8034, w_eco8035, w_eco8036, w_eco8037, w_eco8038, w_eco8039, w_eco8040, w_eco8041, w_eco8042, w_eco8043, w_eco8044, w_eco8045, w_eco8046, w_eco8047, w_eco8048, w_eco8049, w_eco8050, w_eco8051, w_eco8052, w_eco8053, w_eco8054, w_eco8055, w_eco8056, w_eco8057, w_eco8058, w_eco8059, w_eco8060, w_eco8061, w_eco8062, w_eco8063, w_eco8064, w_eco8065, w_eco8066, w_eco8067, w_eco8068, w_eco8069, w_eco8070, w_eco8071, w_eco8072, w_eco8073, w_eco8074, w_eco8075, w_eco8076, w_eco8077, w_eco8078, w_eco8079, w_eco8080, w_eco8081, w_eco8082, w_eco8083, w_eco8084, w_eco8085, w_eco8086, w_eco8087, w_eco8088, w_eco8089, w_eco8090, w_eco8091, w_eco8092, w_eco8093, w_eco8094, w_eco8095, w_eco8096, w_eco8097, w_eco8098, w_eco8099, w_eco8100, w_eco8101, w_eco8102, w_eco8103, w_eco8104, w_eco8105, w_eco8106, w_eco8107, w_eco8108, w_eco8109, w_eco8110, w_eco8111, w_eco8112, w_eco8113, w_eco8114, w_eco8115, w_eco8116, w_eco8117, w_eco8118, w_eco8119, w_eco8120, w_eco8121, w_eco8122, w_eco8123, w_eco8124, w_eco8125, w_eco8126, w_eco8127, w_eco8128, w_eco8129, w_eco8130, w_eco8131, w_eco8132, w_eco8133, w_eco8134, w_eco8135, w_eco8136, w_eco8137, w_eco8138, w_eco8139, w_eco8140, w_eco8141, w_eco8142, w_eco8143, w_eco8144, w_eco8145, w_eco8146, w_eco8147, w_eco8148, w_eco8149, w_eco8150, w_eco8151, w_eco8152, w_eco8153, w_eco8154, w_eco8155, w_eco8156, w_eco8157, w_eco8158, w_eco8159, w_eco8160, w_eco8161, w_eco8162, w_eco8163, w_eco8164, w_eco8165, w_eco8166, w_eco8167, w_eco8168, w_eco8169, w_eco8170, w_eco8171, w_eco8172, w_eco8173, w_eco8174, w_eco8175, w_eco8176, w_eco8177, w_eco8178, w_eco8179, w_eco8180, w_eco8181, w_eco8182, w_eco8183, w_eco8184, w_eco8185, w_eco8186, w_eco8187, w_eco8188, w_eco8189, w_eco8190, w_eco8191, w_eco8192, w_eco8193, w_eco8194, w_eco8195, w_eco8196, w_eco8197, w_eco8198, w_eco8199, w_eco8200, w_eco8201, w_eco8202, w_eco8203, w_eco8204, w_eco8205, w_eco8206, w_eco8207, w_eco8208, w_eco8209, w_eco8210, w_eco8211, w_eco8212, w_eco8213, w_eco8214, w_eco8215, w_eco8216, w_eco8217, w_eco8218, w_eco8219, w_eco8220, w_eco8221, w_eco8222, w_eco8223, w_eco8224, w_eco8225, w_eco8226, w_eco8227, w_eco8228, w_eco8229, w_eco8230, w_eco8231, w_eco8232, w_eco8233, w_eco8234, w_eco8235, w_eco8236, w_eco8237, w_eco8238, w_eco8239, w_eco8240, w_eco8241, w_eco8242, w_eco8243, w_eco8244, w_eco8245, w_eco8246, w_eco8247, w_eco8248, w_eco8249, w_eco8250, w_eco8251, w_eco8252, w_eco8253, w_eco8254, w_eco8255, w_eco8256, w_eco8257, w_eco8258, w_eco8259, w_eco8260, w_eco8261, w_eco8262, w_eco8263, w_eco8264, w_eco8265, w_eco8266, w_eco8267, w_eco8268, w_eco8269, w_eco8270, w_eco8271, w_eco8272, w_eco8273, w_eco8274, w_eco8275, w_eco8276, w_eco8277, w_eco8278, w_eco8279, w_eco8280, w_eco8281, w_eco8282, w_eco8283, w_eco8284, w_eco8285, w_eco8286, w_eco8287, w_eco8288, w_eco8289, w_eco8290, w_eco8291, w_eco8292, w_eco8293, w_eco8294, w_eco8295, w_eco8296, w_eco8297, w_eco8298, w_eco8299, w_eco8300, w_eco8301, w_eco8302, w_eco8303, w_eco8304, w_eco8305, w_eco8306, w_eco8307, w_eco8308, w_eco8309, w_eco8310, w_eco8311, w_eco8312, w_eco8313, w_eco8314, w_eco8315, w_eco8316, w_eco8317, w_eco8318, w_eco8319, w_eco8320, w_eco8321, w_eco8322, w_eco8323, w_eco8324, w_eco8325, w_eco8326, w_eco8327, w_eco8328, w_eco8329, w_eco8330, w_eco8331, w_eco8332, w_eco8333, w_eco8334, w_eco8335, w_eco8336, w_eco8337, w_eco8338, w_eco8339, w_eco8340, w_eco8341, w_eco8342, w_eco8343, w_eco8344, w_eco8345, w_eco8346, w_eco8347, w_eco8348, w_eco8349, w_eco8350, w_eco8351, w_eco8352, w_eco8353, w_eco8354, w_eco8355, w_eco8356, w_eco8357, w_eco8358, w_eco8359, w_eco8360, w_eco8361, w_eco8362, w_eco8363, w_eco8364, w_eco8365, w_eco8366, w_eco8367, w_eco8368, w_eco8369, w_eco8370, w_eco8371, w_eco8372, w_eco8373, w_eco8374, w_eco8375, w_eco8376, w_eco8377, w_eco8378, w_eco8379, w_eco8380, w_eco8381, w_eco8382, w_eco8383, w_eco8384, w_eco8385, w_eco8386, w_eco8387, w_eco8388, w_eco8389, w_eco8390, w_eco8391, w_eco8392, w_eco8393, w_eco8394, w_eco8395, w_eco8396, w_eco8397, w_eco8398, w_eco8399, w_eco8400, w_eco8401, w_eco8402, w_eco8403, w_eco8404, w_eco8405, w_eco8406, w_eco8407, w_eco8408, w_eco8409, w_eco8410, w_eco8411, w_eco8412, w_eco8413, w_eco8414, w_eco8415, w_eco8416, w_eco8417, w_eco8418, w_eco8419, w_eco8420, w_eco8421, w_eco8422, w_eco8423, w_eco8424, w_eco8425, w_eco8426, w_eco8427, w_eco8428, w_eco8429, w_eco8430, w_eco8431, w_eco8432, w_eco8433, w_eco8434, w_eco8435, w_eco8436, w_eco8437, w_eco8438, w_eco8439, w_eco8440, w_eco8441, w_eco8442, w_eco8443, w_eco8444, w_eco8445, w_eco8446, w_eco8447, w_eco8448, w_eco8449, w_eco8450, w_eco8451, w_eco8452, w_eco8453, w_eco8454, w_eco8455, w_eco8456, w_eco8457, w_eco8458, w_eco8459, w_eco8460, w_eco8461, w_eco8462, w_eco8463, w_eco8464, w_eco8465, w_eco8466, w_eco8467, w_eco8468, w_eco8469, w_eco8470, w_eco8471, w_eco8472, w_eco8473, w_eco8474, w_eco8475, w_eco8476, w_eco8477, w_eco8478, w_eco8479, w_eco8480, w_eco8481, w_eco8482, w_eco8483, w_eco8484, w_eco8485, w_eco8486, w_eco8487, w_eco8488, w_eco8489, w_eco8490, w_eco8491, w_eco8492, w_eco8493, w_eco8494, w_eco8495, w_eco8496, w_eco8497, w_eco8498, w_eco8499, w_eco8500, w_eco8501, w_eco8502, w_eco8503, w_eco8504, w_eco8505, w_eco8506, w_eco8507, w_eco8508, w_eco8509, w_eco8510, w_eco8511, w_eco8512, w_eco8513, w_eco8514, w_eco8515, w_eco8516, w_eco8517, w_eco8518, w_eco8519, w_eco8520, w_eco8521, w_eco8522, w_eco8523, w_eco8524, w_eco8525, w_eco8526, w_eco8527, w_eco8528, w_eco8529, w_eco8530, w_eco8531, w_eco8532, w_eco8533, w_eco8534, w_eco8535, w_eco8536, w_eco8537, w_eco8538, w_eco8539, w_eco8540, w_eco8541, w_eco8542, w_eco8543, w_eco8544, w_eco8545, w_eco8546, w_eco8547, w_eco8548, w_eco8549, w_eco8550, w_eco8551, w_eco8552, w_eco8553, w_eco8554, w_eco8555, w_eco8556, w_eco8557, w_eco8558, w_eco8559, w_eco8560, w_eco8561, w_eco8562, w_eco8563, w_eco8564, w_eco8565, w_eco8566, w_eco8567, w_eco8568, w_eco8569, w_eco8570, w_eco8571, w_eco8572, w_eco8573, w_eco8574, w_eco8575, w_eco8576, w_eco8577, w_eco8578, w_eco8579, w_eco8580, w_eco8581, w_eco8582, w_eco8583, w_eco8584, w_eco8585, w_eco8586, w_eco8587, w_eco8588, w_eco8589, w_eco8590, w_eco8591, w_eco8592, w_eco8593, w_eco8594, w_eco8595, w_eco8596, w_eco8597, w_eco8598, w_eco8599, w_eco8600, w_eco8601, w_eco8602, w_eco8603, w_eco8604, w_eco8605, w_eco8606, w_eco8607, w_eco8608, w_eco8609, w_eco8610, w_eco8611, w_eco8612, w_eco8613, w_eco8614, w_eco8615, w_eco8616, w_eco8617, w_eco8618, w_eco8619, w_eco8620, w_eco8621, w_eco8622, w_eco8623, w_eco8624, w_eco8625, w_eco8626, w_eco8627, w_eco8628, w_eco8629, w_eco8630, w_eco8631, w_eco8632, w_eco8633, w_eco8634, w_eco8635, w_eco8636, w_eco8637, w_eco8638, w_eco8639, w_eco8640, w_eco8641, w_eco8642, w_eco8643, w_eco8644, w_eco8645, w_eco8646, w_eco8647, w_eco8648, w_eco8649, w_eco8650, w_eco8651, w_eco8652, w_eco8653, w_eco8654, w_eco8655, w_eco8656, w_eco8657, w_eco8658, w_eco8659, w_eco8660, w_eco8661, w_eco8662, w_eco8663, w_eco8664, w_eco8665, w_eco8666, w_eco8667, w_eco8668, w_eco8669, w_eco8670, w_eco8671, w_eco8672, w_eco8673, w_eco8674, w_eco8675, w_eco8676, w_eco8677, w_eco8678, w_eco8679, w_eco8680, w_eco8681, w_eco8682, w_eco8683, w_eco8684, w_eco8685, w_eco8686, w_eco8687, w_eco8688, w_eco8689, w_eco8690, w_eco8691, w_eco8692, w_eco8693, w_eco8694, w_eco8695, w_eco8696, w_eco8697, w_eco8698, w_eco8699, w_eco8700, w_eco8701, w_eco8702, w_eco8703, w_eco8704, w_eco8705, w_eco8706, w_eco8707, w_eco8708, w_eco8709, w_eco8710, w_eco8711, w_eco8712, w_eco8713, w_eco8714, w_eco8715, w_eco8716, w_eco8717, w_eco8718, w_eco8719, w_eco8720, w_eco8721, w_eco8722, w_eco8723, w_eco8724, w_eco8725, w_eco8726, w_eco8727, w_eco8728, w_eco8729, w_eco8730, w_eco8731, w_eco8732, w_eco8733, w_eco8734, w_eco8735, w_eco8736, w_eco8737, w_eco8738, w_eco8739, w_eco8740, w_eco8741, w_eco8742, w_eco8743, w_eco8744, w_eco8745, w_eco8746, w_eco8747, w_eco8748, w_eco8749, w_eco8750, w_eco8751, w_eco8752, w_eco8753, w_eco8754, w_eco8755, w_eco8756, w_eco8757, w_eco8758, w_eco8759, w_eco8760, w_eco8761, w_eco8762, w_eco8763, w_eco8764, w_eco8765, w_eco8766, w_eco8767, w_eco8768, w_eco8769, w_eco8770, w_eco8771, w_eco8772, w_eco8773, w_eco8774, w_eco8775, w_eco8776, w_eco8777, w_eco8778, w_eco8779, w_eco8780, w_eco8781, w_eco8782, w_eco8783, w_eco8784, w_eco8785, w_eco8786, w_eco8787, w_eco8788, w_eco8789, w_eco8790, w_eco8791, w_eco8792, w_eco8793, w_eco8794, w_eco8795, w_eco8796, w_eco8797, w_eco8798, w_eco8799, w_eco8800, w_eco8801, w_eco8802, w_eco8803, w_eco8804, w_eco8805, w_eco8806, w_eco8807, w_eco8808, w_eco8809, w_eco8810, w_eco8811, w_eco8812, w_eco8813, w_eco8814, w_eco8815, w_eco8816, w_eco8817, w_eco8818, w_eco8819, w_eco8820, w_eco8821, w_eco8822, w_eco8823, w_eco8824, w_eco8825, w_eco8826, w_eco8827, w_eco8828, w_eco8829, w_eco8830, w_eco8831, w_eco8832, w_eco8833, w_eco8834, w_eco8835, w_eco8836, w_eco8837, w_eco8838, w_eco8839, w_eco8840, w_eco8841, w_eco8842, w_eco8843, w_eco8844, w_eco8845, w_eco8846, w_eco8847, w_eco8848, w_eco8849, w_eco8850, w_eco8851, w_eco8852, w_eco8853, w_eco8854, w_eco8855, w_eco8856, w_eco8857, w_eco8858, w_eco8859, w_eco8860, w_eco8861, w_eco8862, w_eco8863, w_eco8864, w_eco8865, w_eco8866, w_eco8867, w_eco8868, w_eco8869, w_eco8870, w_eco8871, w_eco8872, w_eco8873, w_eco8874, w_eco8875, w_eco8876, w_eco8877, w_eco8878, w_eco8879, w_eco8880, w_eco8881, w_eco8882, w_eco8883, w_eco8884, w_eco8885, w_eco8886, w_eco8887, w_eco8888, w_eco8889, w_eco8890, w_eco8891, w_eco8892, w_eco8893, w_eco8894, w_eco8895, w_eco8896, w_eco8897, w_eco8898, w_eco8899, w_eco8900, w_eco8901, w_eco8902, w_eco8903, w_eco8904, w_eco8905, w_eco8906, w_eco8907, w_eco8908, w_eco8909, w_eco8910, w_eco8911, w_eco8912, w_eco8913, w_eco8914, w_eco8915, w_eco8916, w_eco8917, w_eco8918, w_eco8919, w_eco8920, w_eco8921, w_eco8922, w_eco8923, w_eco8924, w_eco8925, w_eco8926, w_eco8927, w_eco8928, w_eco8929, w_eco8930, w_eco8931, w_eco8932, w_eco8933, w_eco8934, w_eco8935, w_eco8936, w_eco8937, w_eco8938, w_eco8939, w_eco8940, w_eco8941, w_eco8942, w_eco8943, w_eco8944, w_eco8945, w_eco8946, w_eco8947, w_eco8948, w_eco8949, w_eco8950, w_eco8951, w_eco8952, w_eco8953, w_eco8954, w_eco8955, w_eco8956, w_eco8957, w_eco8958, w_eco8959, w_eco8960, w_eco8961, w_eco8962, w_eco8963, w_eco8964, w_eco8965, w_eco8966, w_eco8967, w_eco8968, w_eco8969, w_eco8970, w_eco8971, w_eco8972, w_eco8973, w_eco8974, w_eco8975, w_eco8976, w_eco8977, w_eco8978, w_eco8979, w_eco8980, w_eco8981, w_eco8982, w_eco8983, w_eco8984, w_eco8985, w_eco8986, w_eco8987, w_eco8988, w_eco8989, w_eco8990, w_eco8991, w_eco8992, w_eco8993, w_eco8994, w_eco8995, w_eco8996, w_eco8997, w_eco8998, w_eco8999, w_eco9000, w_eco9001, w_eco9002, w_eco9003, w_eco9004, w_eco9005, w_eco9006, w_eco9007, w_eco9008, w_eco9009, w_eco9010, w_eco9011, w_eco9012, w_eco9013, w_eco9014, w_eco9015, w_eco9016, w_eco9017, w_eco9018, w_eco9019, w_eco9020, w_eco9021, w_eco9022, w_eco9023, w_eco9024, w_eco9025, w_eco9026, w_eco9027, w_eco9028, w_eco9029, w_eco9030, w_eco9031, w_eco9032, w_eco9033, w_eco9034, w_eco9035, w_eco9036, w_eco9037, w_eco9038, w_eco9039, w_eco9040, w_eco9041, w_eco9042, w_eco9043, w_eco9044, w_eco9045, w_eco9046, w_eco9047, w_eco9048, w_eco9049, w_eco9050, w_eco9051, w_eco9052, w_eco9053, w_eco9054, w_eco9055, w_eco9056, w_eco9057, w_eco9058, w_eco9059, w_eco9060, w_eco9061, w_eco9062, w_eco9063, w_eco9064, w_eco9065, w_eco9066, w_eco9067, w_eco9068, w_eco9069, w_eco9070, w_eco9071, w_eco9072, w_eco9073, w_eco9074, w_eco9075, w_eco9076, w_eco9077, w_eco9078, w_eco9079, w_eco9080, w_eco9081, w_eco9082, w_eco9083, w_eco9084, w_eco9085, w_eco9086, w_eco9087, w_eco9088, w_eco9089, w_eco9090, w_eco9091, w_eco9092, w_eco9093, w_eco9094, w_eco9095, w_eco9096, w_eco9097, w_eco9098, w_eco9099, w_eco9100, w_eco9101, w_eco9102, w_eco9103, w_eco9104, w_eco9105, w_eco9106, w_eco9107, w_eco9108, w_eco9109, w_eco9110, w_eco9111, w_eco9112, w_eco9113, w_eco9114, w_eco9115, w_eco9116, w_eco9117, w_eco9118, w_eco9119, w_eco9120, w_eco9121, w_eco9122, w_eco9123, w_eco9124, w_eco9125, w_eco9126, w_eco9127, w_eco9128, w_eco9129, w_eco9130, w_eco9131, w_eco9132, w_eco9133, w_eco9134, w_eco9135, w_eco9136, w_eco9137, w_eco9138, w_eco9139, w_eco9140, w_eco9141, w_eco9142, w_eco9143, w_eco9144, w_eco9145, w_eco9146, w_eco9147, w_eco9148, w_eco9149, w_eco9150, w_eco9151, w_eco9152, w_eco9153, w_eco9154, w_eco9155, w_eco9156, w_eco9157, w_eco9158, w_eco9159, w_eco9160, w_eco9161, w_eco9162, w_eco9163, w_eco9164, w_eco9165, w_eco9166, w_eco9167, w_eco9168, w_eco9169, w_eco9170, w_eco9171, w_eco9172, w_eco9173, w_eco9174, w_eco9175, w_eco9176, w_eco9177, w_eco9178, w_eco9179, w_eco9180, w_eco9181, w_eco9182, w_eco9183, w_eco9184, w_eco9185, w_eco9186, w_eco9187, w_eco9188, w_eco9189, w_eco9190, w_eco9191, w_eco9192, w_eco9193, w_eco9194, w_eco9195, w_eco9196, w_eco9197, w_eco9198, w_eco9199, w_eco9200, w_eco9201, w_eco9202, w_eco9203, w_eco9204, w_eco9205, w_eco9206, w_eco9207, w_eco9208, w_eco9209, w_eco9210, w_eco9211, w_eco9212, w_eco9213, w_eco9214, w_eco9215, w_eco9216, w_eco9217, w_eco9218, w_eco9219, w_eco9220, w_eco9221, w_eco9222, w_eco9223, w_eco9224, w_eco9225, w_eco9226, w_eco9227, w_eco9228, w_eco9229, w_eco9230, w_eco9231, w_eco9232, w_eco9233, w_eco9234, w_eco9235, w_eco9236, w_eco9237, w_eco9238, w_eco9239, w_eco9240, w_eco9241, w_eco9242, w_eco9243, w_eco9244, w_eco9245, w_eco9246, w_eco9247, w_eco9248, w_eco9249, w_eco9250, w_eco9251, w_eco9252, w_eco9253, w_eco9254, w_eco9255, w_eco9256, w_eco9257, w_eco9258, w_eco9259, w_eco9260, w_eco9261, w_eco9262, w_eco9263, w_eco9264, w_eco9265, w_eco9266, w_eco9267, w_eco9268, w_eco9269, w_eco9270, w_eco9271, w_eco9272, w_eco9273, w_eco9274, w_eco9275, w_eco9276, w_eco9277, w_eco9278, w_eco9279, w_eco9280, w_eco9281, w_eco9282, w_eco9283, w_eco9284, w_eco9285, w_eco9286, w_eco9287, w_eco9288, w_eco9289, w_eco9290, w_eco9291, w_eco9292, w_eco9293, w_eco9294, w_eco9295, w_eco9296, w_eco9297, w_eco9298, w_eco9299, w_eco9300, w_eco9301, w_eco9302, w_eco9303, w_eco9304, w_eco9305, w_eco9306, w_eco9307, w_eco9308, w_eco9309, w_eco9310, w_eco9311, w_eco9312, w_eco9313, w_eco9314, w_eco9315, w_eco9316, w_eco9317, w_eco9318, w_eco9319, w_eco9320, w_eco9321, w_eco9322, w_eco9323, w_eco9324, w_eco9325, w_eco9326, w_eco9327, w_eco9328, w_eco9329, w_eco9330, w_eco9331, w_eco9332, w_eco9333, w_eco9334, w_eco9335, w_eco9336, w_eco9337, w_eco9338, w_eco9339, w_eco9340, w_eco9341, w_eco9342, w_eco9343, w_eco9344, w_eco9345, w_eco9346, w_eco9347, w_eco9348, w_eco9349, w_eco9350, w_eco9351, w_eco9352, w_eco9353, w_eco9354, w_eco9355, w_eco9356, w_eco9357, w_eco9358, w_eco9359, w_eco9360, w_eco9361, w_eco9362, w_eco9363, w_eco9364, w_eco9365, w_eco9366, w_eco9367, w_eco9368, w_eco9369, w_eco9370, w_eco9371, w_eco9372, w_eco9373, w_eco9374, w_eco9375, w_eco9376, w_eco9377, w_eco9378, w_eco9379, w_eco9380, w_eco9381, w_eco9382, w_eco9383, w_eco9384, w_eco9385, w_eco9386, w_eco9387, w_eco9388, w_eco9389, w_eco9390, w_eco9391, w_eco9392, w_eco9393, w_eco9394, w_eco9395, w_eco9396, w_eco9397, w_eco9398, w_eco9399, w_eco9400, w_eco9401, w_eco9402, w_eco9403, w_eco9404, w_eco9405, w_eco9406, w_eco9407, w_eco9408, w_eco9409, w_eco9410, w_eco9411, w_eco9412, w_eco9413, w_eco9414, w_eco9415, w_eco9416, w_eco9417, w_eco9418, w_eco9419, w_eco9420, w_eco9421, w_eco9422, w_eco9423, w_eco9424, w_eco9425, w_eco9426, w_eco9427, w_eco9428, w_eco9429, w_eco9430, w_eco9431, w_eco9432, w_eco9433, w_eco9434, w_eco9435, w_eco9436, w_eco9437, w_eco9438, w_eco9439, w_eco9440, w_eco9441, w_eco9442, w_eco9443, w_eco9444, w_eco9445, w_eco9446, w_eco9447, w_eco9448, w_eco9449, w_eco9450, w_eco9451, w_eco9452, w_eco9453, w_eco9454, w_eco9455, w_eco9456, w_eco9457, w_eco9458, w_eco9459, w_eco9460, w_eco9461, w_eco9462, w_eco9463, w_eco9464, w_eco9465, w_eco9466, w_eco9467, w_eco9468, w_eco9469, w_eco9470, w_eco9471, w_eco9472, w_eco9473, w_eco9474, w_eco9475, w_eco9476, w_eco9477, w_eco9478, w_eco9479, w_eco9480, w_eco9481, w_eco9482, w_eco9483, w_eco9484, w_eco9485, w_eco9486, w_eco9487, w_eco9488, w_eco9489, w_eco9490, w_eco9491, w_eco9492, w_eco9493, w_eco9494, w_eco9495, w_eco9496, w_eco9497, w_eco9498, w_eco9499, w_eco9500, w_eco9501, w_eco9502, w_eco9503, w_eco9504, w_eco9505, w_eco9506, w_eco9507, w_eco9508, w_eco9509, w_eco9510, w_eco9511, w_eco9512, w_eco9513, w_eco9514, w_eco9515, w_eco9516, w_eco9517, w_eco9518, w_eco9519, w_eco9520, w_eco9521, w_eco9522, w_eco9523, w_eco9524, w_eco9525, w_eco9526, w_eco9527, w_eco9528, w_eco9529, w_eco9530, w_eco9531, w_eco9532, w_eco9533, w_eco9534, w_eco9535, w_eco9536, w_eco9537, w_eco9538, w_eco9539, w_eco9540, w_eco9541, w_eco9542, w_eco9543, w_eco9544, w_eco9545, w_eco9546, w_eco9547, w_eco9548, w_eco9549, w_eco9550, w_eco9551, w_eco9552, w_eco9553, w_eco9554, w_eco9555, w_eco9556, w_eco9557, w_eco9558, w_eco9559, w_eco9560, w_eco9561, w_eco9562, w_eco9563, w_eco9564, w_eco9565, w_eco9566, w_eco9567, w_eco9568, w_eco9569, w_eco9570, w_eco9571, w_eco9572, w_eco9573, w_eco9574, w_eco9575, w_eco9576, w_eco9577, w_eco9578, w_eco9579, w_eco9580, w_eco9581, w_eco9582, w_eco9583, w_eco9584, w_eco9585, w_eco9586, w_eco9587, w_eco9588, w_eco9589, w_eco9590, w_eco9591, w_eco9592, w_eco9593, w_eco9594, w_eco9595, w_eco9596, w_eco9597, w_eco9598, w_eco9599, w_eco9600, w_eco9601, w_eco9602, w_eco9603, w_eco9604, w_eco9605, w_eco9606, w_eco9607, w_eco9608, w_eco9609, w_eco9610, w_eco9611, w_eco9612, w_eco9613, w_eco9614, w_eco9615, w_eco9616, w_eco9617, w_eco9618, w_eco9619, w_eco9620, w_eco9621, w_eco9622, w_eco9623, w_eco9624, w_eco9625, w_eco9626, w_eco9627, w_eco9628, w_eco9629, w_eco9630, w_eco9631, w_eco9632, w_eco9633, w_eco9634, w_eco9635, w_eco9636, w_eco9637, w_eco9638, w_eco9639, w_eco9640, w_eco9641, w_eco9642, w_eco9643, w_eco9644, w_eco9645, w_eco9646, w_eco9647, w_eco9648, w_eco9649, w_eco9650, w_eco9651, w_eco9652, w_eco9653, w_eco9654, w_eco9655, w_eco9656, w_eco9657, w_eco9658, w_eco9659, w_eco9660, w_eco9661, w_eco9662, w_eco9663, w_eco9664, w_eco9665, w_eco9666, w_eco9667, w_eco9668, w_eco9669, w_eco9670, w_eco9671, w_eco9672, w_eco9673, w_eco9674, w_eco9675, w_eco9676, w_eco9677, w_eco9678, w_eco9679, w_eco9680, w_eco9681, w_eco9682, w_eco9683, w_eco9684, w_eco9685, w_eco9686, w_eco9687, w_eco9688, w_eco9689, w_eco9690, w_eco9691, w_eco9692, w_eco9693, w_eco9694, w_eco9695, w_eco9696, w_eco9697, w_eco9698, w_eco9699, w_eco9700, w_eco9701, w_eco9702, w_eco9703, w_eco9704, w_eco9705, w_eco9706, w_eco9707, w_eco9708, w_eco9709, w_eco9710, w_eco9711, w_eco9712, w_eco9713, w_eco9714, w_eco9715, w_eco9716, w_eco9717, w_eco9718, w_eco9719, w_eco9720, w_eco9721, w_eco9722, w_eco9723, w_eco9724, w_eco9725, w_eco9726, w_eco9727, w_eco9728, w_eco9729, w_eco9730, w_eco9731, w_eco9732, w_eco9733, w_eco9734, w_eco9735, w_eco9736, w_eco9737, w_eco9738, w_eco9739, w_eco9740, w_eco9741, w_eco9742, w_eco9743, w_eco9744, w_eco9745, w_eco9746, w_eco9747, w_eco9748, w_eco9749, w_eco9750, w_eco9751, w_eco9752, w_eco9753, w_eco9754, w_eco9755, w_eco9756, w_eco9757, w_eco9758, w_eco9759, w_eco9760, w_eco9761, w_eco9762, w_eco9763, w_eco9764, w_eco9765, w_eco9766, w_eco9767, w_eco9768, w_eco9769, w_eco9770, w_eco9771, w_eco9772, w_eco9773, w_eco9774, w_eco9775, w_eco9776, w_eco9777, w_eco9778, w_eco9779, w_eco9780, w_eco9781, w_eco9782, w_eco9783, w_eco9784, w_eco9785, w_eco9786, w_eco9787, w_eco9788, w_eco9789, w_eco9790, w_eco9791, w_eco9792, w_eco9793, w_eco9794, w_eco9795, w_eco9796, w_eco9797, w_eco9798, w_eco9799, w_eco9800, w_eco9801, w_eco9802, w_eco9803, w_eco9804, w_eco9805, w_eco9806, w_eco9807, w_eco9808, w_eco9809, w_eco9810, w_eco9811, w_eco9812, w_eco9813, w_eco9814, w_eco9815, w_eco9816, w_eco9817, w_eco9818, w_eco9819, w_eco9820, w_eco9821, w_eco9822, w_eco9823, w_eco9824, w_eco9825, w_eco9826, w_eco9827, w_eco9828, w_eco9829, w_eco9830, w_eco9831, w_eco9832, w_eco9833, w_eco9834, w_eco9835, w_eco9836, w_eco9837, w_eco9838, w_eco9839, w_eco9840, w_eco9841, w_eco9842, w_eco9843, w_eco9844, w_eco9845, w_eco9846, w_eco9847, w_eco9848, w_eco9849, w_eco9850, w_eco9851, w_eco9852, w_eco9853, w_eco9854, w_eco9855, w_eco9856, w_eco9857, w_eco9858, w_eco9859, w_eco9860, w_eco9861, w_eco9862, w_eco9863, w_eco9864, w_eco9865, w_eco9866, w_eco9867, w_eco9868, w_eco9869, w_eco9870, w_eco9871, w_eco9872, w_eco9873, w_eco9874, w_eco9875, w_eco9876, w_eco9877, w_eco9878, w_eco9879, w_eco9880, w_eco9881, w_eco9882, w_eco9883, w_eco9884, w_eco9885, w_eco9886, w_eco9887, w_eco9888, w_eco9889, w_eco9890, w_eco9891, w_eco9892, w_eco9893, w_eco9894, w_eco9895, w_eco9896, w_eco9897, w_eco9898, w_eco9899, w_eco9900, w_eco9901, w_eco9902, w_eco9903, w_eco9904, w_eco9905, w_eco9906, w_eco9907, w_eco9908, w_eco9909, w_eco9910, w_eco9911, w_eco9912, w_eco9913, w_eco9914, w_eco9915, w_eco9916, w_eco9917, w_eco9918, w_eco9919, w_eco9920, w_eco9921, w_eco9922, w_eco9923, w_eco9924, w_eco9925, w_eco9926, w_eco9927, w_eco9928, w_eco9929, w_eco9930, w_eco9931, w_eco9932, w_eco9933, w_eco9934, w_eco9935, w_eco9936, w_eco9937, w_eco9938, w_eco9939, w_eco9940, w_eco9941, w_eco9942, w_eco9943, w_eco9944, w_eco9945, w_eco9946, w_eco9947, w_eco9948, w_eco9949, w_eco9950, w_eco9951, w_eco9952, w_eco9953, w_eco9954, w_eco9955, w_eco9956, w_eco9957, w_eco9958, w_eco9959, w_eco9960, w_eco9961, w_eco9962, w_eco9963, w_eco9964, w_eco9965, w_eco9966, w_eco9967, w_eco9968, w_eco9969, w_eco9970, w_eco9971, w_eco9972, w_eco9973, w_eco9974, w_eco9975, w_eco9976, w_eco9977, w_eco9978, w_eco9979, w_eco9980, w_eco9981, w_eco9982, w_eco9983, w_eco9984, w_eco9985, w_eco9986, w_eco9987, w_eco9988, w_eco9989, w_eco9990, w_eco9991, w_eco9992, w_eco9993, w_eco9994, w_eco9995, w_eco9996, w_eco9997, w_eco9998, w_eco9999, w_eco10000, w_eco10001, w_eco10002, w_eco10003, w_eco10004, w_eco10005, w_eco10006, w_eco10007, w_eco10008, w_eco10009, w_eco10010, w_eco10011, w_eco10012, w_eco10013, w_eco10014, w_eco10015, w_eco10016, w_eco10017, w_eco10018, w_eco10019, w_eco10020, w_eco10021, w_eco10022, w_eco10023, w_eco10024, w_eco10025, w_eco10026, w_eco10027, w_eco10028, w_eco10029, w_eco10030, w_eco10031, w_eco10032, w_eco10033, w_eco10034, w_eco10035, w_eco10036, w_eco10037, w_eco10038, w_eco10039, w_eco10040, w_eco10041, w_eco10042, w_eco10043, w_eco10044, w_eco10045, w_eco10046, w_eco10047, w_eco10048, w_eco10049, w_eco10050, w_eco10051, w_eco10052, w_eco10053, w_eco10054, w_eco10055, w_eco10056, w_eco10057, w_eco10058, w_eco10059, w_eco10060, w_eco10061, w_eco10062, w_eco10063, w_eco10064, w_eco10065, w_eco10066, w_eco10067, w_eco10068, w_eco10069, w_eco10070, w_eco10071, w_eco10072, w_eco10073, w_eco10074, w_eco10075, w_eco10076, w_eco10077, w_eco10078, w_eco10079, w_eco10080, w_eco10081, w_eco10082, w_eco10083, w_eco10084, w_eco10085, w_eco10086, w_eco10087, w_eco10088, w_eco10089, w_eco10090, w_eco10091, w_eco10092, w_eco10093, w_eco10094, w_eco10095, w_eco10096, w_eco10097, w_eco10098, w_eco10099, w_eco10100, w_eco10101, w_eco10102, w_eco10103, w_eco10104, w_eco10105, w_eco10106, w_eco10107, w_eco10108, w_eco10109, w_eco10110, w_eco10111, w_eco10112, w_eco10113, w_eco10114, w_eco10115, w_eco10116, w_eco10117, w_eco10118, w_eco10119, w_eco10120, w_eco10121, w_eco10122, w_eco10123, w_eco10124, w_eco10125, w_eco10126, w_eco10127, w_eco10128, w_eco10129, w_eco10130, w_eco10131, w_eco10132, w_eco10133, w_eco10134, w_eco10135, w_eco10136, w_eco10137, w_eco10138, w_eco10139, w_eco10140, w_eco10141, w_eco10142, w_eco10143, w_eco10144, w_eco10145, w_eco10146, w_eco10147, w_eco10148, w_eco10149, w_eco10150, w_eco10151, w_eco10152, w_eco10153, w_eco10154, w_eco10155, w_eco10156, w_eco10157, w_eco10158, w_eco10159, w_eco10160, w_eco10161, w_eco10162, w_eco10163, w_eco10164, w_eco10165, w_eco10166, w_eco10167, w_eco10168, w_eco10169, w_eco10170, w_eco10171, w_eco10172, w_eco10173, w_eco10174, w_eco10175, w_eco10176, w_eco10177, w_eco10178, w_eco10179, w_eco10180, w_eco10181, w_eco10182, w_eco10183, w_eco10184, w_eco10185, w_eco10186, w_eco10187, w_eco10188, w_eco10189, w_eco10190, w_eco10191, w_eco10192, w_eco10193, w_eco10194, w_eco10195, w_eco10196, w_eco10197, w_eco10198, w_eco10199, w_eco10200, w_eco10201, w_eco10202, w_eco10203, w_eco10204, w_eco10205, w_eco10206, w_eco10207, w_eco10208, w_eco10209, w_eco10210, w_eco10211, w_eco10212, w_eco10213, w_eco10214, w_eco10215, w_eco10216, w_eco10217, w_eco10218, w_eco10219, w_eco10220, w_eco10221, w_eco10222, w_eco10223, w_eco10224, w_eco10225, w_eco10226, w_eco10227, w_eco10228, w_eco10229, w_eco10230, w_eco10231, w_eco10232, w_eco10233, w_eco10234, w_eco10235, w_eco10236, w_eco10237, w_eco10238, w_eco10239, w_eco10240, w_eco10241, w_eco10242, w_eco10243, w_eco10244, w_eco10245, w_eco10246, w_eco10247, w_eco10248, w_eco10249, w_eco10250, w_eco10251, w_eco10252, w_eco10253, w_eco10254, w_eco10255, w_eco10256, w_eco10257, w_eco10258, w_eco10259, w_eco10260, w_eco10261, w_eco10262, w_eco10263, w_eco10264, w_eco10265, w_eco10266, w_eco10267, w_eco10268, w_eco10269, w_eco10270, w_eco10271, w_eco10272, w_eco10273, w_eco10274, w_eco10275, w_eco10276, w_eco10277, w_eco10278, w_eco10279, w_eco10280, w_eco10281, w_eco10282, w_eco10283, w_eco10284, w_eco10285, w_eco10286, w_eco10287, w_eco10288, w_eco10289, w_eco10290, w_eco10291, w_eco10292, w_eco10293, w_eco10294, w_eco10295, w_eco10296, w_eco10297, w_eco10298, w_eco10299, w_eco10300, w_eco10301, w_eco10302, w_eco10303, w_eco10304, w_eco10305, w_eco10306, w_eco10307, w_eco10308, w_eco10309, w_eco10310, w_eco10311, w_eco10312, w_eco10313, w_eco10314, w_eco10315, w_eco10316, w_eco10317, w_eco10318, w_eco10319, w_eco10320, w_eco10321, w_eco10322, w_eco10323, w_eco10324, w_eco10325, w_eco10326, w_eco10327, w_eco10328, w_eco10329, w_eco10330, w_eco10331, w_eco10332, w_eco10333, w_eco10334, w_eco10335, w_eco10336, w_eco10337, w_eco10338, w_eco10339, w_eco10340, w_eco10341, w_eco10342, w_eco10343, w_eco10344, w_eco10345, w_eco10346, w_eco10347, w_eco10348, w_eco10349, w_eco10350, w_eco10351, w_eco10352, w_eco10353, w_eco10354, w_eco10355, w_eco10356, w_eco10357, w_eco10358, w_eco10359, w_eco10360, w_eco10361, w_eco10362, w_eco10363, w_eco10364, w_eco10365, w_eco10366, w_eco10367, w_eco10368, w_eco10369, w_eco10370, w_eco10371, w_eco10372, w_eco10373, w_eco10374, w_eco10375, w_eco10376, w_eco10377, w_eco10378, w_eco10379, w_eco10380, w_eco10381, w_eco10382, w_eco10383, w_eco10384, w_eco10385, w_eco10386, w_eco10387, w_eco10388, w_eco10389, w_eco10390, w_eco10391, w_eco10392, w_eco10393, w_eco10394, w_eco10395, w_eco10396, w_eco10397, w_eco10398, w_eco10399, w_eco10400, w_eco10401, w_eco10402, w_eco10403, w_eco10404, w_eco10405, w_eco10406, w_eco10407, w_eco10408, w_eco10409, w_eco10410, w_eco10411, w_eco10412, w_eco10413, w_eco10414, w_eco10415, w_eco10416, w_eco10417, w_eco10418, w_eco10419, w_eco10420, w_eco10421, w_eco10422, w_eco10423, w_eco10424, w_eco10425, w_eco10426, w_eco10427, w_eco10428, w_eco10429, w_eco10430, w_eco10431, w_eco10432, w_eco10433, w_eco10434, w_eco10435, w_eco10436, w_eco10437, w_eco10438, w_eco10439, w_eco10440, w_eco10441, w_eco10442, w_eco10443, w_eco10444, w_eco10445, w_eco10446, w_eco10447, w_eco10448, w_eco10449, w_eco10450, w_eco10451, w_eco10452, w_eco10453, w_eco10454, w_eco10455, w_eco10456, w_eco10457, w_eco10458, w_eco10459, w_eco10460, w_eco10461, w_eco10462, w_eco10463, w_eco10464, w_eco10465, w_eco10466, w_eco10467, w_eco10468, w_eco10469, w_eco10470, w_eco10471, w_eco10472, w_eco10473, w_eco10474, w_eco10475, w_eco10476, w_eco10477, w_eco10478, w_eco10479, w_eco10480, w_eco10481, w_eco10482, w_eco10483, w_eco10484, w_eco10485, w_eco10486, w_eco10487, w_eco10488, w_eco10489, w_eco10490, w_eco10491, w_eco10492, w_eco10493, w_eco10494, w_eco10495, w_eco10496, w_eco10497, w_eco10498, w_eco10499, w_eco10500, w_eco10501, w_eco10502, w_eco10503, w_eco10504, w_eco10505, w_eco10506, w_eco10507, w_eco10508, w_eco10509, w_eco10510, w_eco10511, w_eco10512, w_eco10513, w_eco10514, w_eco10515, w_eco10516, w_eco10517, w_eco10518, w_eco10519, w_eco10520, w_eco10521, w_eco10522, w_eco10523, w_eco10524, w_eco10525, w_eco10526, w_eco10527, w_eco10528, w_eco10529, w_eco10530, w_eco10531, w_eco10532, w_eco10533, w_eco10534, w_eco10535, w_eco10536, w_eco10537, w_eco10538, w_eco10539, w_eco10540, w_eco10541, w_eco10542, w_eco10543, w_eco10544, w_eco10545, w_eco10546, w_eco10547, w_eco10548, w_eco10549, w_eco10550, w_eco10551, w_eco10552, w_eco10553, w_eco10554, w_eco10555, w_eco10556, w_eco10557, w_eco10558, w_eco10559, w_eco10560, w_eco10561, w_eco10562, w_eco10563, w_eco10564, w_eco10565, w_eco10566, w_eco10567, w_eco10568, w_eco10569, w_eco10570, w_eco10571, w_eco10572, w_eco10573, w_eco10574, w_eco10575, w_eco10576, w_eco10577, w_eco10578, w_eco10579, w_eco10580, w_eco10581, w_eco10582, w_eco10583, w_eco10584, w_eco10585, w_eco10586, w_eco10587, w_eco10588, w_eco10589, w_eco10590, w_eco10591, w_eco10592, w_eco10593, w_eco10594, w_eco10595, w_eco10596, w_eco10597, w_eco10598, w_eco10599, w_eco10600, w_eco10601, w_eco10602, w_eco10603, w_eco10604, w_eco10605, w_eco10606, w_eco10607, w_eco10608, w_eco10609, w_eco10610, w_eco10611, w_eco10612, w_eco10613, w_eco10614, w_eco10615, w_eco10616, w_eco10617, w_eco10618, w_eco10619, w_eco10620, w_eco10621, w_eco10622, w_eco10623, w_eco10624, w_eco10625, w_eco10626, w_eco10627, w_eco10628, w_eco10629, w_eco10630, w_eco10631, w_eco10632, w_eco10633, w_eco10634, w_eco10635, w_eco10636, w_eco10637, w_eco10638, w_eco10639, w_eco10640, w_eco10641, w_eco10642, w_eco10643, w_eco10644, w_eco10645, w_eco10646, w_eco10647, w_eco10648, w_eco10649, w_eco10650, w_eco10651, w_eco10652, w_eco10653, w_eco10654, w_eco10655, w_eco10656, w_eco10657, w_eco10658, w_eco10659, w_eco10660, w_eco10661, w_eco10662, w_eco10663, w_eco10664, w_eco10665, w_eco10666, w_eco10667, w_eco10668, w_eco10669, w_eco10670, w_eco10671, w_eco10672, w_eco10673, w_eco10674, w_eco10675, w_eco10676, w_eco10677, w_eco10678, w_eco10679, w_eco10680, w_eco10681, w_eco10682, w_eco10683, w_eco10684, w_eco10685, w_eco10686, w_eco10687, w_eco10688, w_eco10689, w_eco10690, w_eco10691, w_eco10692, w_eco10693, w_eco10694, w_eco10695, w_eco10696, w_eco10697, w_eco10698, w_eco10699, w_eco10700, w_eco10701, w_eco10702, w_eco10703, w_eco10704, w_eco10705, w_eco10706, w_eco10707, w_eco10708, w_eco10709, w_eco10710, w_eco10711, w_eco10712, w_eco10713, w_eco10714, w_eco10715, w_eco10716, w_eco10717, w_eco10718, w_eco10719, w_eco10720, w_eco10721, w_eco10722, w_eco10723, w_eco10724, w_eco10725, w_eco10726, w_eco10727, w_eco10728, w_eco10729, w_eco10730, w_eco10731, w_eco10732, w_eco10733, w_eco10734, w_eco10735, w_eco10736, w_eco10737, w_eco10738, w_eco10739, w_eco10740, w_eco10741, w_eco10742, w_eco10743, w_eco10744, w_eco10745, w_eco10746, w_eco10747, w_eco10748, w_eco10749, w_eco10750, w_eco10751, w_eco10752, w_eco10753, w_eco10754, w_eco10755, w_eco10756, w_eco10757, w_eco10758, w_eco10759, w_eco10760, w_eco10761, w_eco10762, w_eco10763, w_eco10764, w_eco10765, w_eco10766, w_eco10767, w_eco10768, w_eco10769, w_eco10770, w_eco10771, w_eco10772, w_eco10773, w_eco10774, w_eco10775, w_eco10776, w_eco10777, w_eco10778, w_eco10779, w_eco10780, w_eco10781, w_eco10782, w_eco10783, w_eco10784, w_eco10785, w_eco10786, w_eco10787, w_eco10788, w_eco10789, w_eco10790, w_eco10791, w_eco10792, w_eco10793, w_eco10794, w_eco10795, w_eco10796, w_eco10797, w_eco10798, w_eco10799, w_eco10800, w_eco10801, w_eco10802, w_eco10803, w_eco10804, w_eco10805, w_eco10806, w_eco10807, w_eco10808, w_eco10809, w_eco10810, w_eco10811, w_eco10812, w_eco10813, w_eco10814, w_eco10815, w_eco10816, w_eco10817, w_eco10818, w_eco10819, w_eco10820, w_eco10821, w_eco10822, w_eco10823, w_eco10824, w_eco10825, w_eco10826, w_eco10827, w_eco10828, w_eco10829, w_eco10830, w_eco10831, w_eco10832, w_eco10833, w_eco10834, w_eco10835, w_eco10836, w_eco10837, w_eco10838, w_eco10839, w_eco10840, w_eco10841, w_eco10842, w_eco10843, w_eco10844, w_eco10845, w_eco10846, w_eco10847, w_eco10848, w_eco10849, w_eco10850, w_eco10851, w_eco10852, w_eco10853, w_eco10854, w_eco10855, w_eco10856, w_eco10857, w_eco10858, w_eco10859, w_eco10860, w_eco10861, w_eco10862, w_eco10863, w_eco10864, w_eco10865, w_eco10866, w_eco10867, w_eco10868, w_eco10869, w_eco10870, w_eco10871, w_eco10872, w_eco10873, w_eco10874, w_eco10875, w_eco10876, w_eco10877, w_eco10878, w_eco10879, w_eco10880, w_eco10881, w_eco10882, w_eco10883, w_eco10884, w_eco10885, w_eco10886, w_eco10887, w_eco10888, w_eco10889, w_eco10890, w_eco10891, w_eco10892, w_eco10893, w_eco10894, w_eco10895, w_eco10896, w_eco10897, w_eco10898, w_eco10899, w_eco10900, w_eco10901, w_eco10902, w_eco10903, w_eco10904, w_eco10905, w_eco10906, w_eco10907, w_eco10908, w_eco10909, w_eco10910, w_eco10911, w_eco10912, w_eco10913, w_eco10914, w_eco10915, w_eco10916, w_eco10917, w_eco10918, w_eco10919, w_eco10920, w_eco10921, w_eco10922, w_eco10923, w_eco10924, w_eco10925, w_eco10926, w_eco10927, w_eco10928, w_eco10929, w_eco10930, w_eco10931, w_eco10932, w_eco10933, w_eco10934, w_eco10935, w_eco10936, w_eco10937, w_eco10938, w_eco10939, w_eco10940, w_eco10941, w_eco10942, w_eco10943, w_eco10944, w_eco10945, w_eco10946, w_eco10947, w_eco10948, w_eco10949, w_eco10950, w_eco10951, w_eco10952, w_eco10953, w_eco10954, w_eco10955, w_eco10956, w_eco10957, w_eco10958, w_eco10959, w_eco10960, w_eco10961, w_eco10962, w_eco10963, w_eco10964, w_eco10965, w_eco10966, w_eco10967, w_eco10968, w_eco10969, w_eco10970, w_eco10971, w_eco10972, w_eco10973, w_eco10974, w_eco10975, w_eco10976, w_eco10977, w_eco10978, w_eco10979, w_eco10980, w_eco10981, w_eco10982, w_eco10983, w_eco10984, w_eco10985, w_eco10986, w_eco10987, w_eco10988, w_eco10989, w_eco10990, w_eco10991, w_eco10992, w_eco10993, w_eco10994, w_eco10995, w_eco10996, w_eco10997, w_eco10998, w_eco10999, w_eco11000, w_eco11001, w_eco11002, w_eco11003, w_eco11004, w_eco11005, w_eco11006, w_eco11007, w_eco11008, w_eco11009, w_eco11010, w_eco11011, w_eco11012, w_eco11013, w_eco11014, w_eco11015, w_eco11016, w_eco11017, w_eco11018, w_eco11019, w_eco11020, w_eco11021, w_eco11022, w_eco11023, w_eco11024, w_eco11025, w_eco11026, w_eco11027, w_eco11028, w_eco11029, w_eco11030, w_eco11031, w_eco11032, w_eco11033, w_eco11034, w_eco11035, w_eco11036, w_eco11037, w_eco11038, w_eco11039, w_eco11040, w_eco11041, w_eco11042, w_eco11043, w_eco11044, w_eco11045, w_eco11046, w_eco11047, w_eco11048, w_eco11049, w_eco11050, w_eco11051, w_eco11052, w_eco11053, w_eco11054, w_eco11055, w_eco11056, w_eco11057, w_eco11058, w_eco11059, w_eco11060, w_eco11061, w_eco11062, w_eco11063, w_eco11064, w_eco11065, w_eco11066, w_eco11067, w_eco11068, w_eco11069, w_eco11070, w_eco11071, w_eco11072, w_eco11073, w_eco11074, w_eco11075, w_eco11076, w_eco11077, w_eco11078, w_eco11079, w_eco11080, w_eco11081, w_eco11082, w_eco11083, w_eco11084, w_eco11085, w_eco11086, w_eco11087, w_eco11088, w_eco11089, w_eco11090, w_eco11091, w_eco11092, w_eco11093, w_eco11094, w_eco11095, w_eco11096, w_eco11097, w_eco11098, w_eco11099, w_eco11100, w_eco11101, w_eco11102, w_eco11103, w_eco11104, w_eco11105, w_eco11106, w_eco11107, w_eco11108, w_eco11109, w_eco11110, w_eco11111, w_eco11112, w_eco11113, w_eco11114, w_eco11115, w_eco11116, w_eco11117, w_eco11118, w_eco11119, w_eco11120, w_eco11121, w_eco11122, w_eco11123, w_eco11124, w_eco11125, w_eco11126, w_eco11127, w_eco11128, w_eco11129, w_eco11130, w_eco11131, w_eco11132, w_eco11133, w_eco11134, w_eco11135, w_eco11136, w_eco11137, w_eco11138, w_eco11139, w_eco11140, w_eco11141, w_eco11142, w_eco11143, w_eco11144, w_eco11145, w_eco11146, w_eco11147, w_eco11148, w_eco11149, w_eco11150, w_eco11151, w_eco11152, w_eco11153, w_eco11154, w_eco11155, w_eco11156, w_eco11157, w_eco11158, w_eco11159, w_eco11160, w_eco11161, w_eco11162, w_eco11163, w_eco11164, w_eco11165, w_eco11166, w_eco11167, w_eco11168, w_eco11169, w_eco11170, w_eco11171, w_eco11172, w_eco11173, w_eco11174, w_eco11175, w_eco11176, w_eco11177, w_eco11178, w_eco11179, w_eco11180, w_eco11181, w_eco11182, w_eco11183, w_eco11184, w_eco11185, w_eco11186, w_eco11187, w_eco11188, w_eco11189, w_eco11190, w_eco11191, w_eco11192, w_eco11193, w_eco11194, w_eco11195, w_eco11196, w_eco11197, w_eco11198, w_eco11199, w_eco11200, w_eco11201, w_eco11202, w_eco11203, w_eco11204, w_eco11205, w_eco11206, w_eco11207, w_eco11208, w_eco11209, w_eco11210, w_eco11211, w_eco11212, w_eco11213, w_eco11214, w_eco11215, w_eco11216, w_eco11217, w_eco11218, w_eco11219, w_eco11220, w_eco11221, w_eco11222, w_eco11223, w_eco11224, w_eco11225, w_eco11226, w_eco11227, w_eco11228, w_eco11229, w_eco11230, w_eco11231, w_eco11232, w_eco11233, w_eco11234, w_eco11235, w_eco11236, w_eco11237, w_eco11238, w_eco11239, w_eco11240, w_eco11241, w_eco11242, w_eco11243, w_eco11244, w_eco11245, w_eco11246, w_eco11247, w_eco11248, w_eco11249, w_eco11250, w_eco11251, w_eco11252, w_eco11253, w_eco11254, w_eco11255, w_eco11256, w_eco11257, w_eco11258, w_eco11259, w_eco11260, w_eco11261, w_eco11262, w_eco11263, w_eco11264, w_eco11265, w_eco11266, w_eco11267, w_eco11268, w_eco11269, w_eco11270, w_eco11271, w_eco11272, w_eco11273, w_eco11274, w_eco11275, w_eco11276, w_eco11277, w_eco11278, w_eco11279, w_eco11280, w_eco11281, w_eco11282, w_eco11283, w_eco11284, w_eco11285, w_eco11286, w_eco11287, w_eco11288, w_eco11289, w_eco11290, w_eco11291, w_eco11292, w_eco11293, w_eco11294, w_eco11295, w_eco11296, w_eco11297, w_eco11298, w_eco11299, w_eco11300, w_eco11301, w_eco11302, w_eco11303, w_eco11304, w_eco11305, w_eco11306, w_eco11307, w_eco11308, w_eco11309, w_eco11310, w_eco11311, w_eco11312, w_eco11313, w_eco11314, w_eco11315, w_eco11316, w_eco11317, w_eco11318, w_eco11319, w_eco11320, w_eco11321, w_eco11322, w_eco11323, w_eco11324, w_eco11325, w_eco11326, w_eco11327, w_eco11328, w_eco11329, w_eco11330, w_eco11331, w_eco11332, w_eco11333, w_eco11334, w_eco11335, w_eco11336, w_eco11337, w_eco11338, w_eco11339, w_eco11340, w_eco11341, w_eco11342, w_eco11343, w_eco11344, w_eco11345, w_eco11346, w_eco11347, w_eco11348, w_eco11349, w_eco11350, w_eco11351, w_eco11352, w_eco11353, w_eco11354, w_eco11355, w_eco11356, w_eco11357, w_eco11358, w_eco11359, w_eco11360, w_eco11361, w_eco11362, w_eco11363, w_eco11364, w_eco11365, w_eco11366, w_eco11367, w_eco11368, w_eco11369, w_eco11370, w_eco11371, w_eco11372, w_eco11373, w_eco11374, w_eco11375, w_eco11376, w_eco11377, w_eco11378, w_eco11379, w_eco11380, w_eco11381, w_eco11382, w_eco11383, w_eco11384, w_eco11385, w_eco11386, w_eco11387, w_eco11388, w_eco11389, w_eco11390, w_eco11391, w_eco11392, w_eco11393, w_eco11394, w_eco11395, w_eco11396, w_eco11397, w_eco11398, w_eco11399, w_eco11400, w_eco11401, w_eco11402, w_eco11403, w_eco11404, w_eco11405, w_eco11406, w_eco11407, w_eco11408, w_eco11409, w_eco11410, w_eco11411, w_eco11412, w_eco11413, w_eco11414, w_eco11415, w_eco11416, w_eco11417, w_eco11418, w_eco11419, w_eco11420, w_eco11421, w_eco11422, w_eco11423, w_eco11424, w_eco11425, w_eco11426, w_eco11427, w_eco11428, w_eco11429, w_eco11430, w_eco11431, w_eco11432, w_eco11433, w_eco11434, w_eco11435, w_eco11436, w_eco11437, w_eco11438, w_eco11439, w_eco11440, w_eco11441, w_eco11442, w_eco11443, w_eco11444, w_eco11445, w_eco11446, w_eco11447, w_eco11448, w_eco11449, w_eco11450, w_eco11451, w_eco11452, w_eco11453, w_eco11454, w_eco11455, w_eco11456, w_eco11457, w_eco11458, w_eco11459, w_eco11460, w_eco11461, w_eco11462, w_eco11463, w_eco11464, w_eco11465, w_eco11466, w_eco11467, w_eco11468, w_eco11469, w_eco11470, w_eco11471, w_eco11472, w_eco11473, w_eco11474, w_eco11475, w_eco11476, w_eco11477, w_eco11478, w_eco11479, w_eco11480, w_eco11481, w_eco11482, w_eco11483, w_eco11484, w_eco11485, w_eco11486, w_eco11487, w_eco11488, w_eco11489, w_eco11490, w_eco11491, w_eco11492, w_eco11493, w_eco11494, w_eco11495, w_eco11496, w_eco11497, w_eco11498, w_eco11499, w_eco11500, w_eco11501, w_eco11502, w_eco11503, w_eco11504, w_eco11505, w_eco11506, w_eco11507, w_eco11508, w_eco11509, w_eco11510, w_eco11511, w_eco11512, w_eco11513, w_eco11514, w_eco11515, w_eco11516, w_eco11517, w_eco11518, w_eco11519, w_eco11520, w_eco11521, w_eco11522, w_eco11523, w_eco11524, w_eco11525, w_eco11526, w_eco11527, w_eco11528, w_eco11529, w_eco11530, w_eco11531, w_eco11532, w_eco11533, w_eco11534, w_eco11535, w_eco11536, w_eco11537, w_eco11538, w_eco11539, w_eco11540, w_eco11541, w_eco11542, w_eco11543, w_eco11544, w_eco11545, w_eco11546, w_eco11547, w_eco11548, w_eco11549, w_eco11550, w_eco11551, w_eco11552, w_eco11553, w_eco11554, w_eco11555, w_eco11556, w_eco11557, w_eco11558, w_eco11559, w_eco11560, w_eco11561, w_eco11562, w_eco11563, w_eco11564, w_eco11565, w_eco11566, w_eco11567, w_eco11568, w_eco11569, w_eco11570, w_eco11571, w_eco11572, w_eco11573, w_eco11574, w_eco11575, w_eco11576, w_eco11577, w_eco11578, w_eco11579, w_eco11580, w_eco11581, w_eco11582, w_eco11583, w_eco11584, w_eco11585, w_eco11586, w_eco11587, w_eco11588, w_eco11589, w_eco11590, w_eco11591, w_eco11592, w_eco11593, w_eco11594, w_eco11595, w_eco11596, w_eco11597, w_eco11598, w_eco11599, w_eco11600, w_eco11601, w_eco11602, w_eco11603, w_eco11604, w_eco11605, w_eco11606, w_eco11607, w_eco11608, w_eco11609, w_eco11610, w_eco11611, w_eco11612, w_eco11613, w_eco11614, w_eco11615, w_eco11616, w_eco11617, w_eco11618, w_eco11619, w_eco11620, w_eco11621, w_eco11622, w_eco11623, w_eco11624, w_eco11625, w_eco11626, w_eco11627, w_eco11628, w_eco11629, w_eco11630, w_eco11631, w_eco11632, w_eco11633, w_eco11634, w_eco11635, w_eco11636, w_eco11637, w_eco11638, w_eco11639, w_eco11640, w_eco11641, w_eco11642, w_eco11643, w_eco11644, w_eco11645, w_eco11646, w_eco11647, w_eco11648, w_eco11649, w_eco11650, w_eco11651, w_eco11652, w_eco11653, w_eco11654, w_eco11655, w_eco11656, w_eco11657, w_eco11658, w_eco11659, w_eco11660, w_eco11661, w_eco11662, w_eco11663, w_eco11664, w_eco11665, w_eco11666, w_eco11667, w_eco11668, w_eco11669, w_eco11670, w_eco11671, w_eco11672, w_eco11673, w_eco11674, w_eco11675, w_eco11676, w_eco11677, w_eco11678, w_eco11679, w_eco11680, w_eco11681, w_eco11682, w_eco11683, w_eco11684, w_eco11685, w_eco11686, w_eco11687, w_eco11688, w_eco11689, w_eco11690, w_eco11691, w_eco11692, w_eco11693, w_eco11694, w_eco11695, w_eco11696, w_eco11697, w_eco11698, w_eco11699, w_eco11700, w_eco11701, w_eco11702, w_eco11703, w_eco11704, w_eco11705, w_eco11706, w_eco11707, w_eco11708, w_eco11709, w_eco11710, w_eco11711, w_eco11712, w_eco11713, w_eco11714, w_eco11715, w_eco11716, w_eco11717, w_eco11718, w_eco11719, w_eco11720, w_eco11721, w_eco11722, w_eco11723, w_eco11724, w_eco11725, w_eco11726, w_eco11727, w_eco11728, w_eco11729, w_eco11730, w_eco11731, w_eco11732, w_eco11733, w_eco11734, w_eco11735, w_eco11736, w_eco11737, w_eco11738, w_eco11739, w_eco11740, w_eco11741, w_eco11742, w_eco11743, w_eco11744, w_eco11745, w_eco11746, w_eco11747, w_eco11748, w_eco11749, w_eco11750, w_eco11751, w_eco11752, w_eco11753, w_eco11754, w_eco11755, w_eco11756, w_eco11757, w_eco11758, w_eco11759, w_eco11760, w_eco11761, w_eco11762, w_eco11763, w_eco11764, w_eco11765, w_eco11766, w_eco11767, w_eco11768, w_eco11769, w_eco11770, w_eco11771, w_eco11772, w_eco11773, w_eco11774, w_eco11775, w_eco11776, w_eco11777, w_eco11778, w_eco11779, w_eco11780, w_eco11781, w_eco11782, w_eco11783, w_eco11784, w_eco11785, w_eco11786, w_eco11787, w_eco11788, w_eco11789, w_eco11790, w_eco11791, w_eco11792, w_eco11793, w_eco11794, w_eco11795, w_eco11796, w_eco11797, w_eco11798, w_eco11799, w_eco11800, w_eco11801, w_eco11802, w_eco11803, w_eco11804, w_eco11805, w_eco11806, w_eco11807, w_eco11808, w_eco11809, w_eco11810, w_eco11811, w_eco11812, w_eco11813, w_eco11814, w_eco11815, w_eco11816, w_eco11817, w_eco11818, w_eco11819, w_eco11820, w_eco11821, w_eco11822, w_eco11823, w_eco11824, w_eco11825, w_eco11826, w_eco11827, w_eco11828, w_eco11829, w_eco11830, w_eco11831, w_eco11832, w_eco11833, w_eco11834, w_eco11835, w_eco11836, w_eco11837, w_eco11838, w_eco11839, w_eco11840, w_eco11841, w_eco11842, w_eco11843, w_eco11844, w_eco11845, w_eco11846, w_eco11847, w_eco11848, w_eco11849, w_eco11850, w_eco11851, w_eco11852, w_eco11853, w_eco11854, w_eco11855, w_eco11856, w_eco11857, w_eco11858, w_eco11859, w_eco11860, w_eco11861, w_eco11862, w_eco11863, w_eco11864, w_eco11865, w_eco11866, w_eco11867, w_eco11868, w_eco11869, w_eco11870, w_eco11871, w_eco11872, w_eco11873, w_eco11874, w_eco11875, w_eco11876, w_eco11877, w_eco11878, w_eco11879, w_eco11880, w_eco11881, w_eco11882, w_eco11883, w_eco11884, w_eco11885, w_eco11886, w_eco11887, w_eco11888, w_eco11889, w_eco11890, w_eco11891, w_eco11892, w_eco11893, w_eco11894, w_eco11895, w_eco11896, w_eco11897, w_eco11898, w_eco11899, w_eco11900, w_eco11901, w_eco11902, w_eco11903, w_eco11904, w_eco11905, w_eco11906, w_eco11907, w_eco11908, w_eco11909, w_eco11910, w_eco11911, w_eco11912, w_eco11913, w_eco11914, w_eco11915, w_eco11916, w_eco11917, w_eco11918, w_eco11919, w_eco11920, w_eco11921, w_eco11922, w_eco11923, w_eco11924, w_eco11925, w_eco11926, w_eco11927, w_eco11928, w_eco11929, w_eco11930, w_eco11931, w_eco11932, w_eco11933, w_eco11934, w_eco11935, w_eco11936, w_eco11937, w_eco11938, w_eco11939, w_eco11940, w_eco11941, w_eco11942, w_eco11943, w_eco11944, w_eco11945, w_eco11946, w_eco11947, w_eco11948, w_eco11949, w_eco11950, w_eco11951, w_eco11952, w_eco11953, w_eco11954, w_eco11955, w_eco11956, w_eco11957, w_eco11958, w_eco11959, w_eco11960, w_eco11961, w_eco11962, w_eco11963, w_eco11964, w_eco11965, w_eco11966, w_eco11967, w_eco11968, w_eco11969, w_eco11970, w_eco11971, w_eco11972, w_eco11973, w_eco11974, w_eco11975, w_eco11976, w_eco11977, w_eco11978, w_eco11979, w_eco11980, w_eco11981, w_eco11982, w_eco11983, w_eco11984, w_eco11985, w_eco11986, w_eco11987, w_eco11988, w_eco11989, w_eco11990, w_eco11991, w_eco11992, w_eco11993, w_eco11994, w_eco11995, w_eco11996, w_eco11997, w_eco11998, w_eco11999, w_eco12000, w_eco12001, w_eco12002, w_eco12003, w_eco12004, w_eco12005, w_eco12006, w_eco12007, w_eco12008, w_eco12009, w_eco12010, w_eco12011, w_eco12012, w_eco12013, w_eco12014, w_eco12015, w_eco12016, w_eco12017, w_eco12018, w_eco12019, w_eco12020, w_eco12021, w_eco12022, w_eco12023, w_eco12024, w_eco12025, w_eco12026, w_eco12027, w_eco12028, w_eco12029, w_eco12030, w_eco12031, w_eco12032, w_eco12033, w_eco12034, w_eco12035, w_eco12036, w_eco12037, w_eco12038, w_eco12039, w_eco12040, w_eco12041, w_eco12042, w_eco12043, w_eco12044, w_eco12045, w_eco12046, w_eco12047, w_eco12048, w_eco12049, w_eco12050, w_eco12051, w_eco12052, w_eco12053, w_eco12054, w_eco12055, w_eco12056, w_eco12057, w_eco12058, w_eco12059, w_eco12060, w_eco12061, w_eco12062, w_eco12063, w_eco12064, w_eco12065, w_eco12066, w_eco12067, w_eco12068, w_eco12069, w_eco12070, w_eco12071, w_eco12072, w_eco12073, w_eco12074, w_eco12075, w_eco12076, w_eco12077, w_eco12078, w_eco12079, w_eco12080, w_eco12081, w_eco12082, w_eco12083, w_eco12084, w_eco12085, w_eco12086, w_eco12087, w_eco12088, w_eco12089, w_eco12090, w_eco12091, w_eco12092, w_eco12093, w_eco12094, w_eco12095, w_eco12096, w_eco12097, w_eco12098, w_eco12099, w_eco12100, w_eco12101, w_eco12102, w_eco12103, w_eco12104, w_eco12105, w_eco12106, w_eco12107, w_eco12108, w_eco12109, w_eco12110, w_eco12111, w_eco12112, w_eco12113, w_eco12114, w_eco12115, w_eco12116, w_eco12117, w_eco12118, w_eco12119, w_eco12120, w_eco12121, w_eco12122, w_eco12123, w_eco12124, w_eco12125, w_eco12126, w_eco12127, w_eco12128, w_eco12129, w_eco12130, w_eco12131, w_eco12132, w_eco12133, w_eco12134, w_eco12135, w_eco12136, w_eco12137, w_eco12138, w_eco12139, w_eco12140, w_eco12141, w_eco12142, w_eco12143, w_eco12144, w_eco12145, w_eco12146, w_eco12147, w_eco12148, w_eco12149, w_eco12150, w_eco12151, w_eco12152, w_eco12153, w_eco12154, w_eco12155, w_eco12156, w_eco12157, w_eco12158, w_eco12159, w_eco12160, w_eco12161, w_eco12162, w_eco12163, w_eco12164, w_eco12165, w_eco12166, w_eco12167, w_eco12168, w_eco12169, w_eco12170, w_eco12171, w_eco12172, w_eco12173, w_eco12174, w_eco12175, w_eco12176, w_eco12177, w_eco12178, w_eco12179, w_eco12180, w_eco12181, w_eco12182, w_eco12183, w_eco12184, w_eco12185, w_eco12186, w_eco12187, w_eco12188, w_eco12189, w_eco12190, w_eco12191, w_eco12192, w_eco12193, w_eco12194, w_eco12195, w_eco12196, w_eco12197, w_eco12198, w_eco12199, w_eco12200, w_eco12201, w_eco12202, w_eco12203, w_eco12204, w_eco12205, w_eco12206, w_eco12207, w_eco12208, w_eco12209, w_eco12210, w_eco12211, w_eco12212, w_eco12213, w_eco12214, w_eco12215, w_eco12216, w_eco12217, w_eco12218, w_eco12219, w_eco12220, w_eco12221, w_eco12222, w_eco12223, w_eco12224, w_eco12225, w_eco12226, w_eco12227, w_eco12228, w_eco12229, w_eco12230, w_eco12231, w_eco12232, w_eco12233, w_eco12234, w_eco12235, w_eco12236, w_eco12237, w_eco12238, w_eco12239, w_eco12240, w_eco12241, w_eco12242, w_eco12243, w_eco12244, w_eco12245, w_eco12246, w_eco12247, w_eco12248, w_eco12249, w_eco12250, w_eco12251, w_eco12252, w_eco12253, w_eco12254, w_eco12255, w_eco12256, w_eco12257, w_eco12258, w_eco12259, w_eco12260, w_eco12261, w_eco12262, w_eco12263, w_eco12264, w_eco12265, w_eco12266, w_eco12267, w_eco12268, w_eco12269, w_eco12270, w_eco12271, w_eco12272, w_eco12273, w_eco12274, w_eco12275, w_eco12276, w_eco12277, w_eco12278, w_eco12279, w_eco12280, w_eco12281, w_eco12282, w_eco12283, w_eco12284, w_eco12285, w_eco12286, w_eco12287, w_eco12288, w_eco12289, w_eco12290, w_eco12291, w_eco12292, w_eco12293, w_eco12294, w_eco12295, w_eco12296, w_eco12297, w_eco12298, w_eco12299, w_eco12300, w_eco12301, w_eco12302, w_eco12303, w_eco12304, w_eco12305, w_eco12306, w_eco12307, w_eco12308, w_eco12309, w_eco12310, w_eco12311, w_eco12312, w_eco12313, w_eco12314, w_eco12315, w_eco12316, w_eco12317, w_eco12318, w_eco12319, w_eco12320, w_eco12321, w_eco12322, w_eco12323, w_eco12324, w_eco12325, w_eco12326, w_eco12327, w_eco12328, w_eco12329, w_eco12330, w_eco12331, w_eco12332, w_eco12333, w_eco12334, w_eco12335, w_eco12336, w_eco12337, w_eco12338, w_eco12339, w_eco12340, w_eco12341, w_eco12342, w_eco12343, w_eco12344, w_eco12345, w_eco12346, w_eco12347, w_eco12348, w_eco12349, w_eco12350, w_eco12351, w_eco12352, w_eco12353, w_eco12354, w_eco12355, w_eco12356, w_eco12357, w_eco12358, w_eco12359, w_eco12360, w_eco12361, w_eco12362, w_eco12363, w_eco12364, w_eco12365, w_eco12366, w_eco12367, w_eco12368, w_eco12369, w_eco12370, w_eco12371, w_eco12372, w_eco12373, w_eco12374, w_eco12375, w_eco12376, w_eco12377, w_eco12378, w_eco12379, w_eco12380, w_eco12381, w_eco12382, w_eco12383, w_eco12384, w_eco12385, w_eco12386, w_eco12387, w_eco12388, w_eco12389, w_eco12390, w_eco12391, w_eco12392, w_eco12393, w_eco12394, w_eco12395, w_eco12396, w_eco12397, w_eco12398, w_eco12399, w_eco12400, w_eco12401, w_eco12402, w_eco12403, w_eco12404, w_eco12405, w_eco12406, w_eco12407, w_eco12408, w_eco12409, w_eco12410, w_eco12411, w_eco12412, w_eco12413, w_eco12414, w_eco12415, w_eco12416, w_eco12417, w_eco12418, w_eco12419, w_eco12420, w_eco12421, w_eco12422, w_eco12423, w_eco12424, w_eco12425, w_eco12426, w_eco12427, w_eco12428, w_eco12429, w_eco12430, w_eco12431, w_eco12432, w_eco12433, w_eco12434, w_eco12435, w_eco12436, w_eco12437, w_eco12438, w_eco12439, w_eco12440, w_eco12441, w_eco12442, w_eco12443, w_eco12444, w_eco12445, w_eco12446, w_eco12447, w_eco12448, w_eco12449, w_eco12450, w_eco12451, w_eco12452, w_eco12453, w_eco12454, w_eco12455, w_eco12456, w_eco12457, w_eco12458, w_eco12459, w_eco12460, w_eco12461, w_eco12462, w_eco12463, w_eco12464, w_eco12465, w_eco12466, w_eco12467, w_eco12468, w_eco12469, w_eco12470, w_eco12471, w_eco12472, w_eco12473, w_eco12474, w_eco12475, w_eco12476, w_eco12477, w_eco12478, w_eco12479, w_eco12480, w_eco12481, w_eco12482, w_eco12483, w_eco12484, w_eco12485, w_eco12486, w_eco12487, w_eco12488, w_eco12489, w_eco12490, w_eco12491, w_eco12492, w_eco12493, w_eco12494, w_eco12495, w_eco12496, w_eco12497, w_eco12498, w_eco12499, w_eco12500, w_eco12501, w_eco12502, w_eco12503, w_eco12504, w_eco12505, w_eco12506, w_eco12507, w_eco12508, w_eco12509, w_eco12510, w_eco12511, w_eco12512, w_eco12513, w_eco12514, w_eco12515, w_eco12516, w_eco12517, w_eco12518, w_eco12519, w_eco12520, w_eco12521, w_eco12522, w_eco12523, w_eco12524, w_eco12525, w_eco12526, w_eco12527, w_eco12528, w_eco12529, w_eco12530, w_eco12531, w_eco12532, w_eco12533, w_eco12534, w_eco12535, w_eco12536, w_eco12537, w_eco12538, w_eco12539, w_eco12540, w_eco12541, w_eco12542, w_eco12543, w_eco12544, w_eco12545, w_eco12546, w_eco12547, w_eco12548, w_eco12549, w_eco12550, w_eco12551, w_eco12552, w_eco12553, w_eco12554, w_eco12555, w_eco12556, w_eco12557, w_eco12558, w_eco12559, w_eco12560, w_eco12561, w_eco12562, w_eco12563, w_eco12564, w_eco12565, w_eco12566, w_eco12567, w_eco12568, w_eco12569, w_eco12570, w_eco12571, w_eco12572, w_eco12573, w_eco12574, w_eco12575, w_eco12576, w_eco12577, w_eco12578, w_eco12579, w_eco12580, w_eco12581, w_eco12582, w_eco12583, w_eco12584, w_eco12585, w_eco12586, w_eco12587, w_eco12588, w_eco12589, w_eco12590, w_eco12591, w_eco12592, w_eco12593, w_eco12594, w_eco12595, w_eco12596, w_eco12597, w_eco12598, w_eco12599, w_eco12600, w_eco12601, w_eco12602, w_eco12603, w_eco12604, w_eco12605, w_eco12606, w_eco12607, w_eco12608, w_eco12609, w_eco12610, w_eco12611, w_eco12612, w_eco12613, w_eco12614, w_eco12615, w_eco12616, w_eco12617, w_eco12618, w_eco12619, w_eco12620, w_eco12621, w_eco12622, w_eco12623, w_eco12624, w_eco12625, w_eco12626, w_eco12627, w_eco12628, w_eco12629, w_eco12630, w_eco12631, w_eco12632, w_eco12633, w_eco12634, w_eco12635, w_eco12636, w_eco12637, w_eco12638, w_eco12639, w_eco12640, w_eco12641, w_eco12642, w_eco12643, w_eco12644, w_eco12645, w_eco12646, w_eco12647, w_eco12648, w_eco12649, w_eco12650, w_eco12651, w_eco12652, w_eco12653, w_eco12654, w_eco12655, w_eco12656, w_eco12657, w_eco12658, w_eco12659, w_eco12660, w_eco12661, w_eco12662, w_eco12663, w_eco12664, w_eco12665, w_eco12666, w_eco12667, w_eco12668, w_eco12669, w_eco12670, w_eco12671, w_eco12672, w_eco12673, w_eco12674, w_eco12675, w_eco12676, w_eco12677, w_eco12678, w_eco12679, w_eco12680, w_eco12681, w_eco12682, w_eco12683, w_eco12684, w_eco12685, w_eco12686, w_eco12687, w_eco12688, w_eco12689, w_eco12690, w_eco12691, w_eco12692, w_eco12693, w_eco12694, w_eco12695, w_eco12696, w_eco12697, w_eco12698, w_eco12699, w_eco12700, w_eco12701, w_eco12702, w_eco12703, w_eco12704, w_eco12705, w_eco12706, w_eco12707, w_eco12708, w_eco12709, w_eco12710, w_eco12711, w_eco12712, w_eco12713, w_eco12714, w_eco12715, w_eco12716, w_eco12717, w_eco12718, w_eco12719, w_eco12720, w_eco12721, w_eco12722, w_eco12723, w_eco12724, w_eco12725, w_eco12726, w_eco12727, w_eco12728, w_eco12729, w_eco12730, w_eco12731, w_eco12732, w_eco12733, w_eco12734, w_eco12735, w_eco12736, w_eco12737, w_eco12738, w_eco12739, w_eco12740, w_eco12741, w_eco12742, w_eco12743, w_eco12744, w_eco12745, w_eco12746, w_eco12747, w_eco12748, w_eco12749, w_eco12750, w_eco12751, w_eco12752, w_eco12753, w_eco12754, w_eco12755, w_eco12756, w_eco12757, w_eco12758, w_eco12759, w_eco12760, w_eco12761, w_eco12762, w_eco12763, w_eco12764, w_eco12765, w_eco12766, w_eco12767, w_eco12768, w_eco12769, w_eco12770, w_eco12771, w_eco12772, w_eco12773, w_eco12774, w_eco12775, w_eco12776, w_eco12777, w_eco12778, w_eco12779, w_eco12780, w_eco12781, w_eco12782, w_eco12783, w_eco12784, w_eco12785, w_eco12786, w_eco12787, w_eco12788, w_eco12789, w_eco12790, w_eco12791, w_eco12792, w_eco12793, w_eco12794, w_eco12795, w_eco12796, w_eco12797, w_eco12798, w_eco12799, w_eco12800, w_eco12801, w_eco12802, w_eco12803, w_eco12804, w_eco12805, w_eco12806, w_eco12807, w_eco12808, w_eco12809, w_eco12810, w_eco12811, w_eco12812, w_eco12813, w_eco12814, w_eco12815, w_eco12816, w_eco12817, w_eco12818, w_eco12819, w_eco12820, w_eco12821, w_eco12822, w_eco12823, w_eco12824, w_eco12825, w_eco12826, w_eco12827, w_eco12828, w_eco12829, w_eco12830, w_eco12831, w_eco12832, w_eco12833, w_eco12834, w_eco12835, w_eco12836, w_eco12837, w_eco12838, w_eco12839, w_eco12840, w_eco12841, w_eco12842, w_eco12843, w_eco12844, w_eco12845, w_eco12846, w_eco12847, w_eco12848, w_eco12849, w_eco12850, w_eco12851, w_eco12852, w_eco12853, w_eco12854, w_eco12855, w_eco12856, w_eco12857, w_eco12858, w_eco12859, w_eco12860, w_eco12861, w_eco12862, w_eco12863, w_eco12864, w_eco12865, w_eco12866, w_eco12867, w_eco12868, w_eco12869, w_eco12870, w_eco12871, w_eco12872, w_eco12873, w_eco12874, w_eco12875, w_eco12876, w_eco12877, w_eco12878, w_eco12879, w_eco12880, w_eco12881, w_eco12882, w_eco12883, w_eco12884, w_eco12885, w_eco12886, w_eco12887, w_eco12888, w_eco12889, w_eco12890, w_eco12891, w_eco12892, w_eco12893, w_eco12894, w_eco12895, w_eco12896, w_eco12897, w_eco12898, w_eco12899, w_eco12900, w_eco12901, w_eco12902, w_eco12903, w_eco12904, w_eco12905, w_eco12906, w_eco12907, w_eco12908, w_eco12909, w_eco12910, w_eco12911, w_eco12912, w_eco12913, w_eco12914, w_eco12915, w_eco12916, w_eco12917, w_eco12918, w_eco12919, w_eco12920, w_eco12921, w_eco12922, w_eco12923, w_eco12924, w_eco12925, w_eco12926, w_eco12927, w_eco12928, w_eco12929, w_eco12930, w_eco12931, w_eco12932, w_eco12933, w_eco12934, w_eco12935, w_eco12936, w_eco12937, w_eco12938, w_eco12939, w_eco12940, w_eco12941, w_eco12942, w_eco12943, w_eco12944, w_eco12945, w_eco12946, w_eco12947, w_eco12948, w_eco12949, w_eco12950, w_eco12951, w_eco12952, w_eco12953, w_eco12954, w_eco12955, w_eco12956, w_eco12957, w_eco12958, w_eco12959, w_eco12960, w_eco12961, w_eco12962, w_eco12963, w_eco12964, w_eco12965, w_eco12966, w_eco12967, w_eco12968, w_eco12969, w_eco12970, w_eco12971, w_eco12972, w_eco12973, w_eco12974, w_eco12975, w_eco12976, w_eco12977, w_eco12978, w_eco12979, w_eco12980, w_eco12981, w_eco12982, w_eco12983, w_eco12984, w_eco12985, w_eco12986, w_eco12987, w_eco12988, w_eco12989, w_eco12990, w_eco12991, w_eco12992, w_eco12993, w_eco12994, w_eco12995, w_eco12996, w_eco12997, w_eco12998, w_eco12999, w_eco13000, w_eco13001, w_eco13002, w_eco13003, w_eco13004, w_eco13005, w_eco13006, w_eco13007, w_eco13008, w_eco13009, w_eco13010, w_eco13011, w_eco13012, w_eco13013, w_eco13014, w_eco13015, w_eco13016, w_eco13017, w_eco13018, w_eco13019, w_eco13020, w_eco13021, w_eco13022, w_eco13023, w_eco13024, w_eco13025, w_eco13026, w_eco13027, w_eco13028, w_eco13029, w_eco13030, w_eco13031, w_eco13032, w_eco13033, w_eco13034, w_eco13035, w_eco13036, w_eco13037, w_eco13038, w_eco13039, w_eco13040, w_eco13041, w_eco13042, w_eco13043, w_eco13044, w_eco13045, w_eco13046, w_eco13047, w_eco13048, w_eco13049, w_eco13050, w_eco13051, w_eco13052, w_eco13053, w_eco13054, w_eco13055, w_eco13056, w_eco13057, w_eco13058, w_eco13059, w_eco13060, w_eco13061, w_eco13062, w_eco13063, w_eco13064, w_eco13065, w_eco13066, w_eco13067, w_eco13068, w_eco13069, w_eco13070, w_eco13071, w_eco13072, w_eco13073, w_eco13074, w_eco13075, w_eco13076, w_eco13077, w_eco13078, w_eco13079, w_eco13080, w_eco13081, w_eco13082, w_eco13083, w_eco13084, w_eco13085, w_eco13086, w_eco13087, w_eco13088, w_eco13089, w_eco13090, w_eco13091, w_eco13092, w_eco13093, w_eco13094, w_eco13095, w_eco13096, w_eco13097, w_eco13098, w_eco13099, w_eco13100, w_eco13101, w_eco13102, w_eco13103, w_eco13104, w_eco13105, w_eco13106, w_eco13107, w_eco13108, w_eco13109, w_eco13110, w_eco13111, w_eco13112, w_eco13113, w_eco13114, w_eco13115, w_eco13116, w_eco13117, w_eco13118, w_eco13119, w_eco13120, w_eco13121, w_eco13122, w_eco13123, w_eco13124, w_eco13125, w_eco13126, w_eco13127, w_eco13128, w_eco13129, w_eco13130, w_eco13131, w_eco13132, w_eco13133, w_eco13134, w_eco13135, w_eco13136, w_eco13137, w_eco13138, w_eco13139, w_eco13140, w_eco13141, w_eco13142, w_eco13143, w_eco13144, w_eco13145, w_eco13146, w_eco13147, w_eco13148, w_eco13149, w_eco13150, w_eco13151, w_eco13152, w_eco13153, w_eco13154, w_eco13155, w_eco13156, w_eco13157, w_eco13158, w_eco13159, w_eco13160, w_eco13161, w_eco13162, w_eco13163, w_eco13164, w_eco13165, w_eco13166, w_eco13167, w_eco13168, w_eco13169, w_eco13170, w_eco13171, w_eco13172, w_eco13173, w_eco13174, w_eco13175, w_eco13176, w_eco13177, w_eco13178, w_eco13179, w_eco13180, w_eco13181, w_eco13182, w_eco13183, w_eco13184, w_eco13185, w_eco13186, w_eco13187, w_eco13188, w_eco13189, w_eco13190, w_eco13191, w_eco13192, w_eco13193, w_eco13194, w_eco13195, w_eco13196, w_eco13197, w_eco13198, w_eco13199, w_eco13200, w_eco13201, w_eco13202, w_eco13203, w_eco13204, w_eco13205, w_eco13206, w_eco13207, w_eco13208, w_eco13209, w_eco13210, w_eco13211, w_eco13212, w_eco13213, w_eco13214, w_eco13215, w_eco13216, w_eco13217, w_eco13218, w_eco13219, w_eco13220, w_eco13221, w_eco13222, w_eco13223, w_eco13224, w_eco13225, w_eco13226, w_eco13227, w_eco13228, w_eco13229, w_eco13230, w_eco13231, w_eco13232, w_eco13233, w_eco13234, w_eco13235, w_eco13236, w_eco13237, w_eco13238, w_eco13239, w_eco13240, w_eco13241, w_eco13242, w_eco13243, w_eco13244, w_eco13245, w_eco13246, w_eco13247, w_eco13248, w_eco13249, w_eco13250, w_eco13251, w_eco13252, w_eco13253, w_eco13254, w_eco13255, w_eco13256, w_eco13257, w_eco13258, w_eco13259, w_eco13260, w_eco13261, w_eco13262, w_eco13263, w_eco13264, w_eco13265, w_eco13266, w_eco13267, w_eco13268, w_eco13269, w_eco13270, w_eco13271, w_eco13272, w_eco13273, w_eco13274, w_eco13275, w_eco13276, w_eco13277, w_eco13278, w_eco13279, w_eco13280, w_eco13281, w_eco13282, w_eco13283, w_eco13284, w_eco13285, w_eco13286, w_eco13287, w_eco13288, w_eco13289, w_eco13290, w_eco13291, w_eco13292, w_eco13293, w_eco13294, w_eco13295, w_eco13296, w_eco13297, w_eco13298, w_eco13299, w_eco13300, w_eco13301, w_eco13302, w_eco13303, w_eco13304, w_eco13305, w_eco13306, w_eco13307, w_eco13308, w_eco13309, w_eco13310, w_eco13311, w_eco13312, w_eco13313, w_eco13314, w_eco13315, w_eco13316, w_eco13317, w_eco13318, w_eco13319, w_eco13320, w_eco13321, w_eco13322, w_eco13323, w_eco13324, w_eco13325, w_eco13326, w_eco13327, w_eco13328, w_eco13329, w_eco13330, w_eco13331, w_eco13332, w_eco13333, w_eco13334, w_eco13335, w_eco13336, w_eco13337, w_eco13338, w_eco13339, w_eco13340, w_eco13341, w_eco13342, w_eco13343, w_eco13344, w_eco13345, w_eco13346, w_eco13347, w_eco13348, w_eco13349, w_eco13350, w_eco13351, w_eco13352, w_eco13353, w_eco13354, w_eco13355, w_eco13356, w_eco13357, w_eco13358, w_eco13359, w_eco13360, w_eco13361, w_eco13362, w_eco13363, w_eco13364, w_eco13365, w_eco13366, w_eco13367, w_eco13368, w_eco13369, w_eco13370, w_eco13371, w_eco13372, w_eco13373, w_eco13374, w_eco13375, w_eco13376, w_eco13377, w_eco13378, w_eco13379, w_eco13380, w_eco13381, w_eco13382, w_eco13383, w_eco13384, w_eco13385, w_eco13386, w_eco13387, w_eco13388, w_eco13389, w_eco13390, w_eco13391, w_eco13392, w_eco13393, w_eco13394, w_eco13395, w_eco13396, w_eco13397, w_eco13398, w_eco13399, w_eco13400, w_eco13401, w_eco13402, w_eco13403, w_eco13404, w_eco13405, w_eco13406, w_eco13407, w_eco13408, w_eco13409, w_eco13410, w_eco13411, w_eco13412, w_eco13413, w_eco13414, w_eco13415, w_eco13416, w_eco13417, w_eco13418, w_eco13419, w_eco13420, w_eco13421, w_eco13422, w_eco13423, w_eco13424, w_eco13425, w_eco13426, w_eco13427, w_eco13428, w_eco13429, w_eco13430, w_eco13431, w_eco13432, w_eco13433, w_eco13434, w_eco13435, w_eco13436, w_eco13437, w_eco13438, w_eco13439, w_eco13440, w_eco13441, w_eco13442, w_eco13443, w_eco13444, w_eco13445, w_eco13446, w_eco13447, w_eco13448, w_eco13449, w_eco13450, w_eco13451, w_eco13452, w_eco13453, w_eco13454, w_eco13455, w_eco13456, w_eco13457, w_eco13458, w_eco13459, w_eco13460, w_eco13461, w_eco13462, w_eco13463, w_eco13464, w_eco13465, w_eco13466, w_eco13467, w_eco13468, w_eco13469, w_eco13470, w_eco13471, w_eco13472, w_eco13473, w_eco13474, w_eco13475, w_eco13476, w_eco13477, w_eco13478, w_eco13479, w_eco13480, w_eco13481, w_eco13482, w_eco13483, w_eco13484, w_eco13485, w_eco13486, w_eco13487, w_eco13488, w_eco13489, w_eco13490, w_eco13491, w_eco13492, w_eco13493, w_eco13494, w_eco13495, w_eco13496, w_eco13497, w_eco13498, w_eco13499, w_eco13500, w_eco13501, w_eco13502, w_eco13503, w_eco13504, w_eco13505, w_eco13506, w_eco13507, w_eco13508, w_eco13509, w_eco13510, w_eco13511, w_eco13512, w_eco13513, w_eco13514, w_eco13515, w_eco13516, w_eco13517, w_eco13518, w_eco13519, w_eco13520, w_eco13521, w_eco13522, w_eco13523, w_eco13524, w_eco13525, w_eco13526, w_eco13527, w_eco13528, w_eco13529, w_eco13530, w_eco13531, w_eco13532, w_eco13533, w_eco13534, w_eco13535, w_eco13536, w_eco13537, w_eco13538, w_eco13539, w_eco13540, w_eco13541, w_eco13542, w_eco13543, w_eco13544, w_eco13545, w_eco13546, w_eco13547, w_eco13548, w_eco13549, w_eco13550, w_eco13551, w_eco13552, w_eco13553, w_eco13554, w_eco13555, w_eco13556, w_eco13557, w_eco13558, w_eco13559, w_eco13560, w_eco13561, w_eco13562, w_eco13563, w_eco13564, w_eco13565, w_eco13566, w_eco13567, w_eco13568, w_eco13569, w_eco13570, w_eco13571, w_eco13572, w_eco13573, w_eco13574, w_eco13575, w_eco13576, w_eco13577, w_eco13578, w_eco13579, w_eco13580, w_eco13581, w_eco13582, w_eco13583, w_eco13584, w_eco13585, w_eco13586, w_eco13587, w_eco13588, w_eco13589, w_eco13590, w_eco13591, w_eco13592, w_eco13593, w_eco13594, w_eco13595, w_eco13596, w_eco13597, w_eco13598, w_eco13599, w_eco13600, w_eco13601, w_eco13602, w_eco13603, w_eco13604, w_eco13605, w_eco13606, w_eco13607, w_eco13608, w_eco13609, w_eco13610, w_eco13611, w_eco13612, w_eco13613, w_eco13614, w_eco13615, w_eco13616, w_eco13617, w_eco13618, w_eco13619, w_eco13620, w_eco13621, w_eco13622, w_eco13623, w_eco13624, w_eco13625, w_eco13626, w_eco13627, w_eco13628, w_eco13629, w_eco13630, w_eco13631, w_eco13632, w_eco13633, w_eco13634, w_eco13635, w_eco13636, w_eco13637, w_eco13638, w_eco13639, w_eco13640, w_eco13641, w_eco13642, w_eco13643, w_eco13644, w_eco13645, w_eco13646, w_eco13647, w_eco13648, w_eco13649, w_eco13650, w_eco13651, w_eco13652, w_eco13653, w_eco13654, w_eco13655, w_eco13656, w_eco13657, w_eco13658, w_eco13659, w_eco13660, w_eco13661, w_eco13662, w_eco13663, w_eco13664, w_eco13665, w_eco13666, w_eco13667, w_eco13668, w_eco13669, w_eco13670, w_eco13671, w_eco13672, w_eco13673, w_eco13674, w_eco13675, w_eco13676, w_eco13677, w_eco13678, w_eco13679, w_eco13680, w_eco13681, w_eco13682, w_eco13683, w_eco13684, w_eco13685, w_eco13686, w_eco13687, w_eco13688, w_eco13689, w_eco13690, w_eco13691, w_eco13692, w_eco13693, w_eco13694, w_eco13695, w_eco13696, w_eco13697, w_eco13698, w_eco13699, w_eco13700, w_eco13701, w_eco13702, w_eco13703, w_eco13704, w_eco13705, w_eco13706, w_eco13707, w_eco13708, w_eco13709, w_eco13710, w_eco13711, w_eco13712, w_eco13713, w_eco13714, w_eco13715, w_eco13716, w_eco13717, w_eco13718, w_eco13719, w_eco13720, w_eco13721, w_eco13722, w_eco13723, w_eco13724, w_eco13725, w_eco13726, w_eco13727, w_eco13728, w_eco13729, w_eco13730, w_eco13731, w_eco13732, w_eco13733, w_eco13734, w_eco13735, w_eco13736, w_eco13737, w_eco13738, w_eco13739, w_eco13740, w_eco13741, w_eco13742, w_eco13743, w_eco13744, w_eco13745, w_eco13746, w_eco13747, w_eco13748, w_eco13749, w_eco13750, w_eco13751, w_eco13752, w_eco13753, w_eco13754, w_eco13755, w_eco13756, w_eco13757, w_eco13758, w_eco13759, w_eco13760, w_eco13761, w_eco13762, w_eco13763, w_eco13764, w_eco13765, w_eco13766, w_eco13767, w_eco13768, w_eco13769, w_eco13770, w_eco13771, w_eco13772, w_eco13773, w_eco13774, w_eco13775, w_eco13776, w_eco13777, w_eco13778, w_eco13779, w_eco13780, w_eco13781, w_eco13782, w_eco13783, w_eco13784, w_eco13785, w_eco13786, w_eco13787, w_eco13788, w_eco13789, w_eco13790, w_eco13791, w_eco13792, w_eco13793, w_eco13794, w_eco13795, w_eco13796, w_eco13797, w_eco13798, w_eco13799, w_eco13800, w_eco13801, w_eco13802, w_eco13803, w_eco13804, w_eco13805, w_eco13806, w_eco13807, w_eco13808, w_eco13809, w_eco13810, w_eco13811, w_eco13812, w_eco13813, w_eco13814, w_eco13815, w_eco13816, w_eco13817, w_eco13818, w_eco13819, w_eco13820, w_eco13821, w_eco13822, w_eco13823, w_eco13824, w_eco13825, w_eco13826, w_eco13827, w_eco13828, w_eco13829, w_eco13830, w_eco13831, w_eco13832, w_eco13833, w_eco13834, w_eco13835, w_eco13836, w_eco13837, w_eco13838, w_eco13839, w_eco13840, w_eco13841, w_eco13842, w_eco13843, w_eco13844, w_eco13845, w_eco13846, w_eco13847, w_eco13848, w_eco13849, w_eco13850, w_eco13851, w_eco13852, w_eco13853, w_eco13854, w_eco13855, w_eco13856, w_eco13857, w_eco13858, w_eco13859, w_eco13860, w_eco13861, w_eco13862, w_eco13863, w_eco13864, w_eco13865, w_eco13866, w_eco13867, w_eco13868, w_eco13869, w_eco13870, w_eco13871, w_eco13872, w_eco13873, w_eco13874, w_eco13875, w_eco13876, w_eco13877, w_eco13878, w_eco13879, w_eco13880, w_eco13881, w_eco13882, w_eco13883, w_eco13884, w_eco13885, w_eco13886, w_eco13887, w_eco13888, w_eco13889, w_eco13890, w_eco13891, w_eco13892, w_eco13893, w_eco13894, w_eco13895, w_eco13896, w_eco13897, w_eco13898, w_eco13899, w_eco13900, w_eco13901, w_eco13902, w_eco13903, w_eco13904, w_eco13905, w_eco13906, w_eco13907, w_eco13908, w_eco13909, w_eco13910, w_eco13911, w_eco13912, w_eco13913, w_eco13914, w_eco13915, w_eco13916, w_eco13917, w_eco13918, w_eco13919, w_eco13920, w_eco13921, w_eco13922, w_eco13923, w_eco13924, w_eco13925, w_eco13926, w_eco13927, w_eco13928, w_eco13929, w_eco13930, w_eco13931, w_eco13932, w_eco13933, w_eco13934, w_eco13935, w_eco13936, w_eco13937, w_eco13938, w_eco13939, w_eco13940, w_eco13941, w_eco13942, w_eco13943, w_eco13944, w_eco13945, w_eco13946, w_eco13947, w_eco13948, w_eco13949, w_eco13950, w_eco13951, w_eco13952, w_eco13953, w_eco13954, w_eco13955, w_eco13956, w_eco13957, w_eco13958, w_eco13959, w_eco13960, w_eco13961, w_eco13962, w_eco13963, w_eco13964, w_eco13965, w_eco13966, w_eco13967, w_eco13968, w_eco13969, w_eco13970, w_eco13971, w_eco13972, w_eco13973, w_eco13974, w_eco13975, w_eco13976, w_eco13977, w_eco13978, w_eco13979, w_eco13980, w_eco13981, w_eco13982, w_eco13983, w_eco13984, w_eco13985, w_eco13986, w_eco13987, w_eco13988, w_eco13989, w_eco13990, w_eco13991, w_eco13992, w_eco13993, w_eco13994, w_eco13995, w_eco13996, w_eco13997, w_eco13998, w_eco13999, w_eco14000, w_eco14001, w_eco14002, w_eco14003, w_eco14004, w_eco14005, w_eco14006, w_eco14007, w_eco14008, w_eco14009, w_eco14010, w_eco14011, w_eco14012, w_eco14013, w_eco14014, w_eco14015, w_eco14016, w_eco14017, w_eco14018, w_eco14019, w_eco14020, w_eco14021, w_eco14022, w_eco14023, w_eco14024, w_eco14025, w_eco14026, w_eco14027, w_eco14028, w_eco14029, w_eco14030, w_eco14031, w_eco14032, w_eco14033, w_eco14034, w_eco14035, w_eco14036, w_eco14037, w_eco14038, w_eco14039, w_eco14040, w_eco14041, w_eco14042, w_eco14043, w_eco14044, w_eco14045, w_eco14046, w_eco14047, w_eco14048, w_eco14049, w_eco14050, w_eco14051, w_eco14052, w_eco14053, w_eco14054, w_eco14055, w_eco14056, w_eco14057, w_eco14058, w_eco14059, w_eco14060, w_eco14061, w_eco14062, w_eco14063, w_eco14064, w_eco14065, w_eco14066, w_eco14067, w_eco14068, w_eco14069, w_eco14070, w_eco14071, w_eco14072, w_eco14073, w_eco14074, w_eco14075, w_eco14076, w_eco14077, w_eco14078, w_eco14079, w_eco14080, w_eco14081, w_eco14082, w_eco14083, w_eco14084, w_eco14085, w_eco14086, w_eco14087, w_eco14088, w_eco14089, w_eco14090, w_eco14091, w_eco14092, w_eco14093, w_eco14094, w_eco14095, w_eco14096, w_eco14097, w_eco14098, w_eco14099, w_eco14100, w_eco14101, w_eco14102, w_eco14103, w_eco14104, w_eco14105, w_eco14106, w_eco14107, w_eco14108, w_eco14109, w_eco14110, w_eco14111, w_eco14112, w_eco14113, w_eco14114, w_eco14115, w_eco14116, w_eco14117, w_eco14118, w_eco14119, w_eco14120, w_eco14121, w_eco14122, w_eco14123, w_eco14124, w_eco14125, w_eco14126, w_eco14127, w_eco14128, w_eco14129, w_eco14130, w_eco14131, w_eco14132, w_eco14133, w_eco14134, w_eco14135, w_eco14136, w_eco14137, w_eco14138, w_eco14139, w_eco14140, w_eco14141, w_eco14142, w_eco14143, w_eco14144, w_eco14145, w_eco14146, w_eco14147, w_eco14148, w_eco14149, w_eco14150, w_eco14151, w_eco14152, w_eco14153, w_eco14154, w_eco14155, w_eco14156, w_eco14157, w_eco14158, w_eco14159, w_eco14160, w_eco14161, w_eco14162, w_eco14163, w_eco14164, w_eco14165, w_eco14166, w_eco14167, w_eco14168, w_eco14169, w_eco14170, w_eco14171, w_eco14172, w_eco14173, w_eco14174, w_eco14175, w_eco14176, w_eco14177, w_eco14178, w_eco14179, w_eco14180, w_eco14181, w_eco14182, w_eco14183, w_eco14184, w_eco14185, w_eco14186, w_eco14187, w_eco14188, w_eco14189, w_eco14190, w_eco14191, w_eco14192, w_eco14193, w_eco14194, w_eco14195, w_eco14196, w_eco14197, w_eco14198, w_eco14199, w_eco14200, w_eco14201, w_eco14202, w_eco14203, w_eco14204, w_eco14205, w_eco14206, w_eco14207, w_eco14208, w_eco14209, w_eco14210, w_eco14211, w_eco14212, w_eco14213, w_eco14214, w_eco14215, w_eco14216, w_eco14217, w_eco14218, w_eco14219, w_eco14220, w_eco14221, w_eco14222, w_eco14223, w_eco14224, w_eco14225, w_eco14226, w_eco14227, w_eco14228, w_eco14229, w_eco14230, w_eco14231, w_eco14232, w_eco14233, w_eco14234, w_eco14235, w_eco14236, w_eco14237, w_eco14238, w_eco14239, w_eco14240, w_eco14241, w_eco14242, w_eco14243, w_eco14244, w_eco14245, w_eco14246, w_eco14247, w_eco14248, w_eco14249, w_eco14250, w_eco14251, w_eco14252, w_eco14253, w_eco14254, w_eco14255, w_eco14256, w_eco14257, w_eco14258, w_eco14259, w_eco14260, w_eco14261, w_eco14262, w_eco14263, w_eco14264, w_eco14265, w_eco14266, w_eco14267, w_eco14268, w_eco14269, w_eco14270, w_eco14271, w_eco14272, w_eco14273, w_eco14274, w_eco14275, w_eco14276, w_eco14277, w_eco14278, w_eco14279, w_eco14280, w_eco14281, w_eco14282, w_eco14283, w_eco14284, w_eco14285, w_eco14286, w_eco14287, w_eco14288, w_eco14289, w_eco14290, w_eco14291, w_eco14292, w_eco14293, w_eco14294, w_eco14295, w_eco14296, w_eco14297, w_eco14298, w_eco14299, w_eco14300, w_eco14301, w_eco14302, w_eco14303, w_eco14304, w_eco14305, w_eco14306, w_eco14307, w_eco14308, w_eco14309, w_eco14310, w_eco14311, w_eco14312, w_eco14313, w_eco14314, w_eco14315, w_eco14316, w_eco14317, w_eco14318, w_eco14319, w_eco14320, w_eco14321, w_eco14322, w_eco14323, w_eco14324, w_eco14325, w_eco14326, w_eco14327, w_eco14328, w_eco14329, w_eco14330, w_eco14331, w_eco14332, w_eco14333, w_eco14334, w_eco14335, w_eco14336, w_eco14337, w_eco14338, w_eco14339, w_eco14340, w_eco14341, w_eco14342, w_eco14343, w_eco14344, w_eco14345, w_eco14346, w_eco14347, w_eco14348, w_eco14349, w_eco14350, w_eco14351, w_eco14352, w_eco14353, w_eco14354, w_eco14355, w_eco14356, w_eco14357, w_eco14358, w_eco14359, w_eco14360, w_eco14361, w_eco14362, w_eco14363, w_eco14364, w_eco14365, w_eco14366, w_eco14367, w_eco14368, w_eco14369, w_eco14370, w_eco14371, w_eco14372, w_eco14373, w_eco14374, w_eco14375, w_eco14376, w_eco14377, w_eco14378, w_eco14379, w_eco14380, w_eco14381, w_eco14382, w_eco14383, w_eco14384, w_eco14385, w_eco14386, w_eco14387, w_eco14388, w_eco14389, w_eco14390, w_eco14391, w_eco14392, w_eco14393, w_eco14394, w_eco14395, w_eco14396, w_eco14397, w_eco14398, w_eco14399, w_eco14400, w_eco14401, w_eco14402, w_eco14403, w_eco14404, w_eco14405, w_eco14406, w_eco14407, w_eco14408, w_eco14409, w_eco14410, w_eco14411, w_eco14412, w_eco14413, w_eco14414, w_eco14415, w_eco14416, w_eco14417, w_eco14418, w_eco14419, w_eco14420, w_eco14421, w_eco14422, w_eco14423, w_eco14424, w_eco14425, w_eco14426, w_eco14427, w_eco14428, w_eco14429, w_eco14430, w_eco14431, w_eco14432, w_eco14433, w_eco14434, w_eco14435, w_eco14436, w_eco14437, w_eco14438, w_eco14439, w_eco14440, w_eco14441, w_eco14442, w_eco14443, w_eco14444, w_eco14445, w_eco14446, w_eco14447, w_eco14448, w_eco14449, w_eco14450, w_eco14451, w_eco14452, w_eco14453, w_eco14454, w_eco14455, w_eco14456, w_eco14457, w_eco14458, w_eco14459, w_eco14460, w_eco14461, w_eco14462, w_eco14463, w_eco14464, w_eco14465, w_eco14466, w_eco14467, w_eco14468, w_eco14469, w_eco14470, w_eco14471, w_eco14472, w_eco14473, w_eco14474, w_eco14475, w_eco14476, w_eco14477, w_eco14478, w_eco14479, w_eco14480, w_eco14481, w_eco14482, w_eco14483, w_eco14484, w_eco14485, w_eco14486, w_eco14487, w_eco14488, w_eco14489, w_eco14490, w_eco14491, w_eco14492, w_eco14493, w_eco14494, w_eco14495, w_eco14496, w_eco14497, w_eco14498, w_eco14499, w_eco14500, w_eco14501, w_eco14502, w_eco14503, w_eco14504, w_eco14505, w_eco14506, w_eco14507, w_eco14508, w_eco14509, w_eco14510, w_eco14511, w_eco14512, w_eco14513, w_eco14514, w_eco14515, w_eco14516, w_eco14517, w_eco14518, w_eco14519, w_eco14520, w_eco14521, w_eco14522, w_eco14523, w_eco14524, w_eco14525, w_eco14526, w_eco14527, w_eco14528, w_eco14529, w_eco14530, w_eco14531, w_eco14532, w_eco14533, w_eco14534, w_eco14535, w_eco14536, w_eco14537, w_eco14538, w_eco14539, w_eco14540, w_eco14541, w_eco14542, w_eco14543, w_eco14544, w_eco14545, w_eco14546, w_eco14547, w_eco14548, w_eco14549, w_eco14550, w_eco14551, w_eco14552, w_eco14553, w_eco14554, w_eco14555, w_eco14556, w_eco14557, w_eco14558, w_eco14559, w_eco14560, w_eco14561, w_eco14562, w_eco14563, w_eco14564, w_eco14565, w_eco14566, w_eco14567, w_eco14568, w_eco14569, w_eco14570, w_eco14571, w_eco14572, w_eco14573, w_eco14574, w_eco14575, w_eco14576, w_eco14577, w_eco14578, w_eco14579, w_eco14580, w_eco14581, w_eco14582, w_eco14583, w_eco14584, w_eco14585, w_eco14586, w_eco14587, w_eco14588, w_eco14589, w_eco14590, w_eco14591, w_eco14592, w_eco14593, w_eco14594, w_eco14595, w_eco14596, w_eco14597, w_eco14598, w_eco14599, w_eco14600, w_eco14601, w_eco14602, w_eco14603, w_eco14604, w_eco14605, w_eco14606, w_eco14607, w_eco14608, w_eco14609, w_eco14610, w_eco14611, w_eco14612, w_eco14613, w_eco14614, w_eco14615, w_eco14616, w_eco14617, w_eco14618, w_eco14619, w_eco14620, w_eco14621, w_eco14622, w_eco14623, w_eco14624, w_eco14625, w_eco14626, w_eco14627, w_eco14628, w_eco14629, w_eco14630, w_eco14631, w_eco14632, w_eco14633, w_eco14634, w_eco14635, w_eco14636, w_eco14637, w_eco14638, w_eco14639, w_eco14640, w_eco14641, w_eco14642, w_eco14643, w_eco14644, w_eco14645, w_eco14646, w_eco14647, w_eco14648, w_eco14649, w_eco14650, w_eco14651, w_eco14652, w_eco14653, w_eco14654, w_eco14655, w_eco14656, w_eco14657, w_eco14658, w_eco14659, w_eco14660, w_eco14661, w_eco14662, w_eco14663, w_eco14664, w_eco14665, w_eco14666, w_eco14667, w_eco14668, w_eco14669, w_eco14670, w_eco14671, w_eco14672, w_eco14673, w_eco14674, w_eco14675, w_eco14676, w_eco14677, w_eco14678, w_eco14679, w_eco14680, w_eco14681, w_eco14682, w_eco14683, w_eco14684, w_eco14685, w_eco14686, w_eco14687, w_eco14688, w_eco14689, w_eco14690, w_eco14691, w_eco14692, w_eco14693, w_eco14694, w_eco14695, w_eco14696, w_eco14697, w_eco14698, w_eco14699, w_eco14700, w_eco14701, w_eco14702, w_eco14703, w_eco14704, w_eco14705, w_eco14706, w_eco14707, w_eco14708, w_eco14709, w_eco14710, w_eco14711, w_eco14712, w_eco14713, w_eco14714, w_eco14715, w_eco14716, w_eco14717, w_eco14718, w_eco14719, w_eco14720, w_eco14721, w_eco14722, w_eco14723, w_eco14724, w_eco14725, w_eco14726, w_eco14727, w_eco14728, w_eco14729, w_eco14730, w_eco14731, w_eco14732, w_eco14733, w_eco14734, w_eco14735, w_eco14736, w_eco14737, w_eco14738, w_eco14739, w_eco14740, w_eco14741, w_eco14742, w_eco14743, w_eco14744, w_eco14745, w_eco14746, w_eco14747, w_eco14748, w_eco14749, w_eco14750, w_eco14751, w_eco14752, w_eco14753, w_eco14754, w_eco14755, w_eco14756, w_eco14757, w_eco14758, w_eco14759, w_eco14760, w_eco14761, w_eco14762, w_eco14763, w_eco14764, w_eco14765, w_eco14766, w_eco14767, w_eco14768, w_eco14769, w_eco14770, w_eco14771, w_eco14772, w_eco14773, w_eco14774, w_eco14775, w_eco14776, w_eco14777, w_eco14778, w_eco14779, w_eco14780, w_eco14781, w_eco14782, w_eco14783, w_eco14784, w_eco14785, w_eco14786, w_eco14787, w_eco14788, w_eco14789, w_eco14790, w_eco14791, w_eco14792, w_eco14793, w_eco14794, w_eco14795, w_eco14796, w_eco14797, w_eco14798, w_eco14799, w_eco14800, w_eco14801, w_eco14802, w_eco14803, w_eco14804, w_eco14805, w_eco14806, w_eco14807, w_eco14808, w_eco14809, w_eco14810, w_eco14811, w_eco14812, w_eco14813, w_eco14814, w_eco14815, w_eco14816, w_eco14817, w_eco14818, w_eco14819, w_eco14820, w_eco14821, w_eco14822, w_eco14823, w_eco14824, w_eco14825, w_eco14826, w_eco14827, w_eco14828, w_eco14829, w_eco14830, w_eco14831, w_eco14832, w_eco14833, w_eco14834, w_eco14835, w_eco14836, w_eco14837, w_eco14838, w_eco14839, w_eco14840, w_eco14841, w_eco14842, w_eco14843, w_eco14844, w_eco14845, w_eco14846, w_eco14847, w_eco14848, w_eco14849, w_eco14850, w_eco14851, w_eco14852, w_eco14853, w_eco14854, w_eco14855, w_eco14856, w_eco14857, w_eco14858, w_eco14859, w_eco14860, w_eco14861, w_eco14862, w_eco14863, w_eco14864, w_eco14865, w_eco14866, w_eco14867, w_eco14868, w_eco14869, w_eco14870, w_eco14871, w_eco14872, w_eco14873, w_eco14874, w_eco14875, w_eco14876, w_eco14877, w_eco14878, w_eco14879, w_eco14880, w_eco14881, w_eco14882, w_eco14883, w_eco14884, w_eco14885, w_eco14886, w_eco14887, w_eco14888, w_eco14889, w_eco14890, w_eco14891, w_eco14892, w_eco14893, w_eco14894, w_eco14895, w_eco14896, w_eco14897, w_eco14898, w_eco14899, w_eco14900, w_eco14901, w_eco14902, w_eco14903, w_eco14904, w_eco14905, w_eco14906, w_eco14907, w_eco14908, w_eco14909, w_eco14910, w_eco14911, w_eco14912, w_eco14913, w_eco14914, w_eco14915, w_eco14916, w_eco14917, w_eco14918, w_eco14919, w_eco14920, w_eco14921, w_eco14922, w_eco14923, w_eco14924, w_eco14925, w_eco14926, w_eco14927, w_eco14928, w_eco14929, w_eco14930, w_eco14931, w_eco14932, w_eco14933, w_eco14934, w_eco14935, w_eco14936, w_eco14937, w_eco14938, w_eco14939, w_eco14940, w_eco14941, w_eco14942, w_eco14943, w_eco14944, w_eco14945, w_eco14946, w_eco14947, w_eco14948, w_eco14949, w_eco14950, w_eco14951, w_eco14952, w_eco14953, w_eco14954, w_eco14955, w_eco14956, w_eco14957, w_eco14958, w_eco14959, w_eco14960, w_eco14961, w_eco14962, w_eco14963, w_eco14964, w_eco14965, w_eco14966, w_eco14967, w_eco14968, w_eco14969, w_eco14970, w_eco14971, w_eco14972, w_eco14973, w_eco14974, w_eco14975, w_eco14976, w_eco14977, w_eco14978, w_eco14979, w_eco14980, w_eco14981, w_eco14982, w_eco14983, w_eco14984, w_eco14985, w_eco14986, w_eco14987, w_eco14988, w_eco14989, w_eco14990, w_eco14991, w_eco14992, w_eco14993, w_eco14994, w_eco14995, w_eco14996, w_eco14997, w_eco14998, w_eco14999, w_eco15000, w_eco15001, w_eco15002, w_eco15003, w_eco15004, w_eco15005, w_eco15006, w_eco15007, w_eco15008, w_eco15009, w_eco15010, w_eco15011, w_eco15012, w_eco15013, w_eco15014, w_eco15015, w_eco15016, w_eco15017, w_eco15018, w_eco15019, w_eco15020, w_eco15021, w_eco15022, w_eco15023, w_eco15024, w_eco15025, w_eco15026, w_eco15027, w_eco15028, w_eco15029, w_eco15030, w_eco15031, w_eco15032, w_eco15033, w_eco15034, w_eco15035, w_eco15036, w_eco15037, w_eco15038, w_eco15039, w_eco15040, w_eco15041, w_eco15042, w_eco15043, w_eco15044, w_eco15045, w_eco15046, w_eco15047, w_eco15048, w_eco15049, w_eco15050, w_eco15051, w_eco15052, w_eco15053, w_eco15054, w_eco15055, w_eco15056, w_eco15057, w_eco15058, w_eco15059, w_eco15060, w_eco15061, w_eco15062, w_eco15063, w_eco15064, w_eco15065, w_eco15066, w_eco15067, w_eco15068, w_eco15069, w_eco15070, w_eco15071, w_eco15072, w_eco15073, w_eco15074, w_eco15075, w_eco15076, w_eco15077, w_eco15078, w_eco15079, w_eco15080, w_eco15081, w_eco15082, w_eco15083, w_eco15084, w_eco15085, w_eco15086, w_eco15087, w_eco15088, w_eco15089, w_eco15090, w_eco15091, w_eco15092, w_eco15093, w_eco15094, w_eco15095, w_eco15096, w_eco15097, w_eco15098, w_eco15099, w_eco15100, w_eco15101, w_eco15102, w_eco15103, w_eco15104, w_eco15105, w_eco15106, w_eco15107, w_eco15108, w_eco15109, w_eco15110, w_eco15111, w_eco15112, w_eco15113, w_eco15114, w_eco15115, w_eco15116, w_eco15117, w_eco15118, w_eco15119, w_eco15120, w_eco15121, w_eco15122, w_eco15123, w_eco15124, w_eco15125, w_eco15126, w_eco15127, w_eco15128, w_eco15129, w_eco15130, w_eco15131, w_eco15132, w_eco15133, w_eco15134, w_eco15135, w_eco15136, w_eco15137, w_eco15138, w_eco15139, w_eco15140, w_eco15141, w_eco15142, w_eco15143, w_eco15144, w_eco15145, w_eco15146, w_eco15147, w_eco15148, w_eco15149, w_eco15150, w_eco15151, w_eco15152, w_eco15153, w_eco15154, w_eco15155, w_eco15156, w_eco15157, w_eco15158, w_eco15159, w_eco15160, w_eco15161, w_eco15162, w_eco15163, w_eco15164, w_eco15165, w_eco15166, w_eco15167, w_eco15168, w_eco15169, w_eco15170, w_eco15171, w_eco15172, w_eco15173, w_eco15174, w_eco15175, w_eco15176, w_eco15177, w_eco15178, w_eco15179, w_eco15180, w_eco15181, w_eco15182, w_eco15183, w_eco15184, w_eco15185, w_eco15186, w_eco15187, w_eco15188, w_eco15189, w_eco15190, w_eco15191, w_eco15192, w_eco15193, w_eco15194, w_eco15195, w_eco15196, w_eco15197, w_eco15198, w_eco15199, w_eco15200, w_eco15201, w_eco15202, w_eco15203, w_eco15204, w_eco15205, w_eco15206, w_eco15207, w_eco15208, w_eco15209, w_eco15210, w_eco15211, w_eco15212, w_eco15213, w_eco15214, w_eco15215, w_eco15216, w_eco15217, w_eco15218, w_eco15219, w_eco15220, w_eco15221, w_eco15222, w_eco15223, w_eco15224, w_eco15225, w_eco15226, w_eco15227, w_eco15228, w_eco15229, w_eco15230, w_eco15231, w_eco15232, w_eco15233, w_eco15234, w_eco15235, w_eco15236, w_eco15237, w_eco15238, w_eco15239, w_eco15240, w_eco15241, w_eco15242, w_eco15243, w_eco15244, w_eco15245, w_eco15246, w_eco15247, w_eco15248, w_eco15249, w_eco15250, w_eco15251, w_eco15252, w_eco15253, w_eco15254, w_eco15255, w_eco15256, w_eco15257, w_eco15258, w_eco15259, w_eco15260, w_eco15261, w_eco15262, w_eco15263, w_eco15264, w_eco15265, w_eco15266, w_eco15267, w_eco15268, w_eco15269, w_eco15270, w_eco15271, w_eco15272, w_eco15273, w_eco15274, w_eco15275, w_eco15276, w_eco15277, w_eco15278, w_eco15279, w_eco15280, w_eco15281, w_eco15282, w_eco15283, w_eco15284, w_eco15285, w_eco15286, w_eco15287, w_eco15288, w_eco15289, w_eco15290, w_eco15291, w_eco15292, w_eco15293, w_eco15294, w_eco15295, w_eco15296, w_eco15297, w_eco15298, w_eco15299, w_eco15300, w_eco15301, w_eco15302, w_eco15303, w_eco15304, w_eco15305, w_eco15306, w_eco15307, w_eco15308, w_eco15309, w_eco15310, w_eco15311, w_eco15312, w_eco15313, w_eco15314, w_eco15315, w_eco15316, w_eco15317, w_eco15318, w_eco15319, w_eco15320, w_eco15321, w_eco15322, w_eco15323, w_eco15324, w_eco15325, w_eco15326, w_eco15327, w_eco15328, w_eco15329, w_eco15330, w_eco15331, w_eco15332, w_eco15333, w_eco15334, w_eco15335, w_eco15336, w_eco15337, w_eco15338, w_eco15339, w_eco15340, w_eco15341, w_eco15342, w_eco15343, w_eco15344, w_eco15345, w_eco15346, w_eco15347, w_eco15348, w_eco15349, w_eco15350, w_eco15351, w_eco15352, w_eco15353, w_eco15354, w_eco15355, w_eco15356, w_eco15357, w_eco15358, w_eco15359, w_eco15360, w_eco15361, w_eco15362, w_eco15363, w_eco15364, w_eco15365, w_eco15366, w_eco15367, w_eco15368, w_eco15369, w_eco15370, w_eco15371, w_eco15372, w_eco15373, w_eco15374, w_eco15375, w_eco15376, w_eco15377, w_eco15378, w_eco15379, w_eco15380, w_eco15381, w_eco15382, w_eco15383, w_eco15384, w_eco15385, w_eco15386, w_eco15387, w_eco15388, w_eco15389, w_eco15390, w_eco15391, w_eco15392, w_eco15393, w_eco15394, w_eco15395, w_eco15396, w_eco15397, w_eco15398, w_eco15399, w_eco15400, w_eco15401, w_eco15402, w_eco15403, w_eco15404, w_eco15405, w_eco15406, w_eco15407, w_eco15408, w_eco15409, w_eco15410, w_eco15411, w_eco15412, w_eco15413, w_eco15414, w_eco15415, w_eco15416, w_eco15417, w_eco15418, w_eco15419, w_eco15420, w_eco15421, w_eco15422, w_eco15423, w_eco15424, w_eco15425, w_eco15426, w_eco15427, w_eco15428, w_eco15429, w_eco15430, w_eco15431, w_eco15432, w_eco15433, w_eco15434, w_eco15435, w_eco15436, w_eco15437, w_eco15438, w_eco15439, w_eco15440, w_eco15441, w_eco15442, w_eco15443, w_eco15444, w_eco15445, w_eco15446, w_eco15447, w_eco15448, w_eco15449, w_eco15450, w_eco15451, w_eco15452, w_eco15453, w_eco15454, w_eco15455, w_eco15456, w_eco15457, w_eco15458, w_eco15459, w_eco15460, w_eco15461, w_eco15462, w_eco15463, w_eco15464, w_eco15465, w_eco15466, w_eco15467, w_eco15468, w_eco15469, w_eco15470, w_eco15471, w_eco15472, w_eco15473, w_eco15474, w_eco15475, w_eco15476, w_eco15477, w_eco15478, w_eco15479, w_eco15480, w_eco15481, w_eco15482, w_eco15483, w_eco15484, w_eco15485, w_eco15486, w_eco15487, w_eco15488, w_eco15489, w_eco15490, w_eco15491, w_eco15492, w_eco15493, w_eco15494, w_eco15495, w_eco15496, w_eco15497, w_eco15498, w_eco15499, w_eco15500, w_eco15501, w_eco15502, w_eco15503, w_eco15504, w_eco15505, w_eco15506, w_eco15507, w_eco15508, w_eco15509, w_eco15510, w_eco15511, w_eco15512, w_eco15513, w_eco15514, w_eco15515, w_eco15516, w_eco15517, w_eco15518, w_eco15519, w_eco15520, w_eco15521, w_eco15522, w_eco15523, w_eco15524, w_eco15525, w_eco15526, w_eco15527, w_eco15528, w_eco15529, w_eco15530, w_eco15531, w_eco15532, w_eco15533, w_eco15534, w_eco15535, w_eco15536, w_eco15537, w_eco15538, w_eco15539, w_eco15540, w_eco15541, w_eco15542, w_eco15543, w_eco15544, w_eco15545, w_eco15546, w_eco15547, w_eco15548, w_eco15549, w_eco15550, w_eco15551, w_eco15552, w_eco15553, w_eco15554, w_eco15555, w_eco15556, w_eco15557, w_eco15558, w_eco15559, w_eco15560, w_eco15561, w_eco15562, w_eco15563, w_eco15564, w_eco15565, w_eco15566, w_eco15567, w_eco15568, w_eco15569, w_eco15570, w_eco15571, w_eco15572, w_eco15573, w_eco15574, w_eco15575, w_eco15576, w_eco15577, w_eco15578, w_eco15579, w_eco15580, w_eco15581, w_eco15582, w_eco15583, w_eco15584, w_eco15585, w_eco15586, w_eco15587, w_eco15588, w_eco15589, w_eco15590, w_eco15591, w_eco15592, w_eco15593, w_eco15594, w_eco15595, w_eco15596, w_eco15597, w_eco15598, w_eco15599, w_eco15600, w_eco15601, w_eco15602, w_eco15603, w_eco15604, w_eco15605, w_eco15606, w_eco15607, w_eco15608, w_eco15609, w_eco15610, w_eco15611, w_eco15612, w_eco15613, w_eco15614, w_eco15615, w_eco15616, w_eco15617, w_eco15618, w_eco15619, w_eco15620, w_eco15621, w_eco15622, w_eco15623, w_eco15624, w_eco15625, w_eco15626, w_eco15627, w_eco15628, w_eco15629, w_eco15630, w_eco15631, w_eco15632, w_eco15633, w_eco15634, w_eco15635, w_eco15636, w_eco15637, w_eco15638, w_eco15639, w_eco15640, w_eco15641, w_eco15642, w_eco15643, w_eco15644, w_eco15645, w_eco15646, w_eco15647, w_eco15648, w_eco15649, w_eco15650, w_eco15651, w_eco15652, w_eco15653, w_eco15654, w_eco15655, w_eco15656, w_eco15657, w_eco15658, w_eco15659, w_eco15660, w_eco15661, w_eco15662, w_eco15663, w_eco15664, w_eco15665, w_eco15666, w_eco15667, w_eco15668, w_eco15669, w_eco15670, w_eco15671, w_eco15672, w_eco15673, w_eco15674, w_eco15675, w_eco15676, w_eco15677, w_eco15678, w_eco15679, w_eco15680, w_eco15681, w_eco15682, w_eco15683, w_eco15684, w_eco15685, w_eco15686, w_eco15687, w_eco15688, w_eco15689, w_eco15690, w_eco15691, w_eco15692, w_eco15693, w_eco15694, w_eco15695, w_eco15696, w_eco15697, w_eco15698, w_eco15699, w_eco15700, w_eco15701, w_eco15702, w_eco15703, w_eco15704, w_eco15705, w_eco15706, w_eco15707, w_eco15708, w_eco15709, w_eco15710, w_eco15711, w_eco15712, w_eco15713, w_eco15714, w_eco15715, w_eco15716, w_eco15717, w_eco15718, w_eco15719, w_eco15720, w_eco15721, w_eco15722, w_eco15723, w_eco15724, w_eco15725, w_eco15726, w_eco15727, w_eco15728, w_eco15729, w_eco15730, w_eco15731, w_eco15732, w_eco15733, w_eco15734, w_eco15735, w_eco15736, w_eco15737, w_eco15738, w_eco15739, w_eco15740, w_eco15741, w_eco15742, w_eco15743, w_eco15744, w_eco15745, w_eco15746, w_eco15747, w_eco15748, w_eco15749, w_eco15750, w_eco15751, w_eco15752, w_eco15753, w_eco15754, w_eco15755, w_eco15756, w_eco15757, w_eco15758, w_eco15759, w_eco15760, w_eco15761, w_eco15762, w_eco15763, w_eco15764, w_eco15765, w_eco15766, w_eco15767, w_eco15768, w_eco15769, w_eco15770, w_eco15771, w_eco15772, w_eco15773, w_eco15774, w_eco15775, w_eco15776, w_eco15777, w_eco15778, w_eco15779, w_eco15780, w_eco15781, w_eco15782, w_eco15783, w_eco15784, w_eco15785, w_eco15786, w_eco15787, w_eco15788, w_eco15789, w_eco15790, w_eco15791, w_eco15792, w_eco15793, w_eco15794, w_eco15795, w_eco15796, w_eco15797, w_eco15798, w_eco15799, w_eco15800, w_eco15801, w_eco15802, w_eco15803, w_eco15804, w_eco15805, w_eco15806, w_eco15807, w_eco15808, w_eco15809, w_eco15810, w_eco15811, w_eco15812, w_eco15813, w_eco15814, w_eco15815, w_eco15816, w_eco15817, w_eco15818, w_eco15819, w_eco15820, w_eco15821, w_eco15822, w_eco15823, w_eco15824, w_eco15825, w_eco15826, w_eco15827, w_eco15828, w_eco15829, w_eco15830, w_eco15831, w_eco15832, w_eco15833, w_eco15834, w_eco15835, w_eco15836, w_eco15837, w_eco15838, w_eco15839, w_eco15840, w_eco15841, w_eco15842, w_eco15843, w_eco15844, w_eco15845, w_eco15846, w_eco15847, w_eco15848, w_eco15849, w_eco15850, w_eco15851, w_eco15852, w_eco15853, w_eco15854, w_eco15855, w_eco15856, w_eco15857, w_eco15858, w_eco15859, w_eco15860, w_eco15861, w_eco15862, w_eco15863, w_eco15864, w_eco15865, w_eco15866, w_eco15867, w_eco15868, w_eco15869, w_eco15870, w_eco15871, w_eco15872, w_eco15873, w_eco15874, w_eco15875, w_eco15876, w_eco15877, w_eco15878, w_eco15879, w_eco15880, w_eco15881, w_eco15882, w_eco15883, w_eco15884, w_eco15885, w_eco15886, w_eco15887, w_eco15888, w_eco15889, w_eco15890, w_eco15891, w_eco15892, w_eco15893, w_eco15894, w_eco15895, w_eco15896, w_eco15897, w_eco15898, w_eco15899, w_eco15900, w_eco15901, w_eco15902, w_eco15903, w_eco15904, w_eco15905, w_eco15906, w_eco15907, w_eco15908, w_eco15909, w_eco15910, w_eco15911, w_eco15912, w_eco15913, w_eco15914, w_eco15915, w_eco15916, w_eco15917, w_eco15918, w_eco15919, w_eco15920, w_eco15921, w_eco15922, w_eco15923, w_eco15924, w_eco15925, w_eco15926, w_eco15927, w_eco15928, w_eco15929, w_eco15930, w_eco15931, w_eco15932, w_eco15933, w_eco15934, w_eco15935, w_eco15936, w_eco15937, w_eco15938, w_eco15939, w_eco15940, w_eco15941, w_eco15942, w_eco15943, w_eco15944, w_eco15945, w_eco15946, w_eco15947, w_eco15948, w_eco15949, w_eco15950, w_eco15951, w_eco15952, w_eco15953, w_eco15954, w_eco15955, w_eco15956, w_eco15957, w_eco15958, w_eco15959, w_eco15960, w_eco15961, w_eco15962, w_eco15963, w_eco15964, w_eco15965, w_eco15966, w_eco15967, w_eco15968, w_eco15969, w_eco15970, w_eco15971, w_eco15972, w_eco15973, w_eco15974, w_eco15975, w_eco15976, w_eco15977, w_eco15978, w_eco15979, w_eco15980, w_eco15981, w_eco15982, w_eco15983, w_eco15984, w_eco15985, w_eco15986, w_eco15987, w_eco15988, w_eco15989, w_eco15990, w_eco15991, w_eco15992, w_eco15993, w_eco15994, w_eco15995, w_eco15996, w_eco15997, w_eco15998, w_eco15999, w_eco16000, w_eco16001, w_eco16002, w_eco16003, w_eco16004, w_eco16005, w_eco16006, w_eco16007, w_eco16008, w_eco16009, w_eco16010, w_eco16011, w_eco16012, w_eco16013, w_eco16014, w_eco16015, w_eco16016, w_eco16017, w_eco16018, w_eco16019, w_eco16020, w_eco16021, w_eco16022, w_eco16023, w_eco16024, w_eco16025, w_eco16026, w_eco16027, w_eco16028, w_eco16029, w_eco16030, w_eco16031, w_eco16032, w_eco16033, w_eco16034, w_eco16035, w_eco16036, w_eco16037, w_eco16038, w_eco16039, w_eco16040, w_eco16041, w_eco16042, w_eco16043, w_eco16044, w_eco16045, w_eco16046, w_eco16047, w_eco16048, w_eco16049, w_eco16050, w_eco16051, w_eco16052, w_eco16053, w_eco16054, w_eco16055, w_eco16056, w_eco16057, w_eco16058, w_eco16059, w_eco16060, w_eco16061, w_eco16062, w_eco16063, w_eco16064, w_eco16065, w_eco16066, w_eco16067, w_eco16068, w_eco16069, w_eco16070, w_eco16071, w_eco16072, w_eco16073, w_eco16074, w_eco16075, w_eco16076, w_eco16077, w_eco16078, w_eco16079, w_eco16080, w_eco16081, w_eco16082, w_eco16083, w_eco16084, w_eco16085, w_eco16086, w_eco16087, w_eco16088, w_eco16089, w_eco16090, w_eco16091, w_eco16092, w_eco16093, w_eco16094, w_eco16095, w_eco16096, w_eco16097, w_eco16098, w_eco16099, w_eco16100, w_eco16101, w_eco16102, w_eco16103, w_eco16104, w_eco16105, w_eco16106, w_eco16107, w_eco16108, w_eco16109, w_eco16110, w_eco16111, w_eco16112, w_eco16113, w_eco16114, w_eco16115, w_eco16116, w_eco16117, w_eco16118, w_eco16119, w_eco16120, w_eco16121, w_eco16122, w_eco16123, w_eco16124, w_eco16125, w_eco16126, w_eco16127, w_eco16128, w_eco16129, w_eco16130, w_eco16131, w_eco16132, w_eco16133, w_eco16134, w_eco16135, w_eco16136, w_eco16137, w_eco16138, w_eco16139, w_eco16140, w_eco16141, w_eco16142, w_eco16143, w_eco16144, w_eco16145, w_eco16146, w_eco16147, w_eco16148, w_eco16149, w_eco16150, w_eco16151, w_eco16152, w_eco16153, w_eco16154, w_eco16155, w_eco16156, w_eco16157, w_eco16158, w_eco16159, w_eco16160, w_eco16161, w_eco16162, w_eco16163, w_eco16164, w_eco16165, w_eco16166, w_eco16167, w_eco16168, w_eco16169, w_eco16170, w_eco16171, w_eco16172, w_eco16173, w_eco16174, w_eco16175, w_eco16176, w_eco16177, w_eco16178, w_eco16179, w_eco16180, w_eco16181, w_eco16182, w_eco16183, w_eco16184, w_eco16185, w_eco16186, w_eco16187, w_eco16188, w_eco16189, w_eco16190, w_eco16191, w_eco16192, w_eco16193, w_eco16194, w_eco16195, w_eco16196, w_eco16197, w_eco16198, w_eco16199, w_eco16200, w_eco16201, w_eco16202, w_eco16203, w_eco16204, w_eco16205, w_eco16206, w_eco16207, w_eco16208, w_eco16209, w_eco16210, w_eco16211, w_eco16212, w_eco16213, w_eco16214, w_eco16215, w_eco16216, w_eco16217, w_eco16218, w_eco16219, w_eco16220, w_eco16221, w_eco16222, w_eco16223, w_eco16224, w_eco16225, w_eco16226, w_eco16227, w_eco16228, w_eco16229, w_eco16230, w_eco16231, w_eco16232, w_eco16233, w_eco16234, w_eco16235, w_eco16236, w_eco16237, w_eco16238, w_eco16239, w_eco16240, w_eco16241, w_eco16242, w_eco16243, w_eco16244, w_eco16245, w_eco16246, w_eco16247, w_eco16248, w_eco16249, w_eco16250, w_eco16251, w_eco16252, w_eco16253, w_eco16254, w_eco16255, w_eco16256, w_eco16257, w_eco16258, w_eco16259, w_eco16260, w_eco16261, w_eco16262, w_eco16263, w_eco16264, w_eco16265, w_eco16266, w_eco16267, w_eco16268, w_eco16269, w_eco16270, w_eco16271, w_eco16272, w_eco16273, w_eco16274, w_eco16275, w_eco16276, w_eco16277, w_eco16278, w_eco16279, w_eco16280, w_eco16281, w_eco16282, w_eco16283, w_eco16284, w_eco16285, w_eco16286, w_eco16287, w_eco16288, w_eco16289, w_eco16290, w_eco16291, w_eco16292, w_eco16293, w_eco16294, w_eco16295, w_eco16296, w_eco16297, w_eco16298, w_eco16299, w_eco16300, w_eco16301, w_eco16302, w_eco16303, w_eco16304, w_eco16305, w_eco16306, w_eco16307, w_eco16308, w_eco16309, w_eco16310, w_eco16311, w_eco16312, w_eco16313, w_eco16314, w_eco16315, w_eco16316, w_eco16317, w_eco16318, w_eco16319, w_eco16320, w_eco16321, w_eco16322, w_eco16323, w_eco16324, w_eco16325, w_eco16326, w_eco16327, w_eco16328, w_eco16329, w_eco16330, w_eco16331, w_eco16332, w_eco16333, w_eco16334, w_eco16335, w_eco16336, w_eco16337, w_eco16338, w_eco16339, w_eco16340, w_eco16341, w_eco16342, w_eco16343, w_eco16344, w_eco16345, w_eco16346, w_eco16347, w_eco16348, w_eco16349, w_eco16350, w_eco16351, w_eco16352, w_eco16353, w_eco16354, w_eco16355, w_eco16356, w_eco16357, w_eco16358, w_eco16359, w_eco16360, w_eco16361, w_eco16362, w_eco16363, w_eco16364, w_eco16365, w_eco16366, w_eco16367, w_eco16368, w_eco16369, w_eco16370, w_eco16371, w_eco16372, w_eco16373, w_eco16374, w_eco16375, w_eco16376, w_eco16377, w_eco16378, w_eco16379, w_eco16380, w_eco16381, w_eco16382, w_eco16383, w_eco16384, w_eco16385, w_eco16386, w_eco16387, w_eco16388, w_eco16389, w_eco16390, w_eco16391, w_eco16392, w_eco16393, w_eco16394, w_eco16395, w_eco16396, w_eco16397, w_eco16398, w_eco16399, w_eco16400, w_eco16401, w_eco16402, w_eco16403, w_eco16404, w_eco16405, w_eco16406, w_eco16407, w_eco16408, w_eco16409, w_eco16410, w_eco16411, w_eco16412, w_eco16413, w_eco16414, w_eco16415, w_eco16416, w_eco16417, w_eco16418, w_eco16419, w_eco16420, w_eco16421, w_eco16422, w_eco16423, w_eco16424, w_eco16425, w_eco16426, w_eco16427, w_eco16428, w_eco16429, w_eco16430, w_eco16431, w_eco16432, w_eco16433, w_eco16434, w_eco16435, w_eco16436, w_eco16437, w_eco16438, w_eco16439, w_eco16440, w_eco16441, w_eco16442, w_eco16443, w_eco16444, w_eco16445, w_eco16446, w_eco16447, w_eco16448, w_eco16449, w_eco16450, w_eco16451, w_eco16452, w_eco16453, w_eco16454, w_eco16455, w_eco16456, w_eco16457, w_eco16458, w_eco16459, w_eco16460, w_eco16461, w_eco16462, w_eco16463, w_eco16464, w_eco16465, w_eco16466, w_eco16467, w_eco16468, w_eco16469, w_eco16470, w_eco16471, w_eco16472, w_eco16473, w_eco16474, w_eco16475, w_eco16476, w_eco16477, w_eco16478, w_eco16479, w_eco16480, w_eco16481, w_eco16482, w_eco16483, w_eco16484, w_eco16485, w_eco16486, w_eco16487, w_eco16488, w_eco16489, w_eco16490, w_eco16491, w_eco16492, w_eco16493, w_eco16494, w_eco16495, w_eco16496, w_eco16497, w_eco16498, w_eco16499, w_eco16500, w_eco16501, w_eco16502, w_eco16503, w_eco16504, w_eco16505, w_eco16506, w_eco16507, w_eco16508, w_eco16509, w_eco16510, w_eco16511, w_eco16512, w_eco16513, w_eco16514, w_eco16515, w_eco16516, w_eco16517, w_eco16518, w_eco16519, w_eco16520, w_eco16521, w_eco16522, w_eco16523, w_eco16524, w_eco16525, w_eco16526, w_eco16527, w_eco16528, w_eco16529, w_eco16530, w_eco16531, w_eco16532, w_eco16533, w_eco16534, w_eco16535, w_eco16536, w_eco16537, w_eco16538, w_eco16539, w_eco16540, w_eco16541, w_eco16542, w_eco16543, w_eco16544, w_eco16545, w_eco16546, w_eco16547, w_eco16548, w_eco16549, w_eco16550, w_eco16551, w_eco16552, w_eco16553, w_eco16554, w_eco16555, w_eco16556, w_eco16557, w_eco16558, w_eco16559, w_eco16560, w_eco16561, w_eco16562, w_eco16563, w_eco16564, w_eco16565, w_eco16566, w_eco16567, w_eco16568, w_eco16569, w_eco16570, w_eco16571, w_eco16572, w_eco16573, w_eco16574, w_eco16575, w_eco16576, w_eco16577, w_eco16578, w_eco16579, w_eco16580, w_eco16581, w_eco16582, w_eco16583, w_eco16584, w_eco16585, w_eco16586, w_eco16587, w_eco16588, w_eco16589, w_eco16590, w_eco16591, w_eco16592, w_eco16593, w_eco16594, w_eco16595, w_eco16596, w_eco16597, w_eco16598, w_eco16599, w_eco16600, w_eco16601, w_eco16602, w_eco16603, w_eco16604, w_eco16605, w_eco16606, w_eco16607, w_eco16608, w_eco16609, w_eco16610, w_eco16611, w_eco16612, w_eco16613, w_eco16614, w_eco16615, w_eco16616, w_eco16617, w_eco16618, w_eco16619, w_eco16620, w_eco16621, w_eco16622, w_eco16623, w_eco16624, w_eco16625, w_eco16626, w_eco16627, w_eco16628, w_eco16629, w_eco16630, w_eco16631, w_eco16632, w_eco16633, w_eco16634, w_eco16635, w_eco16636, w_eco16637, w_eco16638, w_eco16639, w_eco16640, w_eco16641, w_eco16642, w_eco16643, w_eco16644, w_eco16645, w_eco16646, w_eco16647, w_eco16648, w_eco16649, w_eco16650, w_eco16651, w_eco16652, w_eco16653, w_eco16654, w_eco16655, w_eco16656, w_eco16657, w_eco16658, w_eco16659, w_eco16660, w_eco16661, w_eco16662, w_eco16663, w_eco16664, w_eco16665, w_eco16666, w_eco16667, w_eco16668, w_eco16669, w_eco16670, w_eco16671, w_eco16672, w_eco16673, w_eco16674, w_eco16675, w_eco16676, w_eco16677, w_eco16678, w_eco16679, w_eco16680, w_eco16681, w_eco16682, w_eco16683, w_eco16684, w_eco16685, w_eco16686, w_eco16687, w_eco16688, w_eco16689, w_eco16690, w_eco16691, w_eco16692, w_eco16693, w_eco16694, w_eco16695, w_eco16696, w_eco16697, w_eco16698, w_eco16699, w_eco16700, w_eco16701, w_eco16702, w_eco16703, w_eco16704, w_eco16705, w_eco16706, w_eco16707, w_eco16708, w_eco16709, w_eco16710, w_eco16711, w_eco16712, w_eco16713, w_eco16714, w_eco16715, w_eco16716, w_eco16717, w_eco16718, w_eco16719, w_eco16720, w_eco16721, w_eco16722, w_eco16723, w_eco16724, w_eco16725, w_eco16726, w_eco16727, w_eco16728, w_eco16729, w_eco16730, w_eco16731, w_eco16732, w_eco16733, w_eco16734, w_eco16735, w_eco16736, w_eco16737, w_eco16738, w_eco16739, w_eco16740, w_eco16741, w_eco16742, w_eco16743, w_eco16744, w_eco16745, w_eco16746, w_eco16747, w_eco16748, w_eco16749, w_eco16750, w_eco16751, w_eco16752, w_eco16753, w_eco16754, w_eco16755, w_eco16756, w_eco16757, w_eco16758, w_eco16759, w_eco16760, w_eco16761, w_eco16762, w_eco16763, w_eco16764, w_eco16765, w_eco16766, w_eco16767, w_eco16768, w_eco16769, w_eco16770, w_eco16771, w_eco16772, w_eco16773, w_eco16774, w_eco16775, w_eco16776, w_eco16777, w_eco16778, w_eco16779, w_eco16780, w_eco16781, w_eco16782, w_eco16783, w_eco16784, w_eco16785, w_eco16786, w_eco16787, w_eco16788, w_eco16789, w_eco16790, w_eco16791, w_eco16792, w_eco16793, w_eco16794, w_eco16795, w_eco16796, w_eco16797, w_eco16798, w_eco16799, w_eco16800, w_eco16801, w_eco16802, w_eco16803, w_eco16804, w_eco16805, w_eco16806, w_eco16807, w_eco16808, w_eco16809, w_eco16810, w_eco16811, w_eco16812, w_eco16813, w_eco16814, w_eco16815, w_eco16816, w_eco16817, w_eco16818, w_eco16819, w_eco16820, w_eco16821, w_eco16822, w_eco16823, w_eco16824, w_eco16825, w_eco16826, w_eco16827, w_eco16828, w_eco16829, w_eco16830, w_eco16831, w_eco16832, w_eco16833, w_eco16834, w_eco16835, w_eco16836, w_eco16837, w_eco16838, w_eco16839, w_eco16840, w_eco16841, w_eco16842, w_eco16843, w_eco16844, w_eco16845, w_eco16846, w_eco16847, w_eco16848, w_eco16849, w_eco16850, w_eco16851, w_eco16852, w_eco16853, w_eco16854, w_eco16855, w_eco16856, w_eco16857, w_eco16858, w_eco16859, w_eco16860, w_eco16861, w_eco16862, w_eco16863, w_eco16864, w_eco16865, w_eco16866, w_eco16867, w_eco16868, w_eco16869, w_eco16870, w_eco16871, w_eco16872, w_eco16873, w_eco16874, w_eco16875, w_eco16876, w_eco16877, w_eco16878, w_eco16879, w_eco16880, w_eco16881, w_eco16882, w_eco16883, w_eco16884, w_eco16885, w_eco16886, w_eco16887, w_eco16888, w_eco16889, w_eco16890, w_eco16891, w_eco16892, w_eco16893, w_eco16894, w_eco16895, w_eco16896, w_eco16897, w_eco16898, w_eco16899, w_eco16900, w_eco16901, w_eco16902, w_eco16903, w_eco16904, w_eco16905, w_eco16906, w_eco16907, w_eco16908, w_eco16909, w_eco16910, w_eco16911, w_eco16912, w_eco16913, w_eco16914, w_eco16915, w_eco16916, w_eco16917, w_eco16918, w_eco16919, w_eco16920, w_eco16921, w_eco16922, w_eco16923, w_eco16924, w_eco16925, w_eco16926, w_eco16927, w_eco16928, w_eco16929, w_eco16930, w_eco16931, w_eco16932, w_eco16933, w_eco16934, w_eco16935, w_eco16936, w_eco16937, w_eco16938, w_eco16939, w_eco16940, w_eco16941, w_eco16942, w_eco16943, w_eco16944, w_eco16945, w_eco16946, w_eco16947, w_eco16948, w_eco16949, w_eco16950, w_eco16951, w_eco16952, w_eco16953, w_eco16954, w_eco16955, w_eco16956, w_eco16957, w_eco16958, w_eco16959, w_eco16960, w_eco16961, w_eco16962, w_eco16963, w_eco16964, w_eco16965, w_eco16966, w_eco16967, w_eco16968, w_eco16969, w_eco16970, w_eco16971, w_eco16972, w_eco16973, w_eco16974, w_eco16975, w_eco16976, w_eco16977, w_eco16978, w_eco16979, w_eco16980, w_eco16981, w_eco16982, w_eco16983, w_eco16984, w_eco16985, w_eco16986, w_eco16987, w_eco16988, w_eco16989, w_eco16990, w_eco16991, w_eco16992, w_eco16993, w_eco16994, w_eco16995, w_eco16996, w_eco16997, w_eco16998, w_eco16999, w_eco17000, w_eco17001, w_eco17002, w_eco17003, w_eco17004, w_eco17005, w_eco17006, w_eco17007, w_eco17008, w_eco17009, w_eco17010, w_eco17011, w_eco17012, w_eco17013, w_eco17014, w_eco17015, w_eco17016, w_eco17017, w_eco17018, w_eco17019, w_eco17020, w_eco17021, w_eco17022, w_eco17023, w_eco17024, w_eco17025, w_eco17026, w_eco17027, w_eco17028, w_eco17029, w_eco17030, w_eco17031, w_eco17032, w_eco17033, w_eco17034, w_eco17035, w_eco17036, w_eco17037, w_eco17038, w_eco17039, w_eco17040, w_eco17041, w_eco17042, w_eco17043, w_eco17044, w_eco17045, w_eco17046, w_eco17047, w_eco17048, w_eco17049, w_eco17050, w_eco17051, w_eco17052, w_eco17053, w_eco17054, w_eco17055, w_eco17056, w_eco17057, w_eco17058, w_eco17059, w_eco17060, w_eco17061, w_eco17062, w_eco17063, w_eco17064, w_eco17065, w_eco17066, w_eco17067, w_eco17068, w_eco17069, w_eco17070, w_eco17071, w_eco17072, w_eco17073, w_eco17074, w_eco17075, w_eco17076, w_eco17077, w_eco17078, w_eco17079, w_eco17080, w_eco17081, w_eco17082, w_eco17083, w_eco17084, w_eco17085, w_eco17086, w_eco17087, w_eco17088, w_eco17089, w_eco17090, w_eco17091, w_eco17092, w_eco17093, w_eco17094, w_eco17095, w_eco17096, w_eco17097, w_eco17098, w_eco17099, w_eco17100, w_eco17101, w_eco17102, w_eco17103, w_eco17104, w_eco17105, w_eco17106, w_eco17107, w_eco17108, w_eco17109, w_eco17110, w_eco17111, w_eco17112, w_eco17113, w_eco17114, w_eco17115, w_eco17116, w_eco17117, w_eco17118, w_eco17119, w_eco17120, w_eco17121, w_eco17122, w_eco17123, w_eco17124, w_eco17125, w_eco17126, w_eco17127, w_eco17128, w_eco17129, w_eco17130, w_eco17131, w_eco17132, w_eco17133, w_eco17134, w_eco17135, w_eco17136, w_eco17137, w_eco17138, w_eco17139, w_eco17140, w_eco17141, w_eco17142, w_eco17143, w_eco17144, w_eco17145, w_eco17146, w_eco17147, w_eco17148, w_eco17149, w_eco17150, w_eco17151, w_eco17152, w_eco17153, w_eco17154, w_eco17155, w_eco17156, w_eco17157, w_eco17158, w_eco17159, w_eco17160, w_eco17161, w_eco17162, w_eco17163, w_eco17164, w_eco17165, w_eco17166, w_eco17167, w_eco17168, w_eco17169, w_eco17170, w_eco17171, w_eco17172, w_eco17173, w_eco17174, w_eco17175, w_eco17176, w_eco17177, w_eco17178, w_eco17179, w_eco17180, w_eco17181, w_eco17182, w_eco17183, w_eco17184, w_eco17185, w_eco17186, w_eco17187, w_eco17188, w_eco17189, w_eco17190, w_eco17191, w_eco17192, w_eco17193, w_eco17194, w_eco17195, w_eco17196, w_eco17197, w_eco17198, w_eco17199, w_eco17200, w_eco17201, w_eco17202, w_eco17203, w_eco17204, w_eco17205, w_eco17206, w_eco17207, w_eco17208, w_eco17209, w_eco17210, w_eco17211, w_eco17212, w_eco17213, w_eco17214, w_eco17215, w_eco17216, w_eco17217, w_eco17218, w_eco17219, w_eco17220, w_eco17221, w_eco17222, w_eco17223, w_eco17224, w_eco17225, w_eco17226, w_eco17227, w_eco17228, w_eco17229, w_eco17230, w_eco17231, w_eco17232, w_eco17233, w_eco17234, w_eco17235, w_eco17236, w_eco17237, w_eco17238, w_eco17239, w_eco17240, w_eco17241, w_eco17242, w_eco17243, w_eco17244, w_eco17245, w_eco17246, w_eco17247, w_eco17248, w_eco17249, w_eco17250, w_eco17251, w_eco17252, w_eco17253, w_eco17254, w_eco17255, w_eco17256, w_eco17257, w_eco17258, w_eco17259, w_eco17260, w_eco17261, w_eco17262, w_eco17263, w_eco17264, w_eco17265, w_eco17266, w_eco17267, w_eco17268, w_eco17269, w_eco17270, w_eco17271, w_eco17272, w_eco17273, w_eco17274, w_eco17275, w_eco17276, w_eco17277, w_eco17278, w_eco17279, w_eco17280, w_eco17281, w_eco17282, w_eco17283, w_eco17284, w_eco17285, w_eco17286, w_eco17287, w_eco17288, w_eco17289, w_eco17290, w_eco17291, w_eco17292, w_eco17293, w_eco17294, w_eco17295, w_eco17296, w_eco17297, w_eco17298, w_eco17299, w_eco17300, w_eco17301, w_eco17302, w_eco17303, w_eco17304, w_eco17305, w_eco17306, w_eco17307, w_eco17308, w_eco17309, w_eco17310, w_eco17311, w_eco17312, w_eco17313, w_eco17314, w_eco17315, w_eco17316, w_eco17317, w_eco17318, w_eco17319, w_eco17320, w_eco17321, w_eco17322, w_eco17323, w_eco17324, w_eco17325, w_eco17326, w_eco17327, w_eco17328, w_eco17329, w_eco17330, w_eco17331, w_eco17332, w_eco17333, w_eco17334, w_eco17335, w_eco17336, w_eco17337, w_eco17338, w_eco17339, w_eco17340, w_eco17341, w_eco17342, w_eco17343, w_eco17344, w_eco17345, w_eco17346, w_eco17347, w_eco17348, w_eco17349, w_eco17350, w_eco17351, w_eco17352, w_eco17353, w_eco17354, w_eco17355, w_eco17356, w_eco17357, w_eco17358, w_eco17359, w_eco17360, w_eco17361, w_eco17362, w_eco17363, w_eco17364, w_eco17365, w_eco17366, w_eco17367, w_eco17368, w_eco17369, w_eco17370, w_eco17371, w_eco17372, w_eco17373, w_eco17374, w_eco17375, w_eco17376, w_eco17377, w_eco17378, w_eco17379, w_eco17380, w_eco17381, w_eco17382, w_eco17383, w_eco17384, w_eco17385, w_eco17386, w_eco17387, w_eco17388, w_eco17389, w_eco17390, w_eco17391, w_eco17392, w_eco17393, w_eco17394, w_eco17395, w_eco17396, w_eco17397, w_eco17398, w_eco17399, w_eco17400, w_eco17401, w_eco17402, w_eco17403, w_eco17404, w_eco17405, w_eco17406, w_eco17407, w_eco17408, w_eco17409, w_eco17410, w_eco17411, w_eco17412, w_eco17413, w_eco17414, w_eco17415, w_eco17416, w_eco17417, w_eco17418, w_eco17419, w_eco17420, w_eco17421, w_eco17422, w_eco17423, w_eco17424, w_eco17425, w_eco17426, w_eco17427, w_eco17428, w_eco17429, w_eco17430, w_eco17431, w_eco17432, w_eco17433, w_eco17434, w_eco17435, w_eco17436, w_eco17437, w_eco17438, w_eco17439, w_eco17440, w_eco17441, w_eco17442, w_eco17443, w_eco17444, w_eco17445, w_eco17446, w_eco17447, w_eco17448, w_eco17449, w_eco17450, w_eco17451, w_eco17452, w_eco17453, w_eco17454, w_eco17455, w_eco17456, w_eco17457, w_eco17458, w_eco17459, w_eco17460, w_eco17461, w_eco17462, w_eco17463, w_eco17464, w_eco17465, w_eco17466, w_eco17467, w_eco17468, w_eco17469, w_eco17470, w_eco17471, w_eco17472, w_eco17473, w_eco17474, w_eco17475, w_eco17476, w_eco17477, w_eco17478, w_eco17479, w_eco17480, w_eco17481, w_eco17482, w_eco17483, w_eco17484, w_eco17485, w_eco17486, w_eco17487, w_eco17488, w_eco17489, w_eco17490, w_eco17491, w_eco17492, w_eco17493, w_eco17494, w_eco17495, w_eco17496, w_eco17497, w_eco17498, w_eco17499, w_eco17500, w_eco17501, w_eco17502, w_eco17503, w_eco17504, w_eco17505, w_eco17506, w_eco17507, w_eco17508, w_eco17509, w_eco17510, w_eco17511, w_eco17512, w_eco17513, w_eco17514, w_eco17515, w_eco17516, w_eco17517, w_eco17518, w_eco17519, w_eco17520, w_eco17521, w_eco17522, w_eco17523, w_eco17524, w_eco17525, w_eco17526, w_eco17527, w_eco17528, w_eco17529, w_eco17530, w_eco17531, w_eco17532, w_eco17533, w_eco17534, w_eco17535, w_eco17536, w_eco17537, w_eco17538, w_eco17539, w_eco17540, w_eco17541, w_eco17542, w_eco17543, w_eco17544, w_eco17545, w_eco17546, w_eco17547, w_eco17548, w_eco17549, w_eco17550, w_eco17551, w_eco17552, w_eco17553, w_eco17554, w_eco17555, w_eco17556, w_eco17557, w_eco17558, w_eco17559, w_eco17560, w_eco17561, w_eco17562, w_eco17563, w_eco17564, w_eco17565, w_eco17566, w_eco17567, w_eco17568, w_eco17569, w_eco17570, w_eco17571, w_eco17572, w_eco17573, w_eco17574, w_eco17575, w_eco17576, w_eco17577, w_eco17578, w_eco17579, w_eco17580, w_eco17581, w_eco17582, w_eco17583, w_eco17584, w_eco17585, w_eco17586, w_eco17587, w_eco17588, w_eco17589, w_eco17590, w_eco17591, w_eco17592, w_eco17593, w_eco17594, w_eco17595, w_eco17596, w_eco17597, w_eco17598, w_eco17599, w_eco17600, w_eco17601, w_eco17602, w_eco17603, w_eco17604, w_eco17605, w_eco17606, w_eco17607, w_eco17608, w_eco17609, w_eco17610, w_eco17611, w_eco17612, w_eco17613, w_eco17614, w_eco17615, w_eco17616, w_eco17617, w_eco17618, w_eco17619, w_eco17620, w_eco17621, w_eco17622, w_eco17623, w_eco17624, w_eco17625, w_eco17626, w_eco17627, w_eco17628, w_eco17629, w_eco17630, w_eco17631, w_eco17632, w_eco17633, w_eco17634, w_eco17635, w_eco17636, w_eco17637, w_eco17638, w_eco17639, w_eco17640, w_eco17641, w_eco17642, w_eco17643, w_eco17644, w_eco17645, w_eco17646, w_eco17647, w_eco17648, w_eco17649, w_eco17650, w_eco17651, w_eco17652, w_eco17653, w_eco17654, w_eco17655, w_eco17656, w_eco17657, w_eco17658, w_eco17659, w_eco17660, w_eco17661, w_eco17662, w_eco17663, w_eco17664, w_eco17665, w_eco17666, w_eco17667, w_eco17668, w_eco17669, w_eco17670, w_eco17671, w_eco17672, w_eco17673, w_eco17674, w_eco17675, w_eco17676, w_eco17677, w_eco17678, w_eco17679, w_eco17680, w_eco17681, w_eco17682, w_eco17683, w_eco17684, w_eco17685, w_eco17686, w_eco17687, w_eco17688, w_eco17689, w_eco17690, w_eco17691, w_eco17692, w_eco17693, w_eco17694, w_eco17695, w_eco17696, w_eco17697, w_eco17698, w_eco17699, w_eco17700, w_eco17701, w_eco17702, w_eco17703, w_eco17704, w_eco17705, w_eco17706, w_eco17707, w_eco17708, w_eco17709, w_eco17710, w_eco17711, w_eco17712, w_eco17713, w_eco17714, w_eco17715, w_eco17716, w_eco17717, w_eco17718, w_eco17719, w_eco17720, w_eco17721, w_eco17722, w_eco17723, w_eco17724, w_eco17725, w_eco17726, w_eco17727, w_eco17728, w_eco17729, w_eco17730, w_eco17731, w_eco17732, w_eco17733, w_eco17734, w_eco17735, w_eco17736, w_eco17737, w_eco17738, w_eco17739, w_eco17740, w_eco17741, w_eco17742, w_eco17743, w_eco17744, w_eco17745, w_eco17746, w_eco17747, w_eco17748, w_eco17749, w_eco17750, w_eco17751, w_eco17752, w_eco17753, w_eco17754, w_eco17755, w_eco17756, w_eco17757, w_eco17758, w_eco17759, w_eco17760, w_eco17761, w_eco17762, w_eco17763, w_eco17764, w_eco17765, w_eco17766, w_eco17767, w_eco17768, w_eco17769, w_eco17770, w_eco17771, w_eco17772, w_eco17773, w_eco17774, w_eco17775, w_eco17776, w_eco17777, w_eco17778, w_eco17779, w_eco17780, w_eco17781, w_eco17782, w_eco17783, w_eco17784, w_eco17785, w_eco17786, w_eco17787, w_eco17788, w_eco17789, w_eco17790, w_eco17791, w_eco17792, w_eco17793, w_eco17794, w_eco17795, w_eco17796, w_eco17797, w_eco17798, w_eco17799, w_eco17800, w_eco17801, w_eco17802, w_eco17803, w_eco17804, w_eco17805, w_eco17806, w_eco17807, w_eco17808, w_eco17809, w_eco17810, w_eco17811, w_eco17812, w_eco17813, w_eco17814, w_eco17815, w_eco17816, w_eco17817, w_eco17818, w_eco17819, w_eco17820, w_eco17821, w_eco17822, w_eco17823, w_eco17824, w_eco17825, w_eco17826, w_eco17827, w_eco17828, w_eco17829, w_eco17830, w_eco17831, w_eco17832, w_eco17833, w_eco17834, w_eco17835, w_eco17836, w_eco17837, w_eco17838, w_eco17839, w_eco17840, w_eco17841, w_eco17842, w_eco17843, w_eco17844, w_eco17845, w_eco17846, w_eco17847, w_eco17848, w_eco17849, w_eco17850, w_eco17851, w_eco17852, w_eco17853, w_eco17854, w_eco17855, w_eco17856, w_eco17857, w_eco17858, w_eco17859, w_eco17860, w_eco17861, w_eco17862, w_eco17863, w_eco17864, w_eco17865, w_eco17866, w_eco17867, w_eco17868, w_eco17869, w_eco17870, w_eco17871, w_eco17872, w_eco17873, w_eco17874, w_eco17875, w_eco17876, w_eco17877, w_eco17878, w_eco17879, w_eco17880, w_eco17881, w_eco17882, w_eco17883, w_eco17884, w_eco17885, w_eco17886, w_eco17887, w_eco17888, w_eco17889, w_eco17890, w_eco17891, w_eco17892, w_eco17893, w_eco17894, w_eco17895, w_eco17896, w_eco17897, w_eco17898, w_eco17899, w_eco17900, w_eco17901, w_eco17902, w_eco17903, w_eco17904, w_eco17905, w_eco17906, w_eco17907, w_eco17908, w_eco17909, w_eco17910, w_eco17911, w_eco17912, w_eco17913, w_eco17914, w_eco17915, w_eco17916, w_eco17917, w_eco17918, w_eco17919, w_eco17920, w_eco17921, w_eco17922, w_eco17923, w_eco17924, w_eco17925, w_eco17926, w_eco17927, w_eco17928, w_eco17929, w_eco17930, w_eco17931, w_eco17932, w_eco17933, w_eco17934, w_eco17935, w_eco17936, w_eco17937, w_eco17938, w_eco17939, w_eco17940, w_eco17941, w_eco17942, w_eco17943, w_eco17944, w_eco17945, w_eco17946, w_eco17947, w_eco17948, w_eco17949, w_eco17950, w_eco17951, w_eco17952, w_eco17953, w_eco17954, w_eco17955, w_eco17956, w_eco17957, w_eco17958, w_eco17959, w_eco17960, w_eco17961, w_eco17962, w_eco17963, w_eco17964, w_eco17965, w_eco17966, w_eco17967, w_eco17968, w_eco17969, w_eco17970, w_eco17971, w_eco17972, w_eco17973, w_eco17974, w_eco17975, w_eco17976, w_eco17977, w_eco17978, w_eco17979, w_eco17980, w_eco17981, w_eco17982, w_eco17983, w_eco17984, w_eco17985, w_eco17986, w_eco17987, w_eco17988, w_eco17989, w_eco17990, w_eco17991, w_eco17992, w_eco17993, w_eco17994, w_eco17995, w_eco17996, w_eco17997, w_eco17998, w_eco17999, w_eco18000, w_eco18001, w_eco18002, w_eco18003, w_eco18004, w_eco18005, w_eco18006, w_eco18007, w_eco18008, w_eco18009, w_eco18010, w_eco18011, w_eco18012, w_eco18013, w_eco18014, w_eco18015, w_eco18016, w_eco18017, w_eco18018, w_eco18019, w_eco18020, w_eco18021, w_eco18022, w_eco18023, w_eco18024, w_eco18025, w_eco18026, w_eco18027, w_eco18028, w_eco18029, w_eco18030, w_eco18031, w_eco18032, w_eco18033, w_eco18034, w_eco18035, w_eco18036, w_eco18037, w_eco18038, w_eco18039, w_eco18040, w_eco18041, w_eco18042, w_eco18043, w_eco18044, w_eco18045, w_eco18046, w_eco18047, w_eco18048, w_eco18049, w_eco18050, w_eco18051, w_eco18052, w_eco18053, w_eco18054, w_eco18055, w_eco18056, w_eco18057, w_eco18058, w_eco18059, w_eco18060, w_eco18061, w_eco18062, w_eco18063, w_eco18064, w_eco18065, w_eco18066, w_eco18067, w_eco18068, w_eco18069, w_eco18070, w_eco18071, w_eco18072, w_eco18073, w_eco18074, w_eco18075, w_eco18076, w_eco18077, w_eco18078, w_eco18079, w_eco18080, w_eco18081, w_eco18082, w_eco18083, w_eco18084, w_eco18085, w_eco18086, w_eco18087, w_eco18088, w_eco18089, w_eco18090, w_eco18091, w_eco18092, w_eco18093, w_eco18094, w_eco18095, w_eco18096, w_eco18097, w_eco18098, w_eco18099, w_eco18100, w_eco18101, w_eco18102, w_eco18103, w_eco18104, w_eco18105, w_eco18106, w_eco18107, w_eco18108, w_eco18109, w_eco18110, w_eco18111, w_eco18112, w_eco18113, w_eco18114, w_eco18115, w_eco18116, w_eco18117, w_eco18118, w_eco18119, w_eco18120, w_eco18121, w_eco18122, w_eco18123, w_eco18124, w_eco18125, w_eco18126, w_eco18127, w_eco18128, w_eco18129, w_eco18130, w_eco18131, w_eco18132, w_eco18133, w_eco18134, w_eco18135, w_eco18136, w_eco18137, w_eco18138, w_eco18139, w_eco18140, w_eco18141, w_eco18142, w_eco18143, w_eco18144, w_eco18145, w_eco18146, w_eco18147, w_eco18148, w_eco18149, w_eco18150, w_eco18151, w_eco18152, w_eco18153, w_eco18154, w_eco18155, w_eco18156, w_eco18157, w_eco18158, w_eco18159, w_eco18160, w_eco18161, w_eco18162, w_eco18163, w_eco18164, w_eco18165, w_eco18166, w_eco18167, w_eco18168, w_eco18169, w_eco18170, w_eco18171, w_eco18172, w_eco18173, w_eco18174, w_eco18175, w_eco18176, w_eco18177, w_eco18178, w_eco18179, w_eco18180, w_eco18181, w_eco18182, w_eco18183, w_eco18184, w_eco18185, w_eco18186, w_eco18187, w_eco18188, w_eco18189, w_eco18190, w_eco18191, w_eco18192, w_eco18193, w_eco18194, w_eco18195, w_eco18196, w_eco18197, w_eco18198, w_eco18199, w_eco18200, w_eco18201, w_eco18202, w_eco18203, w_eco18204, w_eco18205, w_eco18206, w_eco18207, w_eco18208, w_eco18209, w_eco18210, w_eco18211, w_eco18212, w_eco18213, w_eco18214, w_eco18215, w_eco18216, w_eco18217, w_eco18218, w_eco18219, w_eco18220, w_eco18221, w_eco18222, w_eco18223, w_eco18224, w_eco18225, w_eco18226, w_eco18227, w_eco18228, w_eco18229, w_eco18230, w_eco18231, w_eco18232, w_eco18233, w_eco18234, w_eco18235, w_eco18236, w_eco18237, w_eco18238, w_eco18239, w_eco18240, w_eco18241, w_eco18242, w_eco18243, w_eco18244, w_eco18245, w_eco18246, w_eco18247, w_eco18248, w_eco18249, w_eco18250, w_eco18251, w_eco18252, w_eco18253, w_eco18254, w_eco18255, w_eco18256, w_eco18257, w_eco18258, w_eco18259, w_eco18260, w_eco18261, w_eco18262, w_eco18263, w_eco18264, w_eco18265, w_eco18266, w_eco18267, w_eco18268, w_eco18269, w_eco18270, w_eco18271, w_eco18272, w_eco18273, w_eco18274, w_eco18275, w_eco18276, w_eco18277, w_eco18278, w_eco18279, w_eco18280, w_eco18281, w_eco18282, w_eco18283, w_eco18284, w_eco18285, w_eco18286, w_eco18287, w_eco18288, w_eco18289, w_eco18290, w_eco18291, w_eco18292, w_eco18293, w_eco18294, w_eco18295, w_eco18296, w_eco18297, w_eco18298, w_eco18299, w_eco18300, w_eco18301, w_eco18302, w_eco18303, w_eco18304, w_eco18305, w_eco18306, w_eco18307, w_eco18308, w_eco18309, w_eco18310, w_eco18311, w_eco18312, w_eco18313, w_eco18314, w_eco18315, w_eco18316, w_eco18317, w_eco18318, w_eco18319, w_eco18320, w_eco18321, w_eco18322, w_eco18323, w_eco18324, w_eco18325, w_eco18326, w_eco18327, w_eco18328, w_eco18329, w_eco18330, w_eco18331, w_eco18332, w_eco18333, w_eco18334, w_eco18335, w_eco18336, w_eco18337, w_eco18338, w_eco18339, w_eco18340, w_eco18341, w_eco18342, w_eco18343, w_eco18344, w_eco18345, w_eco18346, w_eco18347, w_eco18348, w_eco18349, w_eco18350, w_eco18351, w_eco18352, w_eco18353, w_eco18354, w_eco18355, w_eco18356, w_eco18357, w_eco18358, w_eco18359, w_eco18360, w_eco18361, w_eco18362, w_eco18363, w_eco18364, w_eco18365, w_eco18366, w_eco18367, w_eco18368, w_eco18369, w_eco18370, w_eco18371, w_eco18372, w_eco18373, w_eco18374, w_eco18375, w_eco18376, w_eco18377, w_eco18378, w_eco18379, w_eco18380, w_eco18381, w_eco18382, w_eco18383, w_eco18384, w_eco18385, w_eco18386, w_eco18387, w_eco18388, w_eco18389, w_eco18390, w_eco18391, w_eco18392, w_eco18393, w_eco18394, w_eco18395, w_eco18396, w_eco18397, w_eco18398, w_eco18399, w_eco18400, w_eco18401, w_eco18402, w_eco18403, w_eco18404, w_eco18405, w_eco18406, w_eco18407, w_eco18408, w_eco18409, w_eco18410, w_eco18411, w_eco18412, w_eco18413, w_eco18414, w_eco18415, w_eco18416, w_eco18417, w_eco18418, w_eco18419, w_eco18420, w_eco18421, w_eco18422, w_eco18423, w_eco18424, w_eco18425, w_eco18426, w_eco18427, w_eco18428, w_eco18429, w_eco18430, w_eco18431, w_eco18432, w_eco18433, w_eco18434, w_eco18435, w_eco18436, w_eco18437, w_eco18438, w_eco18439, w_eco18440, w_eco18441, w_eco18442, w_eco18443, w_eco18444, w_eco18445, w_eco18446, w_eco18447, w_eco18448, w_eco18449, w_eco18450, w_eco18451, w_eco18452, w_eco18453, w_eco18454, w_eco18455, w_eco18456, w_eco18457, w_eco18458, w_eco18459, w_eco18460, w_eco18461, w_eco18462, w_eco18463, w_eco18464, w_eco18465, w_eco18466, w_eco18467, w_eco18468, w_eco18469, w_eco18470, w_eco18471, w_eco18472, w_eco18473, w_eco18474, w_eco18475, w_eco18476, w_eco18477, w_eco18478, w_eco18479, w_eco18480, w_eco18481, w_eco18482, w_eco18483, w_eco18484, w_eco18485, w_eco18486, w_eco18487, w_eco18488, w_eco18489, w_eco18490, w_eco18491, w_eco18492, w_eco18493, w_eco18494, w_eco18495, w_eco18496, w_eco18497, w_eco18498, w_eco18499, w_eco18500, w_eco18501, w_eco18502, w_eco18503, w_eco18504, w_eco18505, w_eco18506, w_eco18507, w_eco18508, w_eco18509, w_eco18510, w_eco18511, w_eco18512, w_eco18513, w_eco18514, w_eco18515, w_eco18516, w_eco18517, w_eco18518, w_eco18519, w_eco18520, w_eco18521, w_eco18522, w_eco18523, w_eco18524, w_eco18525, w_eco18526, w_eco18527, w_eco18528, w_eco18529, w_eco18530, w_eco18531, w_eco18532, w_eco18533, w_eco18534, w_eco18535, w_eco18536, w_eco18537, w_eco18538, w_eco18539, w_eco18540, w_eco18541, w_eco18542, w_eco18543, w_eco18544, w_eco18545, w_eco18546, w_eco18547, w_eco18548, w_eco18549, w_eco18550, w_eco18551, w_eco18552, w_eco18553, w_eco18554, w_eco18555, w_eco18556, w_eco18557, w_eco18558, w_eco18559, w_eco18560, w_eco18561, w_eco18562, w_eco18563, w_eco18564, w_eco18565, w_eco18566, w_eco18567, w_eco18568, w_eco18569, w_eco18570, w_eco18571, w_eco18572, w_eco18573, w_eco18574, w_eco18575, w_eco18576, w_eco18577, w_eco18578, w_eco18579, w_eco18580, w_eco18581, w_eco18582, w_eco18583, w_eco18584, w_eco18585, w_eco18586, w_eco18587, w_eco18588, w_eco18589, w_eco18590, w_eco18591, w_eco18592, w_eco18593, w_eco18594, w_eco18595, w_eco18596, w_eco18597, w_eco18598, w_eco18599, w_eco18600, w_eco18601, w_eco18602, w_eco18603, w_eco18604, w_eco18605, w_eco18606, w_eco18607, w_eco18608, w_eco18609, w_eco18610, w_eco18611, w_eco18612, w_eco18613, w_eco18614, w_eco18615, w_eco18616, w_eco18617, w_eco18618, w_eco18619, w_eco18620, w_eco18621, w_eco18622, w_eco18623, w_eco18624, w_eco18625, w_eco18626, w_eco18627, w_eco18628, w_eco18629, w_eco18630, w_eco18631, w_eco18632, w_eco18633, w_eco18634, w_eco18635, w_eco18636, w_eco18637, w_eco18638, w_eco18639, w_eco18640, w_eco18641, w_eco18642, w_eco18643, w_eco18644, w_eco18645, w_eco18646, w_eco18647, w_eco18648, w_eco18649, w_eco18650, w_eco18651, w_eco18652, w_eco18653, w_eco18654, w_eco18655, w_eco18656, w_eco18657, w_eco18658, w_eco18659, w_eco18660, w_eco18661, w_eco18662, w_eco18663, w_eco18664, w_eco18665, w_eco18666, w_eco18667, w_eco18668, w_eco18669, w_eco18670, w_eco18671, w_eco18672, w_eco18673, w_eco18674, w_eco18675, w_eco18676, w_eco18677, w_eco18678, w_eco18679, w_eco18680, w_eco18681, w_eco18682, w_eco18683, w_eco18684, w_eco18685, w_eco18686, w_eco18687, w_eco18688, w_eco18689, w_eco18690, w_eco18691, w_eco18692, w_eco18693, w_eco18694, w_eco18695, w_eco18696, w_eco18697, w_eco18698, w_eco18699, w_eco18700, w_eco18701, w_eco18702, w_eco18703, w_eco18704, w_eco18705, w_eco18706, w_eco18707, w_eco18708, w_eco18709, w_eco18710, w_eco18711, w_eco18712, w_eco18713, w_eco18714, w_eco18715, w_eco18716, w_eco18717, w_eco18718, w_eco18719, w_eco18720, w_eco18721, w_eco18722, w_eco18723, w_eco18724, w_eco18725, w_eco18726, w_eco18727, w_eco18728, w_eco18729, w_eco18730, w_eco18731, w_eco18732, w_eco18733, w_eco18734, w_eco18735, w_eco18736, w_eco18737, w_eco18738, w_eco18739, w_eco18740, w_eco18741, w_eco18742, w_eco18743, w_eco18744, w_eco18745, w_eco18746, w_eco18747, w_eco18748, w_eco18749, w_eco18750, w_eco18751, w_eco18752, w_eco18753, w_eco18754, w_eco18755, w_eco18756, w_eco18757, w_eco18758, w_eco18759, w_eco18760, w_eco18761, w_eco18762, w_eco18763, w_eco18764, w_eco18765, w_eco18766, w_eco18767, w_eco18768, w_eco18769, w_eco18770, w_eco18771, w_eco18772, w_eco18773, w_eco18774, w_eco18775, w_eco18776, w_eco18777, w_eco18778, w_eco18779, w_eco18780, w_eco18781, w_eco18782, w_eco18783, w_eco18784, w_eco18785, w_eco18786, w_eco18787, w_eco18788, w_eco18789, w_eco18790, w_eco18791, w_eco18792, w_eco18793, w_eco18794, w_eco18795, w_eco18796, w_eco18797, w_eco18798, w_eco18799, w_eco18800, w_eco18801, w_eco18802, w_eco18803, w_eco18804, w_eco18805, w_eco18806, w_eco18807, w_eco18808, w_eco18809, w_eco18810, w_eco18811, w_eco18812, w_eco18813, w_eco18814, w_eco18815, w_eco18816, w_eco18817, w_eco18818, w_eco18819, w_eco18820, w_eco18821, w_eco18822, w_eco18823, w_eco18824, w_eco18825, w_eco18826, w_eco18827, w_eco18828, w_eco18829, w_eco18830, w_eco18831, w_eco18832, w_eco18833, w_eco18834, w_eco18835, w_eco18836, w_eco18837, w_eco18838, w_eco18839, w_eco18840, w_eco18841, w_eco18842, w_eco18843, w_eco18844, w_eco18845, w_eco18846, w_eco18847, w_eco18848, w_eco18849, w_eco18850, w_eco18851, w_eco18852, w_eco18853, w_eco18854, w_eco18855, w_eco18856, w_eco18857, w_eco18858, w_eco18859, w_eco18860, w_eco18861, w_eco18862, w_eco18863, w_eco18864, w_eco18865, w_eco18866, w_eco18867, w_eco18868, w_eco18869, w_eco18870, w_eco18871, w_eco18872, w_eco18873, w_eco18874, w_eco18875, w_eco18876, w_eco18877, w_eco18878, w_eco18879, w_eco18880, w_eco18881, w_eco18882, w_eco18883, w_eco18884, w_eco18885, w_eco18886, w_eco18887, w_eco18888, w_eco18889, w_eco18890, w_eco18891, w_eco18892, w_eco18893, w_eco18894, w_eco18895, w_eco18896, w_eco18897, w_eco18898, w_eco18899, w_eco18900, w_eco18901, w_eco18902, w_eco18903, w_eco18904, w_eco18905, w_eco18906, w_eco18907, w_eco18908, w_eco18909, w_eco18910, w_eco18911, w_eco18912, w_eco18913, w_eco18914, w_eco18915, w_eco18916, w_eco18917, w_eco18918, w_eco18919, w_eco18920, w_eco18921, w_eco18922, w_eco18923, w_eco18924, w_eco18925, w_eco18926, w_eco18927, w_eco18928, w_eco18929, w_eco18930, w_eco18931, w_eco18932, w_eco18933, w_eco18934, w_eco18935, w_eco18936, w_eco18937, w_eco18938, w_eco18939, w_eco18940, w_eco18941, w_eco18942, w_eco18943, w_eco18944, w_eco18945, w_eco18946, w_eco18947, w_eco18948, w_eco18949, w_eco18950, w_eco18951, w_eco18952, w_eco18953, w_eco18954, w_eco18955, w_eco18956, w_eco18957, w_eco18958, w_eco18959, w_eco18960, w_eco18961, w_eco18962, w_eco18963, w_eco18964, w_eco18965, w_eco18966, w_eco18967, w_eco18968, w_eco18969, w_eco18970, w_eco18971, w_eco18972, w_eco18973, w_eco18974, w_eco18975, w_eco18976, w_eco18977, w_eco18978, w_eco18979, w_eco18980, w_eco18981, w_eco18982, w_eco18983, w_eco18984, w_eco18985, w_eco18986, w_eco18987, w_eco18988, w_eco18989, w_eco18990, w_eco18991, w_eco18992, w_eco18993, w_eco18994, w_eco18995, w_eco18996, w_eco18997, w_eco18998, w_eco18999, w_eco19000, w_eco19001, w_eco19002, w_eco19003, w_eco19004, w_eco19005, w_eco19006, w_eco19007, w_eco19008, w_eco19009, w_eco19010, w_eco19011, w_eco19012, w_eco19013, w_eco19014, w_eco19015, w_eco19016, w_eco19017, w_eco19018, w_eco19019, w_eco19020, w_eco19021, w_eco19022, w_eco19023, w_eco19024, w_eco19025, w_eco19026, w_eco19027, w_eco19028, w_eco19029, w_eco19030, w_eco19031, w_eco19032, w_eco19033, w_eco19034, w_eco19035, w_eco19036, w_eco19037, w_eco19038, w_eco19039, w_eco19040, w_eco19041, w_eco19042, w_eco19043, w_eco19044, w_eco19045, w_eco19046, w_eco19047, w_eco19048, w_eco19049, w_eco19050, w_eco19051, w_eco19052, w_eco19053, w_eco19054, w_eco19055, w_eco19056, w_eco19057, w_eco19058, w_eco19059, w_eco19060, w_eco19061, w_eco19062, w_eco19063, w_eco19064, w_eco19065, w_eco19066, w_eco19067, w_eco19068, w_eco19069, w_eco19070, w_eco19071, w_eco19072, w_eco19073, w_eco19074, w_eco19075, w_eco19076, w_eco19077, w_eco19078, w_eco19079, w_eco19080, w_eco19081, w_eco19082, w_eco19083, w_eco19084, w_eco19085, w_eco19086, w_eco19087, w_eco19088, w_eco19089, w_eco19090, w_eco19091, w_eco19092, w_eco19093, w_eco19094, w_eco19095, w_eco19096, w_eco19097, w_eco19098, w_eco19099, w_eco19100, w_eco19101, w_eco19102, w_eco19103, w_eco19104, w_eco19105, w_eco19106, w_eco19107, w_eco19108, w_eco19109, w_eco19110, w_eco19111, w_eco19112, w_eco19113, w_eco19114, w_eco19115, w_eco19116, w_eco19117, w_eco19118, w_eco19119, w_eco19120, w_eco19121, w_eco19122, w_eco19123, w_eco19124, w_eco19125, w_eco19126, w_eco19127, w_eco19128, w_eco19129, w_eco19130, w_eco19131, w_eco19132, w_eco19133, w_eco19134, w_eco19135, w_eco19136, w_eco19137, w_eco19138, w_eco19139, w_eco19140, w_eco19141, w_eco19142, w_eco19143, w_eco19144, w_eco19145, w_eco19146, w_eco19147, w_eco19148, w_eco19149, w_eco19150, w_eco19151, w_eco19152, w_eco19153, w_eco19154, w_eco19155, w_eco19156, w_eco19157, w_eco19158, w_eco19159, w_eco19160, w_eco19161, w_eco19162, w_eco19163, w_eco19164, w_eco19165, w_eco19166, w_eco19167, w_eco19168, w_eco19169, w_eco19170, w_eco19171, w_eco19172, w_eco19173, w_eco19174, w_eco19175, w_eco19176, w_eco19177, w_eco19178, w_eco19179, w_eco19180, w_eco19181, w_eco19182, w_eco19183, w_eco19184, w_eco19185, w_eco19186, w_eco19187, w_eco19188, w_eco19189, w_eco19190, w_eco19191, w_eco19192, w_eco19193, w_eco19194, w_eco19195, w_eco19196, w_eco19197, w_eco19198, w_eco19199, w_eco19200, w_eco19201, w_eco19202, w_eco19203, w_eco19204, w_eco19205, w_eco19206, w_eco19207, w_eco19208, w_eco19209, w_eco19210, w_eco19211, w_eco19212, w_eco19213, w_eco19214, w_eco19215, w_eco19216, w_eco19217, w_eco19218, w_eco19219, w_eco19220, w_eco19221, w_eco19222, w_eco19223, w_eco19224, w_eco19225, w_eco19226, w_eco19227, w_eco19228, w_eco19229, w_eco19230, w_eco19231, w_eco19232, w_eco19233, w_eco19234, w_eco19235, w_eco19236, w_eco19237, w_eco19238, w_eco19239, w_eco19240, w_eco19241, w_eco19242, w_eco19243, w_eco19244, w_eco19245, w_eco19246, w_eco19247, w_eco19248, w_eco19249, w_eco19250, w_eco19251, w_eco19252, w_eco19253, w_eco19254, w_eco19255, w_eco19256, w_eco19257, w_eco19258, w_eco19259, w_eco19260, w_eco19261, w_eco19262, w_eco19263, w_eco19264, w_eco19265, w_eco19266, w_eco19267, w_eco19268, w_eco19269, w_eco19270, w_eco19271, w_eco19272, w_eco19273, w_eco19274, w_eco19275, w_eco19276, w_eco19277, w_eco19278, w_eco19279, w_eco19280, w_eco19281, w_eco19282, w_eco19283, w_eco19284, w_eco19285, w_eco19286, w_eco19287, w_eco19288, w_eco19289, w_eco19290, w_eco19291, w_eco19292, w_eco19293, w_eco19294, w_eco19295, w_eco19296, w_eco19297, w_eco19298, w_eco19299, w_eco19300, w_eco19301, w_eco19302, w_eco19303, w_eco19304, w_eco19305, w_eco19306, w_eco19307, w_eco19308, w_eco19309, w_eco19310, w_eco19311, w_eco19312, w_eco19313, w_eco19314, w_eco19315, w_eco19316, w_eco19317, w_eco19318, w_eco19319, w_eco19320, w_eco19321, w_eco19322, w_eco19323, w_eco19324, w_eco19325, w_eco19326, w_eco19327, w_eco19328, w_eco19329, w_eco19330, w_eco19331, w_eco19332, w_eco19333, w_eco19334, w_eco19335, w_eco19336, w_eco19337, w_eco19338, w_eco19339, w_eco19340, w_eco19341, w_eco19342, w_eco19343, w_eco19344, w_eco19345, w_eco19346, w_eco19347, w_eco19348, w_eco19349, w_eco19350, w_eco19351, w_eco19352, w_eco19353, w_eco19354, w_eco19355, w_eco19356, w_eco19357, w_eco19358, w_eco19359, w_eco19360, w_eco19361, w_eco19362, w_eco19363, w_eco19364, w_eco19365, w_eco19366, w_eco19367, w_eco19368, w_eco19369, w_eco19370, w_eco19371, w_eco19372, w_eco19373, w_eco19374, w_eco19375, w_eco19376, w_eco19377, w_eco19378, w_eco19379, w_eco19380, w_eco19381, w_eco19382, w_eco19383, w_eco19384, w_eco19385, w_eco19386, w_eco19387, w_eco19388, w_eco19389, w_eco19390, w_eco19391, w_eco19392, w_eco19393, w_eco19394, w_eco19395, w_eco19396, w_eco19397, w_eco19398, w_eco19399, w_eco19400, w_eco19401, w_eco19402, w_eco19403, w_eco19404, w_eco19405, w_eco19406, w_eco19407, w_eco19408, w_eco19409, w_eco19410, w_eco19411, w_eco19412, w_eco19413, w_eco19414, w_eco19415, w_eco19416, w_eco19417, w_eco19418, w_eco19419, w_eco19420, w_eco19421, w_eco19422, w_eco19423, w_eco19424, w_eco19425, w_eco19426, w_eco19427, w_eco19428, w_eco19429, w_eco19430, w_eco19431, w_eco19432, w_eco19433, w_eco19434, w_eco19435, w_eco19436, w_eco19437, w_eco19438, w_eco19439, w_eco19440, w_eco19441, w_eco19442, w_eco19443, w_eco19444, w_eco19445, w_eco19446, w_eco19447, w_eco19448, w_eco19449, w_eco19450, w_eco19451, w_eco19452, w_eco19453, w_eco19454, w_eco19455, w_eco19456, w_eco19457, w_eco19458, w_eco19459, w_eco19460, w_eco19461, w_eco19462, w_eco19463, w_eco19464, w_eco19465, w_eco19466, w_eco19467, w_eco19468, w_eco19469, w_eco19470, w_eco19471, w_eco19472, w_eco19473, w_eco19474, w_eco19475, w_eco19476, w_eco19477, w_eco19478, w_eco19479, w_eco19480, w_eco19481, w_eco19482, w_eco19483, w_eco19484, w_eco19485, w_eco19486, w_eco19487, w_eco19488, w_eco19489, w_eco19490, w_eco19491, w_eco19492, w_eco19493, w_eco19494, w_eco19495, w_eco19496, w_eco19497, w_eco19498, w_eco19499, w_eco19500, w_eco19501, w_eco19502, w_eco19503, w_eco19504, w_eco19505, w_eco19506, w_eco19507, w_eco19508, w_eco19509, w_eco19510, w_eco19511, w_eco19512, w_eco19513, w_eco19514, w_eco19515, w_eco19516, w_eco19517, w_eco19518, w_eco19519, w_eco19520, w_eco19521, w_eco19522, w_eco19523, w_eco19524, w_eco19525, w_eco19526, w_eco19527, w_eco19528, w_eco19529, w_eco19530, w_eco19531, w_eco19532, w_eco19533, w_eco19534, w_eco19535, w_eco19536, w_eco19537, w_eco19538, w_eco19539, w_eco19540, w_eco19541, w_eco19542, w_eco19543, w_eco19544, w_eco19545, w_eco19546, w_eco19547, w_eco19548, w_eco19549, w_eco19550, w_eco19551, w_eco19552, w_eco19553, w_eco19554, w_eco19555, w_eco19556, w_eco19557, w_eco19558, w_eco19559, w_eco19560, w_eco19561, w_eco19562, w_eco19563, w_eco19564, w_eco19565, w_eco19566, w_eco19567, w_eco19568, w_eco19569, w_eco19570, w_eco19571, w_eco19572, w_eco19573, w_eco19574, w_eco19575, w_eco19576, w_eco19577, w_eco19578, w_eco19579, w_eco19580, w_eco19581, w_eco19582, w_eco19583, w_eco19584, w_eco19585, w_eco19586, w_eco19587, w_eco19588, w_eco19589, w_eco19590, w_eco19591, w_eco19592, w_eco19593, w_eco19594, w_eco19595, w_eco19596, w_eco19597, w_eco19598, w_eco19599, w_eco19600, w_eco19601, w_eco19602, w_eco19603, w_eco19604, w_eco19605, w_eco19606, w_eco19607, w_eco19608, w_eco19609, w_eco19610, w_eco19611, w_eco19612, w_eco19613, w_eco19614, w_eco19615, w_eco19616, w_eco19617, w_eco19618, w_eco19619, w_eco19620, w_eco19621, w_eco19622, w_eco19623, w_eco19624, w_eco19625, w_eco19626, w_eco19627, w_eco19628, w_eco19629, w_eco19630, w_eco19631, w_eco19632, w_eco19633, w_eco19634, w_eco19635, w_eco19636, w_eco19637, w_eco19638, w_eco19639, w_eco19640, w_eco19641, w_eco19642, w_eco19643, w_eco19644, w_eco19645, w_eco19646, w_eco19647, w_eco19648, w_eco19649, w_eco19650, w_eco19651, w_eco19652, w_eco19653, w_eco19654, w_eco19655, w_eco19656, w_eco19657, w_eco19658, w_eco19659, w_eco19660, w_eco19661, w_eco19662, w_eco19663, w_eco19664, w_eco19665, w_eco19666, w_eco19667, w_eco19668, w_eco19669, w_eco19670, w_eco19671, w_eco19672, w_eco19673, w_eco19674, w_eco19675, w_eco19676, w_eco19677, w_eco19678, w_eco19679, w_eco19680, w_eco19681, w_eco19682, w_eco19683, w_eco19684, w_eco19685, w_eco19686, w_eco19687, w_eco19688, w_eco19689, w_eco19690, w_eco19691, w_eco19692, w_eco19693, w_eco19694, w_eco19695, w_eco19696, w_eco19697, w_eco19698, w_eco19699, w_eco19700, w_eco19701, w_eco19702, w_eco19703, w_eco19704, w_eco19705, w_eco19706, w_eco19707, w_eco19708, w_eco19709, w_eco19710, w_eco19711, w_eco19712, w_eco19713, w_eco19714, w_eco19715, w_eco19716, w_eco19717, w_eco19718, w_eco19719, w_eco19720, w_eco19721, w_eco19722, w_eco19723, w_eco19724, w_eco19725, w_eco19726, w_eco19727, w_eco19728, w_eco19729, w_eco19730, w_eco19731, w_eco19732, w_eco19733, w_eco19734, w_eco19735, w_eco19736, w_eco19737, w_eco19738, w_eco19739, w_eco19740, w_eco19741, w_eco19742, w_eco19743, w_eco19744, w_eco19745, w_eco19746, w_eco19747, w_eco19748, w_eco19749, w_eco19750, w_eco19751, w_eco19752, w_eco19753, w_eco19754, w_eco19755, w_eco19756, w_eco19757, w_eco19758, w_eco19759, w_eco19760, w_eco19761, w_eco19762, w_eco19763, w_eco19764, w_eco19765, w_eco19766, w_eco19767, w_eco19768, w_eco19769, w_eco19770, w_eco19771, w_eco19772, w_eco19773, w_eco19774, w_eco19775, w_eco19776, w_eco19777, w_eco19778, w_eco19779, w_eco19780, w_eco19781, w_eco19782, w_eco19783, w_eco19784, w_eco19785, w_eco19786, w_eco19787, w_eco19788, w_eco19789, w_eco19790, w_eco19791, w_eco19792, w_eco19793, w_eco19794, w_eco19795, w_eco19796, w_eco19797, w_eco19798, w_eco19799, w_eco19800, w_eco19801, w_eco19802, w_eco19803, w_eco19804, w_eco19805, w_eco19806, w_eco19807, w_eco19808, w_eco19809, w_eco19810, w_eco19811, w_eco19812, w_eco19813, w_eco19814, w_eco19815, w_eco19816, w_eco19817, w_eco19818, w_eco19819, w_eco19820, w_eco19821, w_eco19822, w_eco19823, w_eco19824, w_eco19825, w_eco19826, w_eco19827, w_eco19828, w_eco19829, w_eco19830, w_eco19831, w_eco19832, w_eco19833, w_eco19834, w_eco19835, w_eco19836, w_eco19837, w_eco19838, w_eco19839, w_eco19840, w_eco19841, w_eco19842, w_eco19843, w_eco19844, w_eco19845, w_eco19846, w_eco19847, w_eco19848, w_eco19849, w_eco19850, w_eco19851, w_eco19852, w_eco19853, w_eco19854, w_eco19855, w_eco19856, w_eco19857, w_eco19858, w_eco19859, w_eco19860, w_eco19861, w_eco19862, w_eco19863, w_eco19864, w_eco19865, w_eco19866, w_eco19867, w_eco19868, w_eco19869, w_eco19870, w_eco19871, w_eco19872, w_eco19873, w_eco19874, w_eco19875, w_eco19876, w_eco19877, w_eco19878, w_eco19879, w_eco19880, w_eco19881, w_eco19882, w_eco19883, w_eco19884, w_eco19885, w_eco19886, w_eco19887, w_eco19888, w_eco19889, w_eco19890, w_eco19891, w_eco19892, w_eco19893, w_eco19894, w_eco19895, w_eco19896, w_eco19897, w_eco19898, w_eco19899, w_eco19900, w_eco19901, w_eco19902, w_eco19903, w_eco19904, w_eco19905, w_eco19906, w_eco19907, w_eco19908, w_eco19909, w_eco19910, w_eco19911, w_eco19912, w_eco19913, w_eco19914, w_eco19915, w_eco19916, w_eco19917, w_eco19918, w_eco19919, w_eco19920, w_eco19921, w_eco19922, w_eco19923, w_eco19924, w_eco19925, w_eco19926, w_eco19927, w_eco19928, w_eco19929, w_eco19930, w_eco19931, w_eco19932, w_eco19933, w_eco19934, w_eco19935, w_eco19936, w_eco19937, w_eco19938, w_eco19939, w_eco19940, w_eco19941, w_eco19942, w_eco19943, w_eco19944, w_eco19945, w_eco19946, w_eco19947, w_eco19948, w_eco19949, w_eco19950, w_eco19951, w_eco19952, w_eco19953, w_eco19954, w_eco19955, w_eco19956, w_eco19957, w_eco19958, w_eco19959, w_eco19960, w_eco19961, w_eco19962, w_eco19963, w_eco19964, w_eco19965, w_eco19966, w_eco19967, w_eco19968, w_eco19969, w_eco19970, w_eco19971, w_eco19972, w_eco19973, w_eco19974, w_eco19975, w_eco19976, w_eco19977, w_eco19978, w_eco19979, w_eco19980, w_eco19981, w_eco19982, w_eco19983, w_eco19984, w_eco19985, w_eco19986, w_eco19987, w_eco19988, w_eco19989, w_eco19990, w_eco19991, w_eco19992, w_eco19993, w_eco19994, w_eco19995, w_eco19996, w_eco19997, w_eco19998, w_eco19999, w_eco20000, w_eco20001, w_eco20002, w_eco20003, w_eco20004, w_eco20005, w_eco20006, w_eco20007, w_eco20008, w_eco20009, w_eco20010, w_eco20011, w_eco20012, w_eco20013, w_eco20014, w_eco20015, w_eco20016, w_eco20017, w_eco20018, w_eco20019, w_eco20020, w_eco20021, w_eco20022, w_eco20023, w_eco20024, w_eco20025, w_eco20026, w_eco20027, w_eco20028, w_eco20029, w_eco20030, w_eco20031, w_eco20032, w_eco20033, w_eco20034, w_eco20035, w_eco20036, w_eco20037, w_eco20038, w_eco20039, w_eco20040, w_eco20041, w_eco20042, w_eco20043, w_eco20044, w_eco20045, w_eco20046, w_eco20047, w_eco20048, w_eco20049, w_eco20050, w_eco20051, w_eco20052, w_eco20053, w_eco20054, w_eco20055, w_eco20056, w_eco20057, w_eco20058, w_eco20059, w_eco20060, w_eco20061, w_eco20062, w_eco20063, w_eco20064, w_eco20065, w_eco20066, w_eco20067, w_eco20068, w_eco20069, w_eco20070, w_eco20071, w_eco20072, w_eco20073, w_eco20074, w_eco20075, w_eco20076, w_eco20077, w_eco20078, w_eco20079, w_eco20080, w_eco20081, w_eco20082, w_eco20083, w_eco20084, w_eco20085, w_eco20086, w_eco20087, w_eco20088, w_eco20089, w_eco20090, w_eco20091, w_eco20092, w_eco20093, w_eco20094, w_eco20095, w_eco20096, w_eco20097, w_eco20098, w_eco20099, w_eco20100, w_eco20101, w_eco20102, w_eco20103, w_eco20104, w_eco20105, w_eco20106, w_eco20107, w_eco20108, w_eco20109, w_eco20110, w_eco20111, w_eco20112, w_eco20113, w_eco20114, w_eco20115, w_eco20116, w_eco20117, w_eco20118, w_eco20119, w_eco20120, w_eco20121, w_eco20122, w_eco20123, w_eco20124, w_eco20125, w_eco20126, w_eco20127, w_eco20128, w_eco20129, w_eco20130, w_eco20131, w_eco20132, w_eco20133, w_eco20134, w_eco20135, w_eco20136, w_eco20137, w_eco20138, w_eco20139, w_eco20140, w_eco20141, w_eco20142, w_eco20143, w_eco20144, w_eco20145, w_eco20146, w_eco20147, w_eco20148, w_eco20149, w_eco20150, w_eco20151, w_eco20152, w_eco20153, w_eco20154, w_eco20155, w_eco20156, w_eco20157, w_eco20158, w_eco20159, w_eco20160, w_eco20161, w_eco20162, w_eco20163, w_eco20164, w_eco20165, w_eco20166, w_eco20167, w_eco20168, w_eco20169, w_eco20170, w_eco20171, w_eco20172, w_eco20173, w_eco20174, w_eco20175, w_eco20176, w_eco20177, w_eco20178, w_eco20179, w_eco20180, w_eco20181, w_eco20182, w_eco20183, w_eco20184, w_eco20185, w_eco20186, w_eco20187, w_eco20188, w_eco20189, w_eco20190, w_eco20191, w_eco20192, w_eco20193, w_eco20194, w_eco20195, w_eco20196, w_eco20197, w_eco20198, w_eco20199, w_eco20200, w_eco20201, w_eco20202, w_eco20203, w_eco20204, w_eco20205, w_eco20206, w_eco20207, w_eco20208, w_eco20209, w_eco20210, w_eco20211, w_eco20212, w_eco20213, w_eco20214, w_eco20215, w_eco20216, w_eco20217, w_eco20218, w_eco20219, w_eco20220, w_eco20221, w_eco20222, w_eco20223, w_eco20224, w_eco20225, w_eco20226, w_eco20227, w_eco20228, w_eco20229, w_eco20230, w_eco20231, w_eco20232, w_eco20233, w_eco20234, w_eco20235, w_eco20236, w_eco20237, w_eco20238, w_eco20239, w_eco20240, w_eco20241, w_eco20242, w_eco20243, w_eco20244, w_eco20245, w_eco20246, w_eco20247, w_eco20248, w_eco20249, w_eco20250, w_eco20251, w_eco20252, w_eco20253, w_eco20254, w_eco20255, w_eco20256, w_eco20257, w_eco20258, w_eco20259, w_eco20260, w_eco20261, w_eco20262, w_eco20263, w_eco20264, w_eco20265, w_eco20266, w_eco20267, w_eco20268, w_eco20269, w_eco20270, w_eco20271, w_eco20272, w_eco20273, w_eco20274, w_eco20275, w_eco20276, w_eco20277, w_eco20278, w_eco20279, w_eco20280, w_eco20281, w_eco20282, w_eco20283, w_eco20284, w_eco20285, w_eco20286, w_eco20287, w_eco20288, w_eco20289, w_eco20290, w_eco20291, w_eco20292, w_eco20293, w_eco20294, w_eco20295, w_eco20296, w_eco20297, w_eco20298, w_eco20299, w_eco20300, w_eco20301, w_eco20302, w_eco20303, w_eco20304, w_eco20305, w_eco20306, w_eco20307, w_eco20308, w_eco20309, w_eco20310, w_eco20311, w_eco20312, w_eco20313, w_eco20314, w_eco20315, w_eco20316, w_eco20317, w_eco20318, w_eco20319, w_eco20320, w_eco20321, w_eco20322, w_eco20323, w_eco20324, w_eco20325, w_eco20326, w_eco20327, w_eco20328, w_eco20329, w_eco20330, w_eco20331, w_eco20332, w_eco20333, w_eco20334, w_eco20335, w_eco20336, w_eco20337, w_eco20338, w_eco20339, w_eco20340, w_eco20341, w_eco20342, w_eco20343, w_eco20344, w_eco20345, w_eco20346, w_eco20347, w_eco20348, w_eco20349, w_eco20350, w_eco20351, w_eco20352, w_eco20353, w_eco20354, w_eco20355, w_eco20356, w_eco20357, w_eco20358, w_eco20359, w_eco20360, w_eco20361, w_eco20362, w_eco20363, w_eco20364, w_eco20365, w_eco20366, w_eco20367, w_eco20368, w_eco20369, w_eco20370, w_eco20371, w_eco20372, w_eco20373, w_eco20374, w_eco20375, w_eco20376, w_eco20377, w_eco20378, w_eco20379, w_eco20380, w_eco20381, w_eco20382, w_eco20383, w_eco20384, w_eco20385, w_eco20386, w_eco20387, w_eco20388, w_eco20389, w_eco20390, w_eco20391, w_eco20392, w_eco20393, w_eco20394, w_eco20395, w_eco20396, w_eco20397, w_eco20398, w_eco20399, w_eco20400, w_eco20401, w_eco20402, w_eco20403, w_eco20404, w_eco20405, w_eco20406, w_eco20407, w_eco20408, w_eco20409, w_eco20410, w_eco20411, w_eco20412, w_eco20413, w_eco20414, w_eco20415, w_eco20416, w_eco20417, w_eco20418, w_eco20419, w_eco20420, w_eco20421, w_eco20422, w_eco20423, w_eco20424, w_eco20425, w_eco20426, w_eco20427, w_eco20428, w_eco20429, w_eco20430, w_eco20431, w_eco20432, w_eco20433, w_eco20434, w_eco20435, w_eco20436, w_eco20437, w_eco20438, w_eco20439, w_eco20440, w_eco20441, w_eco20442, w_eco20443, w_eco20444, w_eco20445, w_eco20446, w_eco20447, w_eco20448, w_eco20449, w_eco20450, w_eco20451, w_eco20452, w_eco20453, w_eco20454, w_eco20455, w_eco20456, w_eco20457, w_eco20458, w_eco20459, w_eco20460, w_eco20461, w_eco20462, w_eco20463, w_eco20464, w_eco20465, w_eco20466, w_eco20467, w_eco20468, w_eco20469, w_eco20470, w_eco20471, w_eco20472, w_eco20473, w_eco20474, w_eco20475, w_eco20476, w_eco20477, w_eco20478, w_eco20479, w_eco20480, w_eco20481, w_eco20482, w_eco20483, w_eco20484, w_eco20485, w_eco20486, w_eco20487, w_eco20488, w_eco20489, w_eco20490, w_eco20491, w_eco20492, w_eco20493, w_eco20494, w_eco20495, w_eco20496, w_eco20497, w_eco20498, w_eco20499, w_eco20500, w_eco20501, w_eco20502, w_eco20503, w_eco20504, w_eco20505, w_eco20506, w_eco20507, w_eco20508, w_eco20509, w_eco20510, w_eco20511, w_eco20512, w_eco20513, w_eco20514, w_eco20515, w_eco20516, w_eco20517, w_eco20518, w_eco20519, w_eco20520, w_eco20521, w_eco20522, w_eco20523, w_eco20524, w_eco20525, w_eco20526, w_eco20527, w_eco20528, w_eco20529, w_eco20530, w_eco20531, w_eco20532, w_eco20533, w_eco20534, w_eco20535, w_eco20536, w_eco20537, w_eco20538, w_eco20539, w_eco20540, w_eco20541, w_eco20542, w_eco20543, w_eco20544, w_eco20545, w_eco20546, w_eco20547, w_eco20548, w_eco20549, w_eco20550, w_eco20551, w_eco20552, w_eco20553, w_eco20554, w_eco20555, w_eco20556, w_eco20557, w_eco20558, w_eco20559, w_eco20560, w_eco20561, w_eco20562, w_eco20563, w_eco20564, w_eco20565, w_eco20566, w_eco20567, w_eco20568, w_eco20569, w_eco20570, w_eco20571, w_eco20572, w_eco20573, w_eco20574, w_eco20575, w_eco20576, w_eco20577, w_eco20578, w_eco20579, w_eco20580, w_eco20581, w_eco20582, w_eco20583, w_eco20584, w_eco20585, w_eco20586, w_eco20587, w_eco20588, w_eco20589, w_eco20590, w_eco20591, w_eco20592, w_eco20593, w_eco20594, w_eco20595, w_eco20596, w_eco20597, w_eco20598, w_eco20599, w_eco20600, w_eco20601, w_eco20602, w_eco20603, w_eco20604, w_eco20605, w_eco20606, w_eco20607, w_eco20608, w_eco20609, w_eco20610, w_eco20611, w_eco20612, w_eco20613, w_eco20614, w_eco20615, w_eco20616, w_eco20617, w_eco20618, w_eco20619, w_eco20620, w_eco20621, w_eco20622, w_eco20623, w_eco20624, w_eco20625, w_eco20626, w_eco20627, w_eco20628, w_eco20629, w_eco20630, w_eco20631, w_eco20632, w_eco20633, w_eco20634, w_eco20635, w_eco20636, w_eco20637, w_eco20638, w_eco20639, w_eco20640, w_eco20641, w_eco20642, w_eco20643, w_eco20644, w_eco20645, w_eco20646, w_eco20647, w_eco20648, w_eco20649, w_eco20650, w_eco20651, w_eco20652, w_eco20653, w_eco20654, w_eco20655, w_eco20656, w_eco20657, w_eco20658, w_eco20659, w_eco20660, w_eco20661, w_eco20662, w_eco20663, w_eco20664, w_eco20665, w_eco20666, w_eco20667, w_eco20668, w_eco20669, w_eco20670, w_eco20671, w_eco20672, w_eco20673, w_eco20674, w_eco20675, w_eco20676, w_eco20677, w_eco20678, w_eco20679, w_eco20680, w_eco20681, w_eco20682, w_eco20683, w_eco20684, w_eco20685, w_eco20686, w_eco20687, w_eco20688, w_eco20689, w_eco20690, w_eco20691, w_eco20692, w_eco20693, w_eco20694, w_eco20695, w_eco20696, w_eco20697, w_eco20698, w_eco20699, w_eco20700, w_eco20701, w_eco20702, w_eco20703, w_eco20704, w_eco20705, w_eco20706, w_eco20707, w_eco20708, w_eco20709, w_eco20710, w_eco20711, w_eco20712, w_eco20713, w_eco20714, w_eco20715, w_eco20716, w_eco20717, w_eco20718, w_eco20719, w_eco20720, w_eco20721, w_eco20722, w_eco20723, w_eco20724, w_eco20725, w_eco20726, w_eco20727, w_eco20728, w_eco20729, w_eco20730, w_eco20731, w_eco20732, w_eco20733, w_eco20734, w_eco20735, w_eco20736, w_eco20737, w_eco20738, w_eco20739, w_eco20740, w_eco20741, w_eco20742, w_eco20743, w_eco20744, w_eco20745, w_eco20746, w_eco20747, w_eco20748, w_eco20749, w_eco20750, w_eco20751, w_eco20752, w_eco20753, w_eco20754, w_eco20755, w_eco20756, w_eco20757, w_eco20758, w_eco20759, w_eco20760, w_eco20761, w_eco20762, w_eco20763, w_eco20764, w_eco20765, w_eco20766, w_eco20767, w_eco20768, w_eco20769, w_eco20770, w_eco20771, w_eco20772, w_eco20773, w_eco20774, w_eco20775, w_eco20776, w_eco20777, w_eco20778, w_eco20779, w_eco20780, w_eco20781, w_eco20782, w_eco20783, w_eco20784, w_eco20785, w_eco20786, w_eco20787, w_eco20788, w_eco20789, w_eco20790, w_eco20791, w_eco20792, w_eco20793, w_eco20794, w_eco20795, w_eco20796, w_eco20797, w_eco20798, w_eco20799, w_eco20800, w_eco20801, w_eco20802, w_eco20803, w_eco20804, w_eco20805, w_eco20806, w_eco20807, w_eco20808, w_eco20809, w_eco20810, w_eco20811, w_eco20812, w_eco20813, w_eco20814, w_eco20815, w_eco20816, w_eco20817, w_eco20818, w_eco20819, w_eco20820, w_eco20821, w_eco20822, w_eco20823, w_eco20824, w_eco20825, w_eco20826, w_eco20827, w_eco20828, w_eco20829, w_eco20830, w_eco20831, w_eco20832, w_eco20833, w_eco20834, w_eco20835, w_eco20836, w_eco20837, w_eco20838, w_eco20839, w_eco20840, w_eco20841, w_eco20842, w_eco20843, w_eco20844, w_eco20845, w_eco20846, w_eco20847, w_eco20848, w_eco20849, w_eco20850, w_eco20851, w_eco20852, w_eco20853, w_eco20854, w_eco20855, w_eco20856, w_eco20857, w_eco20858, w_eco20859, w_eco20860, w_eco20861, w_eco20862, w_eco20863, w_eco20864, w_eco20865, w_eco20866, w_eco20867, w_eco20868, w_eco20869, w_eco20870, w_eco20871, w_eco20872, w_eco20873, w_eco20874, w_eco20875, w_eco20876, w_eco20877, w_eco20878, w_eco20879, w_eco20880, w_eco20881, w_eco20882, w_eco20883, w_eco20884, w_eco20885, w_eco20886, w_eco20887, w_eco20888, w_eco20889, w_eco20890, w_eco20891, w_eco20892, w_eco20893, w_eco20894, w_eco20895, w_eco20896, w_eco20897, w_eco20898, w_eco20899, w_eco20900, w_eco20901, w_eco20902, w_eco20903, w_eco20904, w_eco20905, w_eco20906, w_eco20907, w_eco20908, w_eco20909, w_eco20910, w_eco20911, w_eco20912, w_eco20913, w_eco20914, w_eco20915, w_eco20916, w_eco20917, w_eco20918, w_eco20919, w_eco20920, w_eco20921, w_eco20922, w_eco20923, w_eco20924, w_eco20925, w_eco20926, w_eco20927, w_eco20928, w_eco20929, w_eco20930, w_eco20931, w_eco20932, w_eco20933, w_eco20934, w_eco20935, w_eco20936, w_eco20937, w_eco20938, w_eco20939, w_eco20940, w_eco20941, w_eco20942, w_eco20943, w_eco20944, w_eco20945, w_eco20946, w_eco20947, w_eco20948, w_eco20949, w_eco20950, w_eco20951, w_eco20952, w_eco20953, w_eco20954, w_eco20955, w_eco20956, w_eco20957, w_eco20958, w_eco20959, w_eco20960, w_eco20961, w_eco20962, w_eco20963, w_eco20964, w_eco20965, w_eco20966, w_eco20967, w_eco20968, w_eco20969, w_eco20970, w_eco20971, w_eco20972, w_eco20973, w_eco20974, w_eco20975, w_eco20976, w_eco20977, w_eco20978, w_eco20979, w_eco20980, w_eco20981, w_eco20982, w_eco20983, w_eco20984, w_eco20985, w_eco20986, w_eco20987, w_eco20988, w_eco20989, w_eco20990, w_eco20991, w_eco20992, w_eco20993, w_eco20994, w_eco20995, w_eco20996, w_eco20997, w_eco20998, w_eco20999, w_eco21000, w_eco21001, w_eco21002, w_eco21003, w_eco21004, w_eco21005, w_eco21006, w_eco21007, w_eco21008, w_eco21009, w_eco21010, w_eco21011, w_eco21012, w_eco21013, w_eco21014, w_eco21015, w_eco21016, w_eco21017, w_eco21018, w_eco21019, w_eco21020, w_eco21021, w_eco21022, w_eco21023, w_eco21024, w_eco21025, w_eco21026, w_eco21027, w_eco21028, w_eco21029, w_eco21030, w_eco21031, w_eco21032, w_eco21033, w_eco21034, w_eco21035, w_eco21036, w_eco21037, w_eco21038, w_eco21039, w_eco21040, w_eco21041, w_eco21042, w_eco21043, w_eco21044, w_eco21045, w_eco21046, w_eco21047, w_eco21048, w_eco21049, w_eco21050, w_eco21051, w_eco21052, w_eco21053, w_eco21054, w_eco21055, w_eco21056, w_eco21057, w_eco21058, w_eco21059, w_eco21060, w_eco21061, w_eco21062, w_eco21063, w_eco21064, w_eco21065, w_eco21066, w_eco21067, w_eco21068, w_eco21069, w_eco21070, w_eco21071, w_eco21072, w_eco21073, w_eco21074, w_eco21075, w_eco21076, w_eco21077, w_eco21078, w_eco21079, w_eco21080, w_eco21081, w_eco21082, w_eco21083, w_eco21084, w_eco21085, w_eco21086, w_eco21087, w_eco21088, w_eco21089, w_eco21090, w_eco21091, w_eco21092, w_eco21093, w_eco21094, w_eco21095, w_eco21096, w_eco21097, w_eco21098, w_eco21099, w_eco21100, w_eco21101, w_eco21102, w_eco21103, w_eco21104, w_eco21105, w_eco21106, w_eco21107, w_eco21108, w_eco21109, w_eco21110, w_eco21111, w_eco21112, w_eco21113, w_eco21114, w_eco21115, w_eco21116, w_eco21117, w_eco21118, w_eco21119, w_eco21120, w_eco21121, w_eco21122, w_eco21123, w_eco21124, w_eco21125, w_eco21126, w_eco21127, w_eco21128, w_eco21129, w_eco21130, w_eco21131, w_eco21132, w_eco21133, w_eco21134, w_eco21135, w_eco21136, w_eco21137, w_eco21138, w_eco21139, w_eco21140, w_eco21141, w_eco21142, w_eco21143, w_eco21144, w_eco21145, w_eco21146, w_eco21147, w_eco21148, w_eco21149, w_eco21150, w_eco21151, w_eco21152, w_eco21153, w_eco21154, w_eco21155, w_eco21156, w_eco21157, w_eco21158, w_eco21159, w_eco21160, w_eco21161, w_eco21162, w_eco21163, w_eco21164, w_eco21165, w_eco21166, w_eco21167, w_eco21168, w_eco21169, w_eco21170, w_eco21171, w_eco21172, w_eco21173, w_eco21174, w_eco21175, w_eco21176, w_eco21177, w_eco21178, w_eco21179, w_eco21180, w_eco21181, w_eco21182, w_eco21183, w_eco21184, w_eco21185, w_eco21186, w_eco21187, w_eco21188, w_eco21189, w_eco21190, w_eco21191, w_eco21192, w_eco21193, w_eco21194, w_eco21195, w_eco21196, w_eco21197, w_eco21198, w_eco21199, w_eco21200, w_eco21201, w_eco21202, w_eco21203, w_eco21204, w_eco21205, w_eco21206, w_eco21207, w_eco21208, w_eco21209, w_eco21210, w_eco21211, w_eco21212, w_eco21213, w_eco21214, w_eco21215, w_eco21216, w_eco21217, w_eco21218, w_eco21219, w_eco21220, w_eco21221, w_eco21222, w_eco21223, w_eco21224, w_eco21225, w_eco21226, w_eco21227, w_eco21228, w_eco21229, w_eco21230, w_eco21231, w_eco21232, w_eco21233, w_eco21234, w_eco21235, w_eco21236, w_eco21237, w_eco21238, w_eco21239, w_eco21240, w_eco21241, w_eco21242, w_eco21243, w_eco21244, w_eco21245, w_eco21246, w_eco21247, w_eco21248, w_eco21249, w_eco21250, w_eco21251, w_eco21252, w_eco21253, w_eco21254, w_eco21255, w_eco21256, w_eco21257, w_eco21258, w_eco21259, w_eco21260, w_eco21261, w_eco21262, w_eco21263, w_eco21264, w_eco21265, w_eco21266, w_eco21267, w_eco21268, w_eco21269, w_eco21270, w_eco21271, w_eco21272, w_eco21273, w_eco21274, w_eco21275, w_eco21276, w_eco21277, w_eco21278, w_eco21279, w_eco21280, w_eco21281, w_eco21282, w_eco21283, w_eco21284, w_eco21285, w_eco21286, w_eco21287, w_eco21288, w_eco21289, w_eco21290, w_eco21291, w_eco21292, w_eco21293, w_eco21294, w_eco21295, w_eco21296, w_eco21297, w_eco21298, w_eco21299, w_eco21300, w_eco21301, w_eco21302, w_eco21303, w_eco21304, w_eco21305, w_eco21306, w_eco21307, w_eco21308, w_eco21309, w_eco21310, w_eco21311, w_eco21312, w_eco21313, w_eco21314, w_eco21315, w_eco21316, w_eco21317, w_eco21318, w_eco21319, w_eco21320, w_eco21321, w_eco21322, w_eco21323, w_eco21324, w_eco21325, w_eco21326, w_eco21327, w_eco21328, w_eco21329, w_eco21330, w_eco21331, w_eco21332, w_eco21333, w_eco21334, w_eco21335, w_eco21336, w_eco21337, w_eco21338, w_eco21339, w_eco21340, w_eco21341, w_eco21342, w_eco21343, w_eco21344, w_eco21345, w_eco21346, w_eco21347, w_eco21348, w_eco21349, w_eco21350, w_eco21351, w_eco21352, w_eco21353, w_eco21354, w_eco21355, w_eco21356, w_eco21357, w_eco21358, w_eco21359, w_eco21360, w_eco21361, w_eco21362, w_eco21363, w_eco21364, w_eco21365, w_eco21366, w_eco21367, w_eco21368, w_eco21369, w_eco21370, w_eco21371, w_eco21372, w_eco21373, w_eco21374, w_eco21375, w_eco21376, w_eco21377, w_eco21378, w_eco21379, w_eco21380, w_eco21381, w_eco21382, w_eco21383, w_eco21384, w_eco21385, w_eco21386, w_eco21387, w_eco21388, w_eco21389, w_eco21390, w_eco21391, w_eco21392, w_eco21393, w_eco21394, w_eco21395, w_eco21396, w_eco21397, w_eco21398, w_eco21399, w_eco21400, w_eco21401, w_eco21402, w_eco21403, w_eco21404, w_eco21405, w_eco21406, w_eco21407, w_eco21408, w_eco21409, w_eco21410, w_eco21411, w_eco21412, w_eco21413, w_eco21414, w_eco21415, w_eco21416, w_eco21417, w_eco21418, w_eco21419, w_eco21420, w_eco21421, w_eco21422, w_eco21423, w_eco21424, w_eco21425, w_eco21426, w_eco21427, w_eco21428, w_eco21429, w_eco21430, w_eco21431, w_eco21432, w_eco21433, w_eco21434, w_eco21435, w_eco21436, w_eco21437, w_eco21438, w_eco21439, w_eco21440, w_eco21441, w_eco21442, w_eco21443, w_eco21444, w_eco21445, w_eco21446, w_eco21447, w_eco21448, w_eco21449, w_eco21450, w_eco21451, w_eco21452, w_eco21453, w_eco21454, w_eco21455, w_eco21456, w_eco21457, w_eco21458, w_eco21459, w_eco21460, w_eco21461, w_eco21462, w_eco21463, w_eco21464, w_eco21465, w_eco21466, w_eco21467, w_eco21468, w_eco21469, w_eco21470, w_eco21471, w_eco21472, w_eco21473, w_eco21474, w_eco21475, w_eco21476, w_eco21477, w_eco21478, w_eco21479, w_eco21480, w_eco21481, w_eco21482, w_eco21483, w_eco21484, w_eco21485, w_eco21486, w_eco21487, w_eco21488, w_eco21489, w_eco21490, w_eco21491, w_eco21492, w_eco21493, w_eco21494, w_eco21495, w_eco21496, w_eco21497, w_eco21498, w_eco21499, w_eco21500, w_eco21501, w_eco21502, w_eco21503, w_eco21504, w_eco21505, w_eco21506, w_eco21507, w_eco21508, w_eco21509, w_eco21510, w_eco21511, w_eco21512, w_eco21513, w_eco21514, w_eco21515, w_eco21516, w_eco21517, w_eco21518, w_eco21519, w_eco21520, w_eco21521, w_eco21522, w_eco21523, w_eco21524, w_eco21525, w_eco21526, w_eco21527, w_eco21528, w_eco21529, w_eco21530, w_eco21531, w_eco21532, w_eco21533, w_eco21534, w_eco21535, w_eco21536, w_eco21537, w_eco21538, w_eco21539, w_eco21540, w_eco21541, w_eco21542, w_eco21543, w_eco21544, w_eco21545, w_eco21546, w_eco21547, w_eco21548, w_eco21549, w_eco21550, w_eco21551, w_eco21552, w_eco21553, w_eco21554, w_eco21555, w_eco21556, w_eco21557, w_eco21558, w_eco21559, w_eco21560, w_eco21561, w_eco21562, w_eco21563, w_eco21564, w_eco21565, w_eco21566, w_eco21567, w_eco21568, w_eco21569, w_eco21570, w_eco21571, w_eco21572, w_eco21573, w_eco21574, w_eco21575, w_eco21576, w_eco21577, w_eco21578, w_eco21579, w_eco21580, w_eco21581, w_eco21582, w_eco21583, w_eco21584, w_eco21585, w_eco21586, w_eco21587, w_eco21588, w_eco21589, w_eco21590, w_eco21591, w_eco21592, w_eco21593, w_eco21594, w_eco21595, w_eco21596, w_eco21597, w_eco21598, w_eco21599, w_eco21600, w_eco21601, w_eco21602, w_eco21603, w_eco21604, w_eco21605, w_eco21606, w_eco21607, w_eco21608, w_eco21609, w_eco21610, w_eco21611, w_eco21612, w_eco21613, w_eco21614, w_eco21615, w_eco21616, w_eco21617, w_eco21618, w_eco21619, w_eco21620, w_eco21621, w_eco21622, w_eco21623, w_eco21624, w_eco21625, w_eco21626, w_eco21627, w_eco21628, w_eco21629, w_eco21630, w_eco21631, w_eco21632, w_eco21633, w_eco21634, w_eco21635, w_eco21636, w_eco21637, w_eco21638, w_eco21639, w_eco21640, w_eco21641, w_eco21642, w_eco21643, w_eco21644, w_eco21645, w_eco21646, w_eco21647, w_eco21648, w_eco21649, w_eco21650, w_eco21651, w_eco21652, w_eco21653, w_eco21654, w_eco21655, w_eco21656, w_eco21657, w_eco21658, w_eco21659, w_eco21660, w_eco21661, w_eco21662, w_eco21663, w_eco21664, w_eco21665, w_eco21666, w_eco21667, w_eco21668, w_eco21669, w_eco21670, w_eco21671, w_eco21672, w_eco21673, w_eco21674, w_eco21675, w_eco21676, w_eco21677, w_eco21678, w_eco21679, w_eco21680, w_eco21681, w_eco21682, w_eco21683, w_eco21684, w_eco21685, w_eco21686, w_eco21687, w_eco21688, w_eco21689, w_eco21690, w_eco21691, w_eco21692, w_eco21693, w_eco21694, w_eco21695, w_eco21696, w_eco21697, w_eco21698, w_eco21699, w_eco21700, w_eco21701, w_eco21702, w_eco21703, w_eco21704, w_eco21705, w_eco21706, w_eco21707, w_eco21708, w_eco21709, w_eco21710, w_eco21711, w_eco21712, w_eco21713, w_eco21714, w_eco21715, w_eco21716, w_eco21717, w_eco21718, w_eco21719, w_eco21720, w_eco21721, w_eco21722, w_eco21723, w_eco21724, w_eco21725, w_eco21726, w_eco21727, w_eco21728, w_eco21729, w_eco21730, w_eco21731, w_eco21732, w_eco21733, w_eco21734, w_eco21735, w_eco21736, w_eco21737, w_eco21738, w_eco21739, w_eco21740, w_eco21741, w_eco21742, w_eco21743, w_eco21744, w_eco21745, w_eco21746, w_eco21747, w_eco21748, w_eco21749, w_eco21750, w_eco21751, w_eco21752, w_eco21753, w_eco21754, w_eco21755, w_eco21756, w_eco21757, w_eco21758, w_eco21759, w_eco21760, w_eco21761, w_eco21762, w_eco21763, w_eco21764, w_eco21765, w_eco21766, w_eco21767, w_eco21768, w_eco21769, w_eco21770, w_eco21771, w_eco21772, w_eco21773, w_eco21774, w_eco21775, w_eco21776, w_eco21777, w_eco21778, w_eco21779, w_eco21780, w_eco21781, w_eco21782, w_eco21783, w_eco21784, w_eco21785, w_eco21786, w_eco21787, w_eco21788, w_eco21789, w_eco21790, w_eco21791, w_eco21792, w_eco21793, w_eco21794, w_eco21795, w_eco21796, w_eco21797, w_eco21798, w_eco21799, w_eco21800, w_eco21801, w_eco21802, w_eco21803, w_eco21804, w_eco21805, w_eco21806, w_eco21807, w_eco21808, w_eco21809, w_eco21810, w_eco21811, w_eco21812, w_eco21813, w_eco21814, w_eco21815, w_eco21816, w_eco21817, w_eco21818, w_eco21819, w_eco21820, w_eco21821, w_eco21822, w_eco21823, w_eco21824, w_eco21825, w_eco21826, w_eco21827, w_eco21828, w_eco21829, w_eco21830, w_eco21831, w_eco21832, w_eco21833, w_eco21834, w_eco21835, w_eco21836, w_eco21837, w_eco21838, w_eco21839, w_eco21840, w_eco21841, w_eco21842, w_eco21843, w_eco21844, w_eco21845, w_eco21846, w_eco21847, w_eco21848, w_eco21849, w_eco21850, w_eco21851, w_eco21852, w_eco21853, w_eco21854, w_eco21855, w_eco21856, w_eco21857, w_eco21858, w_eco21859, w_eco21860, w_eco21861, w_eco21862, w_eco21863, w_eco21864, w_eco21865, w_eco21866, w_eco21867, w_eco21868, w_eco21869, w_eco21870, w_eco21871, w_eco21872, w_eco21873, w_eco21874, w_eco21875, w_eco21876, w_eco21877, w_eco21878, w_eco21879, w_eco21880, w_eco21881, w_eco21882, w_eco21883, w_eco21884, w_eco21885, w_eco21886, w_eco21887, w_eco21888, w_eco21889, w_eco21890, w_eco21891, w_eco21892, w_eco21893, w_eco21894, w_eco21895, w_eco21896, w_eco21897, w_eco21898, w_eco21899, w_eco21900, w_eco21901, w_eco21902, w_eco21903, w_eco21904, w_eco21905, w_eco21906, w_eco21907, w_eco21908, w_eco21909, w_eco21910, w_eco21911, w_eco21912, w_eco21913, w_eco21914, w_eco21915, w_eco21916, w_eco21917, w_eco21918, w_eco21919, w_eco21920, w_eco21921, w_eco21922, w_eco21923, w_eco21924, w_eco21925, w_eco21926, w_eco21927, w_eco21928, w_eco21929, w_eco21930, w_eco21931, w_eco21932, w_eco21933, w_eco21934, w_eco21935, w_eco21936, w_eco21937, w_eco21938, w_eco21939, w_eco21940, w_eco21941, w_eco21942, w_eco21943, w_eco21944, w_eco21945, w_eco21946, w_eco21947, w_eco21948, w_eco21949, w_eco21950, w_eco21951, w_eco21952, w_eco21953, w_eco21954, w_eco21955, w_eco21956, w_eco21957, w_eco21958, w_eco21959, w_eco21960, w_eco21961, w_eco21962, w_eco21963, w_eco21964, w_eco21965, w_eco21966, w_eco21967, w_eco21968, w_eco21969, w_eco21970, w_eco21971, w_eco21972, w_eco21973, w_eco21974, w_eco21975, w_eco21976, w_eco21977, w_eco21978, w_eco21979, w_eco21980, w_eco21981, w_eco21982, w_eco21983, w_eco21984, w_eco21985, w_eco21986, w_eco21987, w_eco21988, w_eco21989, w_eco21990, w_eco21991, w_eco21992, w_eco21993, w_eco21994, w_eco21995, w_eco21996, w_eco21997, w_eco21998, w_eco21999, w_eco22000, w_eco22001, w_eco22002, w_eco22003, w_eco22004, w_eco22005, w_eco22006, w_eco22007, w_eco22008, w_eco22009, w_eco22010, w_eco22011, w_eco22012, w_eco22013, w_eco22014, w_eco22015, w_eco22016, w_eco22017, w_eco22018, w_eco22019, w_eco22020, w_eco22021, w_eco22022, w_eco22023, w_eco22024, w_eco22025, w_eco22026, w_eco22027, w_eco22028, w_eco22029, w_eco22030, w_eco22031, w_eco22032, w_eco22033, w_eco22034, w_eco22035, w_eco22036, w_eco22037, w_eco22038, w_eco22039, w_eco22040, w_eco22041, w_eco22042, w_eco22043, w_eco22044, w_eco22045, w_eco22046, w_eco22047, w_eco22048, w_eco22049, w_eco22050, w_eco22051, w_eco22052, w_eco22053, w_eco22054, w_eco22055, w_eco22056, w_eco22057, w_eco22058, w_eco22059, w_eco22060, w_eco22061, w_eco22062, w_eco22063, w_eco22064, w_eco22065, w_eco22066, w_eco22067, w_eco22068, w_eco22069, w_eco22070, w_eco22071, w_eco22072, w_eco22073, w_eco22074, w_eco22075, w_eco22076, w_eco22077, w_eco22078, w_eco22079, w_eco22080, w_eco22081, w_eco22082, w_eco22083, w_eco22084, w_eco22085, w_eco22086, w_eco22087, w_eco22088, w_eco22089, w_eco22090, w_eco22091, w_eco22092, w_eco22093, w_eco22094, w_eco22095, w_eco22096, w_eco22097, w_eco22098, w_eco22099, w_eco22100, w_eco22101, w_eco22102, w_eco22103, w_eco22104, w_eco22105, w_eco22106, w_eco22107, w_eco22108, w_eco22109, w_eco22110, w_eco22111, w_eco22112, w_eco22113, w_eco22114, w_eco22115, w_eco22116, w_eco22117, w_eco22118, w_eco22119, w_eco22120, w_eco22121, w_eco22122, w_eco22123, w_eco22124, w_eco22125, w_eco22126, w_eco22127, w_eco22128, w_eco22129, w_eco22130, w_eco22131, w_eco22132, w_eco22133, w_eco22134, w_eco22135, w_eco22136, w_eco22137, w_eco22138, w_eco22139, w_eco22140, w_eco22141, w_eco22142, w_eco22143, w_eco22144, w_eco22145, w_eco22146, w_eco22147, w_eco22148, w_eco22149, w_eco22150, w_eco22151, w_eco22152, w_eco22153, w_eco22154, w_eco22155, w_eco22156, w_eco22157, w_eco22158, w_eco22159, w_eco22160, w_eco22161, w_eco22162, w_eco22163, w_eco22164, w_eco22165, w_eco22166, w_eco22167, w_eco22168, w_eco22169, w_eco22170, w_eco22171, w_eco22172, w_eco22173, w_eco22174, w_eco22175, w_eco22176, w_eco22177, w_eco22178, w_eco22179, w_eco22180, w_eco22181, w_eco22182, w_eco22183, w_eco22184, w_eco22185, w_eco22186, w_eco22187, w_eco22188, w_eco22189, w_eco22190, w_eco22191, w_eco22192, w_eco22193, w_eco22194, w_eco22195, w_eco22196, w_eco22197, w_eco22198, w_eco22199, w_eco22200, w_eco22201, w_eco22202, w_eco22203, w_eco22204, w_eco22205, w_eco22206, w_eco22207, w_eco22208, w_eco22209, w_eco22210, w_eco22211, w_eco22212, w_eco22213, w_eco22214, w_eco22215, w_eco22216, w_eco22217, w_eco22218, w_eco22219, w_eco22220, w_eco22221, w_eco22222, w_eco22223, w_eco22224, w_eco22225, w_eco22226, w_eco22227, w_eco22228, w_eco22229, w_eco22230, w_eco22231, w_eco22232, w_eco22233, w_eco22234, w_eco22235, w_eco22236, w_eco22237, w_eco22238, w_eco22239, w_eco22240, w_eco22241, w_eco22242, w_eco22243, w_eco22244, w_eco22245, w_eco22246, w_eco22247, w_eco22248, w_eco22249, w_eco22250, w_eco22251, w_eco22252, w_eco22253, w_eco22254, w_eco22255, w_eco22256, w_eco22257, w_eco22258, w_eco22259, w_eco22260, w_eco22261, w_eco22262, w_eco22263, w_eco22264, w_eco22265, w_eco22266, w_eco22267, w_eco22268, w_eco22269, w_eco22270, w_eco22271, w_eco22272, w_eco22273, w_eco22274, w_eco22275, w_eco22276, w_eco22277, w_eco22278, w_eco22279, w_eco22280, w_eco22281, w_eco22282, w_eco22283, w_eco22284, w_eco22285, w_eco22286, w_eco22287, w_eco22288, w_eco22289, w_eco22290, w_eco22291, w_eco22292, w_eco22293, w_eco22294, w_eco22295, w_eco22296, w_eco22297, w_eco22298, w_eco22299, w_eco22300, w_eco22301, w_eco22302, w_eco22303, w_eco22304, w_eco22305, w_eco22306, w_eco22307, w_eco22308, w_eco22309, w_eco22310, w_eco22311, w_eco22312, w_eco22313, w_eco22314, w_eco22315, w_eco22316, w_eco22317, w_eco22318, w_eco22319, w_eco22320, w_eco22321, w_eco22322, w_eco22323, w_eco22324, w_eco22325, w_eco22326, w_eco22327, w_eco22328, w_eco22329, w_eco22330, w_eco22331, w_eco22332, w_eco22333, w_eco22334, w_eco22335, w_eco22336, w_eco22337, w_eco22338, w_eco22339, w_eco22340, w_eco22341, w_eco22342, w_eco22343, w_eco22344, w_eco22345, w_eco22346, w_eco22347, w_eco22348, w_eco22349, w_eco22350, w_eco22351, w_eco22352, w_eco22353, w_eco22354, w_eco22355, w_eco22356, w_eco22357, w_eco22358, w_eco22359, w_eco22360, w_eco22361, w_eco22362, w_eco22363, w_eco22364, w_eco22365, w_eco22366, w_eco22367, w_eco22368, w_eco22369, w_eco22370, w_eco22371, w_eco22372, w_eco22373, w_eco22374, w_eco22375, w_eco22376, w_eco22377, w_eco22378, w_eco22379, w_eco22380, w_eco22381, w_eco22382, w_eco22383, w_eco22384, w_eco22385, w_eco22386, w_eco22387, w_eco22388, w_eco22389, w_eco22390, w_eco22391, w_eco22392, w_eco22393, w_eco22394, w_eco22395, w_eco22396, w_eco22397, w_eco22398, w_eco22399, w_eco22400, w_eco22401, w_eco22402, w_eco22403, w_eco22404, w_eco22405, w_eco22406, w_eco22407, w_eco22408, w_eco22409, w_eco22410, w_eco22411, w_eco22412, w_eco22413, w_eco22414, w_eco22415, w_eco22416, w_eco22417, w_eco22418, w_eco22419, w_eco22420, w_eco22421, w_eco22422, w_eco22423, w_eco22424, w_eco22425, w_eco22426, w_eco22427, w_eco22428, w_eco22429, w_eco22430, w_eco22431, w_eco22432, w_eco22433, w_eco22434, w_eco22435, w_eco22436, w_eco22437, w_eco22438, w_eco22439, w_eco22440, w_eco22441, w_eco22442, w_eco22443, w_eco22444, w_eco22445, w_eco22446, w_eco22447, w_eco22448, w_eco22449, w_eco22450, w_eco22451, w_eco22452, w_eco22453, w_eco22454, w_eco22455, w_eco22456, w_eco22457, w_eco22458, w_eco22459, w_eco22460, w_eco22461, w_eco22462, w_eco22463, w_eco22464, w_eco22465, w_eco22466, w_eco22467, w_eco22468, w_eco22469, w_eco22470, w_eco22471, w_eco22472, w_eco22473, w_eco22474, w_eco22475, w_eco22476, w_eco22477, w_eco22478, w_eco22479, w_eco22480, w_eco22481, w_eco22482, w_eco22483, w_eco22484, w_eco22485, w_eco22486, w_eco22487, w_eco22488, w_eco22489, w_eco22490, w_eco22491, w_eco22492, w_eco22493, w_eco22494, w_eco22495, w_eco22496, w_eco22497, w_eco22498, w_eco22499, w_eco22500, w_eco22501, w_eco22502, w_eco22503, w_eco22504, w_eco22505, w_eco22506, w_eco22507, w_eco22508, w_eco22509, w_eco22510, w_eco22511, w_eco22512, w_eco22513, w_eco22514, w_eco22515, w_eco22516, w_eco22517, w_eco22518, w_eco22519, w_eco22520, w_eco22521, w_eco22522, w_eco22523, w_eco22524, w_eco22525, w_eco22526, w_eco22527, w_eco22528, w_eco22529, w_eco22530, w_eco22531, w_eco22532, w_eco22533, w_eco22534, w_eco22535, w_eco22536, w_eco22537, w_eco22538, w_eco22539, w_eco22540, w_eco22541, w_eco22542, w_eco22543, w_eco22544, w_eco22545, w_eco22546, w_eco22547, w_eco22548, w_eco22549, w_eco22550, w_eco22551, w_eco22552, w_eco22553, w_eco22554, w_eco22555, w_eco22556, w_eco22557, w_eco22558, w_eco22559, w_eco22560, w_eco22561, w_eco22562, w_eco22563, w_eco22564, w_eco22565, w_eco22566, w_eco22567, w_eco22568, w_eco22569, w_eco22570, w_eco22571, w_eco22572, w_eco22573, w_eco22574, w_eco22575, w_eco22576, w_eco22577, w_eco22578, w_eco22579, w_eco22580, w_eco22581, w_eco22582, w_eco22583, w_eco22584, w_eco22585, w_eco22586, w_eco22587, w_eco22588, w_eco22589, w_eco22590, w_eco22591, w_eco22592, w_eco22593, w_eco22594, w_eco22595, w_eco22596, w_eco22597, w_eco22598, w_eco22599, w_eco22600, w_eco22601, w_eco22602, w_eco22603, w_eco22604, w_eco22605, w_eco22606, w_eco22607, w_eco22608, w_eco22609, w_eco22610, w_eco22611, w_eco22612, w_eco22613, w_eco22614, w_eco22615, w_eco22616, w_eco22617, w_eco22618, w_eco22619, w_eco22620, w_eco22621, w_eco22622, w_eco22623, w_eco22624, w_eco22625, w_eco22626, w_eco22627, w_eco22628, w_eco22629, w_eco22630, w_eco22631, w_eco22632, w_eco22633, w_eco22634, w_eco22635, w_eco22636, w_eco22637, w_eco22638, w_eco22639, w_eco22640, w_eco22641, w_eco22642, w_eco22643, w_eco22644, w_eco22645, w_eco22646, w_eco22647, w_eco22648, w_eco22649, w_eco22650, w_eco22651, w_eco22652, w_eco22653, w_eco22654, w_eco22655, w_eco22656, w_eco22657, w_eco22658, w_eco22659, w_eco22660, w_eco22661, w_eco22662, w_eco22663, w_eco22664, w_eco22665, w_eco22666, w_eco22667, w_eco22668, w_eco22669, w_eco22670, w_eco22671, w_eco22672, w_eco22673, w_eco22674, w_eco22675, w_eco22676, w_eco22677, w_eco22678, w_eco22679, w_eco22680, w_eco22681, w_eco22682, w_eco22683, w_eco22684, w_eco22685, w_eco22686, w_eco22687, w_eco22688, w_eco22689, w_eco22690, w_eco22691, w_eco22692, w_eco22693, w_eco22694, w_eco22695, w_eco22696, w_eco22697, w_eco22698, w_eco22699, w_eco22700, w_eco22701, w_eco22702, w_eco22703, w_eco22704, w_eco22705, w_eco22706, w_eco22707, w_eco22708, w_eco22709, w_eco22710, w_eco22711, w_eco22712, w_eco22713, w_eco22714, w_eco22715, w_eco22716, w_eco22717, w_eco22718, w_eco22719, w_eco22720, w_eco22721, w_eco22722, w_eco22723, w_eco22724, w_eco22725, w_eco22726, w_eco22727, w_eco22728, w_eco22729, w_eco22730, w_eco22731, w_eco22732, w_eco22733, w_eco22734, w_eco22735, w_eco22736, w_eco22737, w_eco22738, w_eco22739, w_eco22740, w_eco22741, w_eco22742, w_eco22743, w_eco22744, w_eco22745, w_eco22746, w_eco22747, w_eco22748, w_eco22749, w_eco22750, w_eco22751, w_eco22752, w_eco22753, w_eco22754, w_eco22755, w_eco22756, w_eco22757, w_eco22758, w_eco22759, w_eco22760, w_eco22761, w_eco22762, w_eco22763, w_eco22764, w_eco22765, w_eco22766, w_eco22767, w_eco22768, w_eco22769, w_eco22770, w_eco22771, w_eco22772, w_eco22773, w_eco22774, w_eco22775, w_eco22776, w_eco22777, w_eco22778, w_eco22779, w_eco22780, w_eco22781, w_eco22782, w_eco22783, w_eco22784, w_eco22785, w_eco22786, w_eco22787, w_eco22788, w_eco22789, w_eco22790, w_eco22791, w_eco22792, w_eco22793, w_eco22794, w_eco22795, w_eco22796, w_eco22797, w_eco22798, w_eco22799, w_eco22800, w_eco22801, w_eco22802, w_eco22803, w_eco22804, w_eco22805, w_eco22806, w_eco22807, w_eco22808, w_eco22809, w_eco22810, w_eco22811, w_eco22812, w_eco22813, w_eco22814, w_eco22815, w_eco22816, w_eco22817, w_eco22818, w_eco22819, w_eco22820, w_eco22821, w_eco22822, w_eco22823, w_eco22824, w_eco22825, w_eco22826, w_eco22827, w_eco22828, w_eco22829, w_eco22830, w_eco22831, w_eco22832, w_eco22833, w_eco22834, w_eco22835, w_eco22836, w_eco22837, w_eco22838, w_eco22839, w_eco22840, w_eco22841, w_eco22842, w_eco22843, w_eco22844, w_eco22845, w_eco22846, w_eco22847, w_eco22848, w_eco22849, w_eco22850, w_eco22851, w_eco22852, w_eco22853, w_eco22854, w_eco22855, w_eco22856, w_eco22857, w_eco22858, w_eco22859, w_eco22860, w_eco22861, w_eco22862, w_eco22863, w_eco22864, w_eco22865, w_eco22866, w_eco22867, w_eco22868, w_eco22869, w_eco22870, w_eco22871, w_eco22872, w_eco22873, w_eco22874, w_eco22875, w_eco22876, w_eco22877, w_eco22878, w_eco22879, w_eco22880, w_eco22881, w_eco22882, w_eco22883, w_eco22884, w_eco22885, w_eco22886, w_eco22887, w_eco22888, w_eco22889, w_eco22890, w_eco22891, w_eco22892, w_eco22893, w_eco22894, w_eco22895, w_eco22896, w_eco22897, w_eco22898, w_eco22899, w_eco22900, w_eco22901, w_eco22902, w_eco22903, w_eco22904, w_eco22905, w_eco22906, w_eco22907, w_eco22908, w_eco22909, w_eco22910, w_eco22911, w_eco22912, w_eco22913, w_eco22914, w_eco22915, w_eco22916, w_eco22917, w_eco22918, w_eco22919, w_eco22920, w_eco22921, w_eco22922, w_eco22923, w_eco22924, w_eco22925, w_eco22926, w_eco22927, w_eco22928, w_eco22929, w_eco22930, w_eco22931, w_eco22932, w_eco22933, w_eco22934, w_eco22935, w_eco22936, w_eco22937, w_eco22938, w_eco22939, w_eco22940, w_eco22941, w_eco22942, w_eco22943, w_eco22944, w_eco22945, w_eco22946, w_eco22947, w_eco22948, w_eco22949, w_eco22950, w_eco22951, w_eco22952, w_eco22953, w_eco22954, w_eco22955, w_eco22956, w_eco22957, w_eco22958, w_eco22959, w_eco22960, w_eco22961, w_eco22962, w_eco22963, w_eco22964, w_eco22965, w_eco22966, w_eco22967, w_eco22968, w_eco22969, w_eco22970, w_eco22971, w_eco22972, w_eco22973, w_eco22974, w_eco22975, w_eco22976, w_eco22977, w_eco22978, w_eco22979, w_eco22980, w_eco22981, w_eco22982, w_eco22983, w_eco22984, w_eco22985, w_eco22986, w_eco22987, w_eco22988, w_eco22989, w_eco22990, w_eco22991, w_eco22992, w_eco22993, w_eco22994, w_eco22995, w_eco22996, w_eco22997, w_eco22998, w_eco22999, w_eco23000, w_eco23001, w_eco23002, w_eco23003, w_eco23004, w_eco23005, w_eco23006, w_eco23007, w_eco23008, w_eco23009, w_eco23010, w_eco23011, w_eco23012, w_eco23013, w_eco23014, w_eco23015, w_eco23016, w_eco23017, w_eco23018, w_eco23019, w_eco23020, w_eco23021, w_eco23022, w_eco23023, w_eco23024, w_eco23025, w_eco23026, w_eco23027, w_eco23028, w_eco23029, w_eco23030, w_eco23031, w_eco23032, w_eco23033, w_eco23034, w_eco23035, w_eco23036, w_eco23037, w_eco23038, w_eco23039, w_eco23040, w_eco23041, w_eco23042, w_eco23043, w_eco23044, w_eco23045, w_eco23046, w_eco23047, w_eco23048, w_eco23049, w_eco23050, w_eco23051, w_eco23052, w_eco23053, w_eco23054, w_eco23055, w_eco23056, w_eco23057, w_eco23058, w_eco23059, w_eco23060, w_eco23061, w_eco23062, w_eco23063, w_eco23064, w_eco23065, w_eco23066, w_eco23067, w_eco23068, w_eco23069, w_eco23070, w_eco23071, w_eco23072, w_eco23073, w_eco23074, w_eco23075, w_eco23076, w_eco23077, w_eco23078, w_eco23079, w_eco23080, w_eco23081, w_eco23082, w_eco23083, w_eco23084, w_eco23085, w_eco23086, w_eco23087, w_eco23088, w_eco23089, w_eco23090, w_eco23091, w_eco23092, w_eco23093, w_eco23094, w_eco23095, w_eco23096, w_eco23097, w_eco23098, w_eco23099, w_eco23100, w_eco23101, w_eco23102, w_eco23103, w_eco23104, w_eco23105, w_eco23106, w_eco23107, w_eco23108, w_eco23109, w_eco23110, w_eco23111, w_eco23112, w_eco23113, w_eco23114, w_eco23115, w_eco23116, w_eco23117, w_eco23118, w_eco23119, w_eco23120, w_eco23121, w_eco23122, w_eco23123, w_eco23124, w_eco23125, w_eco23126, w_eco23127, w_eco23128, w_eco23129, w_eco23130, w_eco23131, w_eco23132, w_eco23133, w_eco23134, w_eco23135, w_eco23136, w_eco23137, w_eco23138, w_eco23139, w_eco23140, w_eco23141, w_eco23142, w_eco23143, w_eco23144, w_eco23145, w_eco23146, w_eco23147, w_eco23148, w_eco23149, w_eco23150, w_eco23151, w_eco23152, w_eco23153, w_eco23154, w_eco23155, w_eco23156, w_eco23157, w_eco23158, w_eco23159, w_eco23160, w_eco23161, w_eco23162, w_eco23163, w_eco23164, w_eco23165, w_eco23166, w_eco23167, w_eco23168, w_eco23169, w_eco23170, w_eco23171, w_eco23172, w_eco23173, w_eco23174, w_eco23175, w_eco23176, w_eco23177, w_eco23178, w_eco23179, w_eco23180, w_eco23181, w_eco23182, w_eco23183, w_eco23184, w_eco23185, w_eco23186, w_eco23187, w_eco23188, w_eco23189, w_eco23190, w_eco23191, w_eco23192, w_eco23193, w_eco23194, w_eco23195, w_eco23196, w_eco23197, w_eco23198, w_eco23199, w_eco23200, w_eco23201, w_eco23202, w_eco23203, w_eco23204, w_eco23205, w_eco23206, w_eco23207, w_eco23208, w_eco23209, w_eco23210, w_eco23211, w_eco23212, w_eco23213, w_eco23214, w_eco23215, w_eco23216, w_eco23217, w_eco23218, w_eco23219, w_eco23220, w_eco23221, w_eco23222, w_eco23223, w_eco23224, w_eco23225, w_eco23226, w_eco23227, w_eco23228, w_eco23229, w_eco23230, w_eco23231, w_eco23232, w_eco23233, w_eco23234, w_eco23235, w_eco23236, w_eco23237, w_eco23238, w_eco23239, w_eco23240, w_eco23241, w_eco23242, w_eco23243, w_eco23244, w_eco23245, w_eco23246, w_eco23247, w_eco23248, w_eco23249, w_eco23250, w_eco23251, w_eco23252, w_eco23253, w_eco23254, w_eco23255, w_eco23256, w_eco23257, w_eco23258, w_eco23259, w_eco23260, w_eco23261, w_eco23262, w_eco23263, w_eco23264, w_eco23265, w_eco23266, w_eco23267, w_eco23268, w_eco23269, w_eco23270, w_eco23271, w_eco23272, w_eco23273, w_eco23274, w_eco23275, w_eco23276, w_eco23277, w_eco23278, w_eco23279, w_eco23280, w_eco23281, w_eco23282, w_eco23283, w_eco23284, w_eco23285, w_eco23286, w_eco23287, w_eco23288, w_eco23289, w_eco23290, w_eco23291, w_eco23292, w_eco23293, w_eco23294, w_eco23295, w_eco23296, w_eco23297, w_eco23298, w_eco23299, w_eco23300, w_eco23301, w_eco23302, w_eco23303, w_eco23304, w_eco23305, w_eco23306, w_eco23307, w_eco23308, w_eco23309, w_eco23310, w_eco23311, w_eco23312, w_eco23313, w_eco23314, w_eco23315, w_eco23316, w_eco23317, w_eco23318, w_eco23319, w_eco23320, w_eco23321, w_eco23322, w_eco23323, w_eco23324, w_eco23325, w_eco23326, w_eco23327, w_eco23328, w_eco23329, w_eco23330, w_eco23331, w_eco23332, w_eco23333, w_eco23334, w_eco23335, w_eco23336, w_eco23337, w_eco23338, w_eco23339, w_eco23340, w_eco23341, w_eco23342, w_eco23343, w_eco23344, w_eco23345, w_eco23346, w_eco23347, w_eco23348, w_eco23349, w_eco23350, w_eco23351, w_eco23352, w_eco23353, w_eco23354, w_eco23355, w_eco23356, w_eco23357, w_eco23358, w_eco23359, w_eco23360, w_eco23361, w_eco23362, w_eco23363, w_eco23364, w_eco23365, w_eco23366, w_eco23367, w_eco23368, w_eco23369, w_eco23370, w_eco23371, w_eco23372, w_eco23373, w_eco23374, w_eco23375, w_eco23376, w_eco23377, w_eco23378, w_eco23379, w_eco23380, w_eco23381, w_eco23382, w_eco23383, w_eco23384, w_eco23385, w_eco23386, w_eco23387, w_eco23388, w_eco23389, w_eco23390, w_eco23391, w_eco23392, w_eco23393, w_eco23394, w_eco23395, w_eco23396, w_eco23397, w_eco23398, w_eco23399, w_eco23400, w_eco23401, w_eco23402, w_eco23403, w_eco23404, w_eco23405, w_eco23406, w_eco23407, w_eco23408, w_eco23409, w_eco23410, w_eco23411, w_eco23412, w_eco23413, w_eco23414, w_eco23415, w_eco23416, w_eco23417, w_eco23418, w_eco23419, w_eco23420, w_eco23421, w_eco23422, w_eco23423, w_eco23424, w_eco23425, w_eco23426, w_eco23427, w_eco23428, w_eco23429, w_eco23430, w_eco23431, w_eco23432, w_eco23433, w_eco23434, w_eco23435, w_eco23436, w_eco23437, w_eco23438, w_eco23439, w_eco23440, w_eco23441, w_eco23442, w_eco23443, w_eco23444, w_eco23445, w_eco23446, w_eco23447, w_eco23448, w_eco23449, w_eco23450, w_eco23451, w_eco23452, w_eco23453, w_eco23454, w_eco23455, w_eco23456, w_eco23457, w_eco23458, w_eco23459, w_eco23460, w_eco23461, w_eco23462, w_eco23463, w_eco23464, w_eco23465, w_eco23466, w_eco23467, w_eco23468, w_eco23469, w_eco23470, w_eco23471, w_eco23472, w_eco23473, w_eco23474, w_eco23475, w_eco23476, w_eco23477, w_eco23478, w_eco23479, w_eco23480, w_eco23481, w_eco23482, w_eco23483, w_eco23484, w_eco23485, w_eco23486, w_eco23487, w_eco23488, w_eco23489, w_eco23490, w_eco23491, w_eco23492, w_eco23493, w_eco23494, w_eco23495, w_eco23496, w_eco23497, w_eco23498, w_eco23499, w_eco23500, w_eco23501, w_eco23502, w_eco23503, w_eco23504, w_eco23505, w_eco23506, w_eco23507, w_eco23508, w_eco23509, w_eco23510, w_eco23511, w_eco23512, w_eco23513, w_eco23514, w_eco23515, w_eco23516, w_eco23517, w_eco23518, w_eco23519, w_eco23520, w_eco23521, w_eco23522, w_eco23523, w_eco23524, w_eco23525, w_eco23526, w_eco23527, w_eco23528, w_eco23529, w_eco23530, w_eco23531, w_eco23532, w_eco23533, w_eco23534, w_eco23535, w_eco23536, w_eco23537, w_eco23538, w_eco23539, w_eco23540, w_eco23541, w_eco23542, w_eco23543, w_eco23544, w_eco23545, w_eco23546, w_eco23547, w_eco23548, w_eco23549, w_eco23550, w_eco23551, w_eco23552, w_eco23553, w_eco23554, w_eco23555, w_eco23556, w_eco23557, w_eco23558, w_eco23559, w_eco23560, w_eco23561, w_eco23562, w_eco23563, w_eco23564, w_eco23565, w_eco23566, w_eco23567, w_eco23568, w_eco23569, w_eco23570, w_eco23571, w_eco23572, w_eco23573, w_eco23574, w_eco23575, w_eco23576, w_eco23577, w_eco23578, w_eco23579, w_eco23580, w_eco23581, w_eco23582, w_eco23583, w_eco23584, w_eco23585, w_eco23586, w_eco23587, w_eco23588, w_eco23589, w_eco23590, w_eco23591, w_eco23592, w_eco23593, w_eco23594, w_eco23595, w_eco23596, w_eco23597, w_eco23598, w_eco23599, w_eco23600, w_eco23601, w_eco23602, w_eco23603, w_eco23604, w_eco23605, w_eco23606, w_eco23607, w_eco23608, w_eco23609, w_eco23610, w_eco23611, w_eco23612, w_eco23613, w_eco23614, w_eco23615, w_eco23616, w_eco23617, w_eco23618, w_eco23619, w_eco23620, w_eco23621, w_eco23622, w_eco23623, w_eco23624, w_eco23625, w_eco23626, w_eco23627, w_eco23628, w_eco23629, w_eco23630, w_eco23631, w_eco23632, w_eco23633, w_eco23634, w_eco23635, w_eco23636, w_eco23637, w_eco23638, w_eco23639, w_eco23640, w_eco23641, w_eco23642, w_eco23643, w_eco23644, w_eco23645, w_eco23646, w_eco23647, w_eco23648, w_eco23649, w_eco23650, w_eco23651, w_eco23652, w_eco23653, w_eco23654, w_eco23655, w_eco23656, w_eco23657, w_eco23658, w_eco23659, w_eco23660, w_eco23661, w_eco23662, w_eco23663, w_eco23664, w_eco23665, w_eco23666, w_eco23667, w_eco23668, w_eco23669, w_eco23670, w_eco23671, w_eco23672, w_eco23673, w_eco23674, w_eco23675, w_eco23676, w_eco23677, w_eco23678, w_eco23679, w_eco23680, w_eco23681, w_eco23682, w_eco23683, w_eco23684, w_eco23685, w_eco23686, w_eco23687, w_eco23688, w_eco23689, w_eco23690, w_eco23691, w_eco23692, w_eco23693, w_eco23694, w_eco23695, w_eco23696, w_eco23697, w_eco23698, w_eco23699, w_eco23700, w_eco23701, w_eco23702, w_eco23703, w_eco23704, w_eco23705, w_eco23706, w_eco23707, w_eco23708, w_eco23709, w_eco23710, w_eco23711, w_eco23712, w_eco23713, w_eco23714, w_eco23715, w_eco23716, w_eco23717, w_eco23718, w_eco23719, w_eco23720, w_eco23721, w_eco23722, w_eco23723, w_eco23724, w_eco23725, w_eco23726, w_eco23727, w_eco23728, w_eco23729, w_eco23730, w_eco23731, w_eco23732, w_eco23733, w_eco23734, w_eco23735, w_eco23736, w_eco23737, w_eco23738, w_eco23739, w_eco23740, w_eco23741, w_eco23742, w_eco23743, w_eco23744, w_eco23745, w_eco23746, w_eco23747, w_eco23748, w_eco23749, w_eco23750, w_eco23751, w_eco23752, w_eco23753, w_eco23754, w_eco23755, w_eco23756, w_eco23757, w_eco23758, w_eco23759, w_eco23760, w_eco23761, w_eco23762, w_eco23763, w_eco23764, w_eco23765, w_eco23766, w_eco23767, w_eco23768, w_eco23769, w_eco23770, w_eco23771, w_eco23772, w_eco23773, w_eco23774, w_eco23775, w_eco23776, w_eco23777, w_eco23778, w_eco23779, w_eco23780, w_eco23781, w_eco23782, w_eco23783, w_eco23784, w_eco23785, w_eco23786, w_eco23787, w_eco23788, w_eco23789, w_eco23790, w_eco23791, w_eco23792, w_eco23793, w_eco23794, w_eco23795, w_eco23796, w_eco23797, w_eco23798, w_eco23799, w_eco23800, w_eco23801, w_eco23802, w_eco23803, w_eco23804, w_eco23805, w_eco23806, w_eco23807, w_eco23808, w_eco23809, w_eco23810, w_eco23811, w_eco23812, w_eco23813, w_eco23814, w_eco23815, w_eco23816, w_eco23817, w_eco23818, w_eco23819, w_eco23820, w_eco23821, w_eco23822, w_eco23823, w_eco23824, w_eco23825, w_eco23826, w_eco23827, w_eco23828, w_eco23829, w_eco23830, w_eco23831, w_eco23832, w_eco23833, w_eco23834, w_eco23835, w_eco23836, w_eco23837, w_eco23838, w_eco23839, w_eco23840, w_eco23841, w_eco23842, w_eco23843, w_eco23844, w_eco23845, w_eco23846, w_eco23847, w_eco23848, w_eco23849, w_eco23850, w_eco23851, w_eco23852, w_eco23853, w_eco23854, w_eco23855, w_eco23856, w_eco23857, w_eco23858, w_eco23859, w_eco23860, w_eco23861, w_eco23862, w_eco23863, w_eco23864, w_eco23865, w_eco23866, w_eco23867, w_eco23868, w_eco23869, w_eco23870, w_eco23871, w_eco23872, w_eco23873, w_eco23874, w_eco23875, w_eco23876, w_eco23877, w_eco23878, w_eco23879, w_eco23880, w_eco23881, w_eco23882, w_eco23883, w_eco23884, w_eco23885, w_eco23886, w_eco23887, w_eco23888, w_eco23889, w_eco23890, w_eco23891, w_eco23892, w_eco23893, w_eco23894, w_eco23895, w_eco23896, w_eco23897, w_eco23898, w_eco23899, w_eco23900, w_eco23901, w_eco23902, w_eco23903, w_eco23904, w_eco23905, w_eco23906, w_eco23907, w_eco23908, w_eco23909, w_eco23910, w_eco23911, w_eco23912, w_eco23913, w_eco23914, w_eco23915, w_eco23916, w_eco23917, w_eco23918, w_eco23919, w_eco23920, w_eco23921, w_eco23922, w_eco23923, w_eco23924, w_eco23925, w_eco23926, w_eco23927, w_eco23928, w_eco23929, w_eco23930, w_eco23931, w_eco23932, w_eco23933, w_eco23934, w_eco23935, w_eco23936, w_eco23937, w_eco23938, w_eco23939, w_eco23940, w_eco23941, w_eco23942, w_eco23943, w_eco23944, w_eco23945, w_eco23946, w_eco23947, w_eco23948, w_eco23949, w_eco23950, w_eco23951, w_eco23952, w_eco23953, w_eco23954, w_eco23955, w_eco23956, w_eco23957, w_eco23958, w_eco23959, w_eco23960, w_eco23961, w_eco23962, w_eco23963, w_eco23964, w_eco23965, w_eco23966, w_eco23967, w_eco23968, w_eco23969, w_eco23970, w_eco23971, w_eco23972, w_eco23973, w_eco23974, w_eco23975, w_eco23976, w_eco23977, w_eco23978, w_eco23979, w_eco23980, w_eco23981, w_eco23982, w_eco23983, w_eco23984, w_eco23985, w_eco23986, w_eco23987, w_eco23988, w_eco23989, w_eco23990, w_eco23991, w_eco23992, w_eco23993, w_eco23994, w_eco23995, w_eco23996, w_eco23997, w_eco23998, w_eco23999, w_eco24000, w_eco24001, w_eco24002, w_eco24003, w_eco24004, w_eco24005, w_eco24006, w_eco24007, w_eco24008, w_eco24009, w_eco24010, w_eco24011, w_eco24012, w_eco24013, w_eco24014, w_eco24015, w_eco24016, w_eco24017, w_eco24018, w_eco24019, w_eco24020, w_eco24021, w_eco24022, w_eco24023, w_eco24024, w_eco24025, w_eco24026, w_eco24027, w_eco24028, w_eco24029, w_eco24030, w_eco24031, w_eco24032, w_eco24033, w_eco24034, w_eco24035, w_eco24036, w_eco24037, w_eco24038, w_eco24039, w_eco24040, w_eco24041, w_eco24042, w_eco24043, w_eco24044, w_eco24045, w_eco24046, w_eco24047, w_eco24048, w_eco24049, w_eco24050, w_eco24051, w_eco24052, w_eco24053, w_eco24054, w_eco24055, w_eco24056, w_eco24057, w_eco24058, w_eco24059, w_eco24060, w_eco24061, w_eco24062, w_eco24063, w_eco24064, w_eco24065, w_eco24066, w_eco24067, w_eco24068, w_eco24069, w_eco24070, w_eco24071, w_eco24072, w_eco24073, w_eco24074, w_eco24075, w_eco24076, w_eco24077, w_eco24078, w_eco24079, w_eco24080, w_eco24081, w_eco24082, w_eco24083, w_eco24084, w_eco24085, w_eco24086, w_eco24087, w_eco24088, w_eco24089, w_eco24090, w_eco24091, w_eco24092, w_eco24093, w_eco24094, w_eco24095, w_eco24096, w_eco24097, w_eco24098, w_eco24099, w_eco24100, w_eco24101, w_eco24102, w_eco24103, w_eco24104, w_eco24105, w_eco24106, w_eco24107, w_eco24108, w_eco24109, w_eco24110, w_eco24111, w_eco24112, w_eco24113, w_eco24114, w_eco24115, w_eco24116, w_eco24117, w_eco24118, w_eco24119, w_eco24120, w_eco24121, w_eco24122, w_eco24123, w_eco24124, w_eco24125, w_eco24126, w_eco24127, w_eco24128, w_eco24129, w_eco24130, w_eco24131, w_eco24132, w_eco24133, w_eco24134, w_eco24135, w_eco24136, w_eco24137, w_eco24138, w_eco24139, w_eco24140, w_eco24141, w_eco24142, w_eco24143, w_eco24144, w_eco24145, w_eco24146, w_eco24147, w_eco24148, w_eco24149, w_eco24150, w_eco24151, w_eco24152, w_eco24153, w_eco24154, w_eco24155, w_eco24156, w_eco24157, w_eco24158, w_eco24159, w_eco24160, w_eco24161, w_eco24162, w_eco24163, w_eco24164, w_eco24165, w_eco24166, w_eco24167, w_eco24168, w_eco24169, w_eco24170, w_eco24171, w_eco24172, w_eco24173, w_eco24174, w_eco24175, w_eco24176, w_eco24177, w_eco24178, w_eco24179, w_eco24180, w_eco24181, w_eco24182, w_eco24183, w_eco24184, w_eco24185, w_eco24186, w_eco24187, w_eco24188, w_eco24189, w_eco24190, w_eco24191, w_eco24192, w_eco24193, w_eco24194, w_eco24195, w_eco24196, w_eco24197, w_eco24198, w_eco24199, w_eco24200, w_eco24201, w_eco24202, w_eco24203, w_eco24204, w_eco24205, w_eco24206, w_eco24207, w_eco24208, w_eco24209, w_eco24210, w_eco24211, w_eco24212, w_eco24213, w_eco24214, w_eco24215, w_eco24216, w_eco24217, w_eco24218, w_eco24219, w_eco24220, w_eco24221, w_eco24222, w_eco24223, w_eco24224, w_eco24225, w_eco24226, w_eco24227, w_eco24228, w_eco24229, w_eco24230, w_eco24231, w_eco24232, w_eco24233, w_eco24234, w_eco24235, w_eco24236, w_eco24237, w_eco24238, w_eco24239, w_eco24240, w_eco24241, w_eco24242, w_eco24243, w_eco24244, w_eco24245, w_eco24246, w_eco24247, w_eco24248, w_eco24249, w_eco24250, w_eco24251, w_eco24252, w_eco24253, w_eco24254, w_eco24255, w_eco24256, w_eco24257, w_eco24258, w_eco24259, w_eco24260, w_eco24261, w_eco24262, w_eco24263, w_eco24264, w_eco24265, w_eco24266, w_eco24267, w_eco24268, w_eco24269, w_eco24270, w_eco24271, w_eco24272, w_eco24273, w_eco24274, w_eco24275, w_eco24276, w_eco24277, w_eco24278, w_eco24279, w_eco24280, w_eco24281, w_eco24282, w_eco24283, w_eco24284, w_eco24285, w_eco24286, w_eco24287, w_eco24288, w_eco24289, w_eco24290, w_eco24291, w_eco24292, w_eco24293, w_eco24294, w_eco24295, w_eco24296, w_eco24297, w_eco24298, w_eco24299, w_eco24300, w_eco24301, w_eco24302, w_eco24303, w_eco24304, w_eco24305, w_eco24306, w_eco24307, w_eco24308, w_eco24309, w_eco24310, w_eco24311, w_eco24312, w_eco24313, w_eco24314, w_eco24315, w_eco24316, w_eco24317, w_eco24318, w_eco24319, w_eco24320, w_eco24321, w_eco24322, w_eco24323, w_eco24324, w_eco24325, w_eco24326, w_eco24327, w_eco24328, w_eco24329, w_eco24330, w_eco24331, w_eco24332, w_eco24333, w_eco24334, w_eco24335, w_eco24336, w_eco24337, w_eco24338, w_eco24339, w_eco24340, w_eco24341, w_eco24342, w_eco24343, w_eco24344, w_eco24345, w_eco24346, w_eco24347, w_eco24348, w_eco24349, w_eco24350, w_eco24351, w_eco24352, w_eco24353, w_eco24354, w_eco24355, w_eco24356, w_eco24357, w_eco24358, w_eco24359, w_eco24360, w_eco24361, w_eco24362, w_eco24363, w_eco24364, w_eco24365, w_eco24366, w_eco24367, w_eco24368, w_eco24369, w_eco24370, w_eco24371, w_eco24372, w_eco24373, w_eco24374, w_eco24375, w_eco24376, w_eco24377, w_eco24378, w_eco24379, w_eco24380, w_eco24381, w_eco24382, w_eco24383, w_eco24384, w_eco24385, w_eco24386, w_eco24387, w_eco24388, w_eco24389, w_eco24390, w_eco24391, w_eco24392, w_eco24393, w_eco24394, w_eco24395, w_eco24396, w_eco24397, w_eco24398, w_eco24399, w_eco24400, w_eco24401, w_eco24402, w_eco24403, w_eco24404, w_eco24405, w_eco24406, w_eco24407, w_eco24408, w_eco24409, w_eco24410, w_eco24411, w_eco24412, w_eco24413, w_eco24414, w_eco24415, w_eco24416, w_eco24417, w_eco24418, w_eco24419, w_eco24420, w_eco24421, w_eco24422, w_eco24423, w_eco24424, w_eco24425, w_eco24426, w_eco24427, w_eco24428, w_eco24429, w_eco24430, w_eco24431, w_eco24432, w_eco24433, w_eco24434, w_eco24435, w_eco24436, w_eco24437, w_eco24438, w_eco24439, w_eco24440, w_eco24441, w_eco24442, w_eco24443, w_eco24444, w_eco24445, w_eco24446, w_eco24447, w_eco24448, w_eco24449, w_eco24450, w_eco24451, w_eco24452, w_eco24453, w_eco24454, w_eco24455, w_eco24456, w_eco24457, w_eco24458, w_eco24459, w_eco24460, w_eco24461, w_eco24462, w_eco24463, w_eco24464, w_eco24465, w_eco24466, w_eco24467, w_eco24468, w_eco24469, w_eco24470, w_eco24471, w_eco24472, w_eco24473, w_eco24474, w_eco24475, w_eco24476, w_eco24477, w_eco24478, w_eco24479, w_eco24480, w_eco24481, w_eco24482, w_eco24483, w_eco24484, w_eco24485, w_eco24486, w_eco24487, w_eco24488, w_eco24489, w_eco24490, w_eco24491, w_eco24492, w_eco24493, w_eco24494, w_eco24495, w_eco24496, w_eco24497, w_eco24498, w_eco24499, w_eco24500, w_eco24501, w_eco24502, w_eco24503, w_eco24504, w_eco24505, w_eco24506, w_eco24507, w_eco24508, w_eco24509, w_eco24510, w_eco24511, w_eco24512, w_eco24513, w_eco24514, w_eco24515, w_eco24516, w_eco24517, w_eco24518, w_eco24519, w_eco24520, w_eco24521, w_eco24522, w_eco24523, w_eco24524, w_eco24525, w_eco24526, w_eco24527, w_eco24528, w_eco24529, w_eco24530, w_eco24531, w_eco24532, w_eco24533, w_eco24534, w_eco24535, w_eco24536, w_eco24537, w_eco24538, w_eco24539, w_eco24540, w_eco24541, w_eco24542, w_eco24543, w_eco24544, w_eco24545, w_eco24546, w_eco24547, w_eco24548, w_eco24549, w_eco24550, w_eco24551, w_eco24552, w_eco24553, w_eco24554, w_eco24555, w_eco24556, w_eco24557, w_eco24558, w_eco24559, w_eco24560, w_eco24561, w_eco24562, w_eco24563, w_eco24564, w_eco24565, w_eco24566, w_eco24567, w_eco24568, w_eco24569, w_eco24570, w_eco24571, w_eco24572, w_eco24573, w_eco24574, w_eco24575, w_eco24576, w_eco24577, w_eco24578, w_eco24579, w_eco24580, w_eco24581, w_eco24582, w_eco24583, w_eco24584, w_eco24585, w_eco24586, w_eco24587, w_eco24588, w_eco24589, w_eco24590, w_eco24591, w_eco24592, w_eco24593, w_eco24594, w_eco24595, w_eco24596, w_eco24597, w_eco24598, w_eco24599, w_eco24600, w_eco24601, w_eco24602, w_eco24603, w_eco24604, w_eco24605, w_eco24606, w_eco24607, w_eco24608, w_eco24609, w_eco24610, w_eco24611, w_eco24612, w_eco24613, w_eco24614, w_eco24615, w_eco24616, w_eco24617, w_eco24618, w_eco24619, w_eco24620, w_eco24621, w_eco24622, w_eco24623, w_eco24624, w_eco24625, w_eco24626, w_eco24627, w_eco24628, w_eco24629, w_eco24630, w_eco24631, w_eco24632, w_eco24633, w_eco24634, w_eco24635, w_eco24636, w_eco24637, w_eco24638, w_eco24639, w_eco24640, w_eco24641, w_eco24642, w_eco24643, w_eco24644, w_eco24645, w_eco24646, w_eco24647, w_eco24648, w_eco24649, w_eco24650, w_eco24651, w_eco24652, w_eco24653, w_eco24654, w_eco24655, w_eco24656, w_eco24657, w_eco24658, w_eco24659, w_eco24660, w_eco24661, w_eco24662, w_eco24663, w_eco24664, w_eco24665, w_eco24666, w_eco24667, w_eco24668, w_eco24669, w_eco24670, w_eco24671, w_eco24672, w_eco24673, w_eco24674, w_eco24675, w_eco24676, w_eco24677, w_eco24678, w_eco24679, w_eco24680, w_eco24681, w_eco24682, w_eco24683, w_eco24684, w_eco24685, w_eco24686, w_eco24687, w_eco24688, w_eco24689, w_eco24690, w_eco24691, w_eco24692, w_eco24693, w_eco24694, w_eco24695, w_eco24696, w_eco24697, w_eco24698, w_eco24699, w_eco24700, w_eco24701, w_eco24702, w_eco24703, w_eco24704, w_eco24705, w_eco24706, w_eco24707, w_eco24708, w_eco24709, w_eco24710, w_eco24711, w_eco24712, w_eco24713, w_eco24714, w_eco24715, w_eco24716, w_eco24717, w_eco24718, w_eco24719, w_eco24720, w_eco24721, w_eco24722, w_eco24723, w_eco24724, w_eco24725, w_eco24726, w_eco24727, w_eco24728, w_eco24729, w_eco24730, w_eco24731, w_eco24732, w_eco24733, w_eco24734, w_eco24735, w_eco24736, w_eco24737, w_eco24738, w_eco24739, w_eco24740, w_eco24741, w_eco24742, w_eco24743, w_eco24744, w_eco24745, w_eco24746, w_eco24747, w_eco24748, w_eco24749, w_eco24750, w_eco24751, w_eco24752, w_eco24753, w_eco24754, w_eco24755, w_eco24756, w_eco24757, w_eco24758, w_eco24759, w_eco24760, w_eco24761, w_eco24762, w_eco24763, w_eco24764, w_eco24765, w_eco24766, w_eco24767, w_eco24768, w_eco24769, w_eco24770, w_eco24771, w_eco24772, w_eco24773, w_eco24774, w_eco24775, w_eco24776, w_eco24777, w_eco24778, w_eco24779, w_eco24780, w_eco24781, w_eco24782, w_eco24783, w_eco24784, w_eco24785, w_eco24786, w_eco24787, w_eco24788, w_eco24789, w_eco24790, w_eco24791, w_eco24792, w_eco24793, w_eco24794, w_eco24795, w_eco24796, w_eco24797, w_eco24798, w_eco24799, w_eco24800, w_eco24801, w_eco24802, w_eco24803, w_eco24804, w_eco24805, w_eco24806, w_eco24807, w_eco24808, w_eco24809, w_eco24810, w_eco24811, w_eco24812, w_eco24813, w_eco24814, w_eco24815, w_eco24816, w_eco24817, w_eco24818, w_eco24819, w_eco24820, w_eco24821, w_eco24822, w_eco24823, w_eco24824, w_eco24825, w_eco24826, w_eco24827, w_eco24828, w_eco24829, w_eco24830, w_eco24831, w_eco24832, w_eco24833, w_eco24834, w_eco24835, w_eco24836, w_eco24837, w_eco24838, w_eco24839, w_eco24840, w_eco24841, w_eco24842, w_eco24843, w_eco24844, w_eco24845, w_eco24846, w_eco24847, w_eco24848, w_eco24849, w_eco24850, w_eco24851, w_eco24852, w_eco24853, w_eco24854, w_eco24855, w_eco24856, w_eco24857, w_eco24858, w_eco24859, w_eco24860, w_eco24861, w_eco24862, w_eco24863, w_eco24864, w_eco24865, w_eco24866, w_eco24867, w_eco24868, w_eco24869, w_eco24870, w_eco24871, w_eco24872, w_eco24873, w_eco24874, w_eco24875, w_eco24876, w_eco24877, w_eco24878, w_eco24879, w_eco24880, w_eco24881, w_eco24882, w_eco24883, w_eco24884, w_eco24885, w_eco24886, w_eco24887, w_eco24888, w_eco24889, w_eco24890, w_eco24891, w_eco24892, w_eco24893, w_eco24894, w_eco24895, w_eco24896, w_eco24897, w_eco24898, w_eco24899, w_eco24900, w_eco24901, w_eco24902, w_eco24903, w_eco24904, w_eco24905, w_eco24906, w_eco24907, w_eco24908, w_eco24909, w_eco24910, w_eco24911, w_eco24912, w_eco24913, w_eco24914, w_eco24915, w_eco24916, w_eco24917, w_eco24918, w_eco24919, w_eco24920, w_eco24921, w_eco24922, w_eco24923, w_eco24924, w_eco24925, w_eco24926, w_eco24927, w_eco24928, w_eco24929, w_eco24930, w_eco24931, w_eco24932, w_eco24933, w_eco24934, w_eco24935, w_eco24936, w_eco24937, w_eco24938, w_eco24939, w_eco24940, w_eco24941, w_eco24942, w_eco24943, w_eco24944, w_eco24945, w_eco24946, w_eco24947, w_eco24948, w_eco24949, w_eco24950, w_eco24951, w_eco24952, w_eco24953, w_eco24954, w_eco24955, w_eco24956, w_eco24957, w_eco24958, w_eco24959, w_eco24960, w_eco24961, w_eco24962, w_eco24963, w_eco24964, w_eco24965, w_eco24966, w_eco24967, w_eco24968, w_eco24969, w_eco24970, w_eco24971, w_eco24972, w_eco24973, w_eco24974, w_eco24975, w_eco24976, w_eco24977, w_eco24978, w_eco24979, w_eco24980, w_eco24981, w_eco24982, w_eco24983, w_eco24984, w_eco24985, w_eco24986, w_eco24987, w_eco24988, w_eco24989, w_eco24990, w_eco24991, w_eco24992, w_eco24993, w_eco24994, w_eco24995, w_eco24996, w_eco24997, w_eco24998, w_eco24999, w_eco25000, w_eco25001, w_eco25002, w_eco25003, w_eco25004, w_eco25005, w_eco25006, w_eco25007, w_eco25008, w_eco25009, w_eco25010, w_eco25011, w_eco25012, w_eco25013, w_eco25014, w_eco25015, w_eco25016, w_eco25017, w_eco25018, w_eco25019, w_eco25020, w_eco25021, w_eco25022, w_eco25023, w_eco25024, w_eco25025, w_eco25026, w_eco25027, w_eco25028, w_eco25029, w_eco25030, w_eco25031, w_eco25032, w_eco25033, w_eco25034, w_eco25035, w_eco25036, w_eco25037, w_eco25038, w_eco25039, w_eco25040, w_eco25041, w_eco25042, w_eco25043, w_eco25044, w_eco25045, w_eco25046, w_eco25047, w_eco25048, w_eco25049, w_eco25050, w_eco25051, w_eco25052, w_eco25053, w_eco25054, w_eco25055, w_eco25056, w_eco25057, w_eco25058, w_eco25059, w_eco25060, w_eco25061, w_eco25062, w_eco25063, w_eco25064, w_eco25065, w_eco25066, w_eco25067, w_eco25068, w_eco25069, w_eco25070, w_eco25071, w_eco25072, w_eco25073, w_eco25074, w_eco25075, w_eco25076, w_eco25077, w_eco25078, w_eco25079, w_eco25080, w_eco25081, w_eco25082, w_eco25083, w_eco25084, w_eco25085, w_eco25086, w_eco25087, w_eco25088, w_eco25089, w_eco25090, w_eco25091, w_eco25092, w_eco25093, w_eco25094, w_eco25095, w_eco25096, w_eco25097, w_eco25098, w_eco25099, w_eco25100, w_eco25101, w_eco25102, w_eco25103, w_eco25104, w_eco25105, w_eco25106, w_eco25107, w_eco25108, w_eco25109, w_eco25110, w_eco25111, w_eco25112, w_eco25113, w_eco25114, w_eco25115, w_eco25116, w_eco25117, w_eco25118, w_eco25119, w_eco25120, w_eco25121, w_eco25122, w_eco25123, w_eco25124, w_eco25125, w_eco25126, w_eco25127, w_eco25128, w_eco25129, w_eco25130, w_eco25131, w_eco25132, w_eco25133, w_eco25134, w_eco25135, w_eco25136, w_eco25137, w_eco25138, w_eco25139, w_eco25140, w_eco25141, w_eco25142, w_eco25143, w_eco25144, w_eco25145, w_eco25146, w_eco25147, w_eco25148, w_eco25149, w_eco25150, w_eco25151, w_eco25152, w_eco25153, w_eco25154, w_eco25155, w_eco25156, w_eco25157, w_eco25158, w_eco25159, w_eco25160, w_eco25161, w_eco25162, w_eco25163, w_eco25164, w_eco25165, w_eco25166, w_eco25167, w_eco25168, w_eco25169, w_eco25170, w_eco25171, w_eco25172, w_eco25173, w_eco25174, w_eco25175, w_eco25176, w_eco25177, w_eco25178, w_eco25179, w_eco25180, w_eco25181, w_eco25182, w_eco25183, w_eco25184, w_eco25185, w_eco25186, w_eco25187, w_eco25188, w_eco25189, w_eco25190, w_eco25191, w_eco25192, w_eco25193, w_eco25194, w_eco25195, w_eco25196, w_eco25197, w_eco25198, w_eco25199, w_eco25200, w_eco25201, w_eco25202, w_eco25203, w_eco25204, w_eco25205, w_eco25206, w_eco25207, w_eco25208, w_eco25209, w_eco25210, w_eco25211, w_eco25212, w_eco25213, w_eco25214, w_eco25215, w_eco25216, w_eco25217, w_eco25218, w_eco25219, w_eco25220, w_eco25221, w_eco25222, w_eco25223, w_eco25224, w_eco25225, w_eco25226, w_eco25227, w_eco25228, w_eco25229, w_eco25230, w_eco25231, w_eco25232, w_eco25233, w_eco25234, w_eco25235, w_eco25236, w_eco25237, w_eco25238, w_eco25239, w_eco25240, w_eco25241, w_eco25242, w_eco25243, w_eco25244, w_eco25245, w_eco25246, w_eco25247, w_eco25248, w_eco25249, w_eco25250, w_eco25251, w_eco25252, w_eco25253, w_eco25254, w_eco25255, w_eco25256, w_eco25257, w_eco25258, w_eco25259, w_eco25260, w_eco25261, w_eco25262, w_eco25263, w_eco25264, w_eco25265, w_eco25266, w_eco25267, w_eco25268, w_eco25269, w_eco25270, w_eco25271, w_eco25272, w_eco25273, w_eco25274, w_eco25275, w_eco25276, w_eco25277, w_eco25278, w_eco25279, w_eco25280, w_eco25281, w_eco25282, w_eco25283, w_eco25284, w_eco25285, w_eco25286, w_eco25287, w_eco25288, w_eco25289, w_eco25290, w_eco25291, w_eco25292, w_eco25293, w_eco25294, w_eco25295, w_eco25296, w_eco25297, w_eco25298, w_eco25299, w_eco25300, w_eco25301, w_eco25302, w_eco25303, w_eco25304, w_eco25305, w_eco25306, w_eco25307, w_eco25308, w_eco25309, w_eco25310, w_eco25311, w_eco25312, w_eco25313, w_eco25314, w_eco25315, w_eco25316, w_eco25317, w_eco25318, w_eco25319, w_eco25320, w_eco25321, w_eco25322, w_eco25323, w_eco25324, w_eco25325, w_eco25326, w_eco25327, w_eco25328, w_eco25329, w_eco25330, w_eco25331, w_eco25332, w_eco25333, w_eco25334, w_eco25335, w_eco25336, w_eco25337, w_eco25338, w_eco25339, w_eco25340, w_eco25341, w_eco25342, w_eco25343, w_eco25344, w_eco25345, w_eco25346, w_eco25347, w_eco25348, w_eco25349, w_eco25350, w_eco25351, w_eco25352, w_eco25353, w_eco25354, w_eco25355, w_eco25356, w_eco25357, w_eco25358, w_eco25359, w_eco25360, w_eco25361, w_eco25362, w_eco25363, w_eco25364, w_eco25365, w_eco25366, w_eco25367, w_eco25368, w_eco25369, w_eco25370, w_eco25371, w_eco25372, w_eco25373, w_eco25374, w_eco25375, w_eco25376, w_eco25377, w_eco25378, w_eco25379, w_eco25380, w_eco25381, w_eco25382, w_eco25383, w_eco25384, w_eco25385, w_eco25386, w_eco25387, w_eco25388, w_eco25389, w_eco25390, w_eco25391, w_eco25392, w_eco25393, w_eco25394, w_eco25395, w_eco25396, w_eco25397, w_eco25398, w_eco25399, w_eco25400, w_eco25401, w_eco25402, w_eco25403, w_eco25404, w_eco25405, w_eco25406, w_eco25407, w_eco25408, w_eco25409, w_eco25410, w_eco25411, w_eco25412, w_eco25413, w_eco25414, w_eco25415, w_eco25416, w_eco25417, w_eco25418, w_eco25419, w_eco25420, w_eco25421, w_eco25422, w_eco25423, w_eco25424, w_eco25425, w_eco25426, w_eco25427, w_eco25428, w_eco25429, w_eco25430, w_eco25431, w_eco25432, w_eco25433, w_eco25434, w_eco25435, w_eco25436, w_eco25437, w_eco25438, w_eco25439, w_eco25440, w_eco25441, w_eco25442, w_eco25443, w_eco25444, w_eco25445, w_eco25446, w_eco25447, w_eco25448, w_eco25449, w_eco25450, w_eco25451, w_eco25452, w_eco25453, w_eco25454, w_eco25455, w_eco25456, w_eco25457, w_eco25458, w_eco25459, w_eco25460, w_eco25461, w_eco25462, w_eco25463, w_eco25464, w_eco25465, w_eco25466, w_eco25467, w_eco25468, w_eco25469, w_eco25470, w_eco25471, w_eco25472, w_eco25473, w_eco25474, w_eco25475, w_eco25476, w_eco25477, w_eco25478, w_eco25479, w_eco25480, w_eco25481, w_eco25482, w_eco25483, w_eco25484, w_eco25485, w_eco25486, w_eco25487, w_eco25488, w_eco25489, w_eco25490, w_eco25491, w_eco25492, w_eco25493, w_eco25494, w_eco25495, w_eco25496, w_eco25497, w_eco25498, w_eco25499, w_eco25500, w_eco25501, w_eco25502, w_eco25503, w_eco25504, w_eco25505, w_eco25506, w_eco25507, w_eco25508, w_eco25509, w_eco25510, w_eco25511, w_eco25512, w_eco25513, w_eco25514, w_eco25515, w_eco25516, w_eco25517, w_eco25518, w_eco25519, w_eco25520, w_eco25521, w_eco25522, w_eco25523, w_eco25524, w_eco25525, w_eco25526, w_eco25527, w_eco25528, w_eco25529, w_eco25530, w_eco25531, w_eco25532, w_eco25533, w_eco25534, w_eco25535, w_eco25536, w_eco25537, w_eco25538, w_eco25539, w_eco25540, w_eco25541, w_eco25542, w_eco25543, w_eco25544, w_eco25545, w_eco25546, w_eco25547, w_eco25548, w_eco25549, w_eco25550, w_eco25551, w_eco25552, w_eco25553, w_eco25554, w_eco25555, w_eco25556, w_eco25557, w_eco25558, w_eco25559, w_eco25560, w_eco25561, w_eco25562, w_eco25563, w_eco25564, w_eco25565, w_eco25566, w_eco25567, w_eco25568, w_eco25569, w_eco25570, w_eco25571, w_eco25572, w_eco25573, w_eco25574, w_eco25575, w_eco25576, w_eco25577, w_eco25578, w_eco25579, w_eco25580, w_eco25581, w_eco25582, w_eco25583, w_eco25584, w_eco25585, w_eco25586, w_eco25587, w_eco25588, w_eco25589, w_eco25590, w_eco25591, w_eco25592, w_eco25593, w_eco25594, w_eco25595, w_eco25596, w_eco25597, w_eco25598, w_eco25599, w_eco25600, w_eco25601, w_eco25602, w_eco25603, w_eco25604, w_eco25605, w_eco25606, w_eco25607, w_eco25608, w_eco25609, w_eco25610, w_eco25611, w_eco25612, w_eco25613, w_eco25614, w_eco25615, w_eco25616, w_eco25617, w_eco25618, w_eco25619, w_eco25620, w_eco25621, w_eco25622, w_eco25623, w_eco25624, w_eco25625, w_eco25626, w_eco25627, w_eco25628, w_eco25629, w_eco25630, w_eco25631, w_eco25632, w_eco25633, w_eco25634, w_eco25635, w_eco25636, w_eco25637, w_eco25638, w_eco25639, w_eco25640, w_eco25641, w_eco25642, w_eco25643, w_eco25644, w_eco25645, w_eco25646, w_eco25647, w_eco25648, w_eco25649, w_eco25650, w_eco25651, w_eco25652, w_eco25653, w_eco25654, w_eco25655, w_eco25656, w_eco25657, w_eco25658, w_eco25659, w_eco25660, w_eco25661, w_eco25662, w_eco25663, w_eco25664, w_eco25665, w_eco25666, w_eco25667, w_eco25668, w_eco25669, w_eco25670, w_eco25671, w_eco25672, w_eco25673, w_eco25674, w_eco25675, w_eco25676, w_eco25677, w_eco25678, w_eco25679, w_eco25680, w_eco25681, w_eco25682, w_eco25683, w_eco25684, w_eco25685, w_eco25686, w_eco25687, w_eco25688, w_eco25689, w_eco25690, w_eco25691, w_eco25692, w_eco25693, w_eco25694, w_eco25695, w_eco25696, w_eco25697, w_eco25698, w_eco25699, w_eco25700, w_eco25701, w_eco25702, w_eco25703, w_eco25704, w_eco25705, w_eco25706, w_eco25707, w_eco25708, w_eco25709, w_eco25710, w_eco25711, w_eco25712, w_eco25713, w_eco25714, w_eco25715, w_eco25716, w_eco25717, w_eco25718, w_eco25719, w_eco25720, w_eco25721, w_eco25722, w_eco25723, w_eco25724, w_eco25725, w_eco25726, w_eco25727, w_eco25728, w_eco25729, w_eco25730, w_eco25731, w_eco25732, w_eco25733, w_eco25734, w_eco25735, w_eco25736, w_eco25737, w_eco25738, w_eco25739, w_eco25740, w_eco25741, w_eco25742, w_eco25743, w_eco25744, w_eco25745, w_eco25746, w_eco25747, w_eco25748, w_eco25749, w_eco25750, w_eco25751, w_eco25752, w_eco25753, w_eco25754, w_eco25755, w_eco25756, w_eco25757, w_eco25758, w_eco25759, w_eco25760, w_eco25761, w_eco25762, w_eco25763, w_eco25764, w_eco25765, w_eco25766, w_eco25767, w_eco25768, w_eco25769, w_eco25770, w_eco25771, w_eco25772, w_eco25773, w_eco25774, w_eco25775, w_eco25776, w_eco25777, w_eco25778, w_eco25779, w_eco25780, w_eco25781, w_eco25782, w_eco25783, w_eco25784, w_eco25785, w_eco25786, w_eco25787, w_eco25788, w_eco25789, w_eco25790, w_eco25791, w_eco25792, w_eco25793, w_eco25794, w_eco25795, w_eco25796, w_eco25797, w_eco25798, w_eco25799, w_eco25800, w_eco25801, w_eco25802, w_eco25803, w_eco25804, w_eco25805, w_eco25806, w_eco25807, w_eco25808, w_eco25809, w_eco25810, w_eco25811, w_eco25812, w_eco25813, w_eco25814, w_eco25815, w_eco25816, w_eco25817, w_eco25818, w_eco25819, w_eco25820, w_eco25821, w_eco25822, w_eco25823, w_eco25824, w_eco25825, w_eco25826, w_eco25827, w_eco25828, w_eco25829, w_eco25830, w_eco25831, w_eco25832, w_eco25833, w_eco25834, w_eco25835, w_eco25836, w_eco25837, w_eco25838, w_eco25839, w_eco25840, w_eco25841, w_eco25842, w_eco25843, w_eco25844, w_eco25845, w_eco25846, w_eco25847, w_eco25848, w_eco25849, w_eco25850, w_eco25851, w_eco25852, w_eco25853, w_eco25854, w_eco25855, w_eco25856, w_eco25857, w_eco25858, w_eco25859, w_eco25860, w_eco25861, w_eco25862, w_eco25863, w_eco25864, w_eco25865, w_eco25866, w_eco25867, w_eco25868, w_eco25869, w_eco25870, w_eco25871, w_eco25872, w_eco25873, w_eco25874, w_eco25875, w_eco25876, w_eco25877, w_eco25878, w_eco25879, w_eco25880, w_eco25881, w_eco25882, w_eco25883, w_eco25884, w_eco25885, w_eco25886, w_eco25887, w_eco25888, w_eco25889, w_eco25890, w_eco25891, w_eco25892, w_eco25893, w_eco25894, w_eco25895, w_eco25896, w_eco25897, w_eco25898, w_eco25899, w_eco25900, w_eco25901, w_eco25902, w_eco25903, w_eco25904, w_eco25905, w_eco25906, w_eco25907, w_eco25908, w_eco25909, w_eco25910, w_eco25911, w_eco25912, w_eco25913, w_eco25914, w_eco25915, w_eco25916, w_eco25917, w_eco25918, w_eco25919, w_eco25920, w_eco25921, w_eco25922, w_eco25923, w_eco25924, w_eco25925, w_eco25926, w_eco25927, w_eco25928, w_eco25929, w_eco25930, w_eco25931, w_eco25932, w_eco25933, w_eco25934, w_eco25935, w_eco25936, w_eco25937, w_eco25938, w_eco25939, w_eco25940, w_eco25941, w_eco25942, w_eco25943, w_eco25944, w_eco25945, w_eco25946, w_eco25947, w_eco25948, w_eco25949, w_eco25950, w_eco25951, w_eco25952, w_eco25953, w_eco25954, w_eco25955, w_eco25956, w_eco25957, w_eco25958, w_eco25959, w_eco25960, w_eco25961, w_eco25962, w_eco25963, w_eco25964, w_eco25965, w_eco25966, w_eco25967, w_eco25968, w_eco25969, w_eco25970, w_eco25971, w_eco25972, w_eco25973, w_eco25974, w_eco25975, w_eco25976, w_eco25977, w_eco25978, w_eco25979, w_eco25980, w_eco25981, w_eco25982, w_eco25983, w_eco25984, w_eco25985, w_eco25986, w_eco25987, w_eco25988, w_eco25989, w_eco25990, w_eco25991, w_eco25992, w_eco25993, w_eco25994, w_eco25995, w_eco25996, w_eco25997, w_eco25998, w_eco25999, w_eco26000, w_eco26001, w_eco26002, w_eco26003, w_eco26004, w_eco26005, w_eco26006, w_eco26007, w_eco26008, w_eco26009, w_eco26010, w_eco26011, w_eco26012, w_eco26013, w_eco26014, w_eco26015, w_eco26016, w_eco26017, w_eco26018, w_eco26019, w_eco26020, w_eco26021, w_eco26022, w_eco26023, w_eco26024, w_eco26025, w_eco26026, w_eco26027, w_eco26028, w_eco26029, w_eco26030, w_eco26031, w_eco26032, w_eco26033, w_eco26034, w_eco26035, w_eco26036, w_eco26037, w_eco26038, w_eco26039, w_eco26040, w_eco26041, w_eco26042, w_eco26043, w_eco26044, w_eco26045, w_eco26046, w_eco26047, w_eco26048, w_eco26049, w_eco26050, w_eco26051, w_eco26052, w_eco26053, w_eco26054, w_eco26055, w_eco26056, w_eco26057, w_eco26058, w_eco26059, w_eco26060, w_eco26061, w_eco26062, w_eco26063, w_eco26064, w_eco26065, w_eco26066, w_eco26067, w_eco26068, w_eco26069, w_eco26070, w_eco26071, w_eco26072, w_eco26073, w_eco26074, w_eco26075, w_eco26076, w_eco26077, w_eco26078, w_eco26079, w_eco26080, w_eco26081, w_eco26082, w_eco26083, w_eco26084, w_eco26085, w_eco26086, w_eco26087, w_eco26088, w_eco26089, w_eco26090, w_eco26091, w_eco26092, w_eco26093, w_eco26094, w_eco26095, w_eco26096, w_eco26097, w_eco26098, w_eco26099, w_eco26100, w_eco26101, w_eco26102, w_eco26103, w_eco26104, w_eco26105, w_eco26106, w_eco26107, w_eco26108, w_eco26109, w_eco26110, w_eco26111, w_eco26112, w_eco26113, w_eco26114, w_eco26115, w_eco26116, w_eco26117, w_eco26118, w_eco26119, w_eco26120, w_eco26121, w_eco26122, w_eco26123, w_eco26124, w_eco26125, w_eco26126, w_eco26127, w_eco26128, w_eco26129, w_eco26130, w_eco26131, w_eco26132, w_eco26133, w_eco26134, w_eco26135, w_eco26136, w_eco26137, w_eco26138, w_eco26139, w_eco26140, w_eco26141, w_eco26142, w_eco26143, w_eco26144, w_eco26145, w_eco26146, w_eco26147, w_eco26148, w_eco26149, w_eco26150, w_eco26151, w_eco26152, w_eco26153, w_eco26154, w_eco26155, w_eco26156, w_eco26157, w_eco26158, w_eco26159, w_eco26160, w_eco26161, w_eco26162, w_eco26163, w_eco26164, w_eco26165, w_eco26166, w_eco26167, w_eco26168, w_eco26169, w_eco26170, w_eco26171, w_eco26172, w_eco26173, w_eco26174, w_eco26175, w_eco26176, w_eco26177, w_eco26178, w_eco26179, w_eco26180, w_eco26181, w_eco26182, w_eco26183, w_eco26184, w_eco26185, w_eco26186, w_eco26187, w_eco26188, w_eco26189, w_eco26190, w_eco26191, w_eco26192, w_eco26193, w_eco26194, w_eco26195, w_eco26196, w_eco26197, w_eco26198, w_eco26199, w_eco26200, w_eco26201, w_eco26202, w_eco26203, w_eco26204, w_eco26205, w_eco26206, w_eco26207, w_eco26208, w_eco26209, w_eco26210, w_eco26211, w_eco26212, w_eco26213, w_eco26214, w_eco26215, w_eco26216, w_eco26217, w_eco26218, w_eco26219, w_eco26220, w_eco26221, w_eco26222, w_eco26223, w_eco26224, w_eco26225, w_eco26226, w_eco26227, w_eco26228, w_eco26229, w_eco26230, w_eco26231, w_eco26232, w_eco26233, w_eco26234, w_eco26235, w_eco26236, w_eco26237, w_eco26238, w_eco26239, w_eco26240, w_eco26241, w_eco26242, w_eco26243, w_eco26244, w_eco26245, w_eco26246, w_eco26247, w_eco26248, w_eco26249, w_eco26250, w_eco26251, w_eco26252, w_eco26253, w_eco26254, w_eco26255, w_eco26256, w_eco26257, w_eco26258, w_eco26259, w_eco26260, w_eco26261, w_eco26262, w_eco26263, w_eco26264, w_eco26265, w_eco26266, w_eco26267, w_eco26268, w_eco26269, w_eco26270, w_eco26271, w_eco26272, w_eco26273, w_eco26274, w_eco26275, w_eco26276, w_eco26277, w_eco26278, w_eco26279, w_eco26280, w_eco26281, w_eco26282, w_eco26283, w_eco26284, w_eco26285, w_eco26286, w_eco26287, w_eco26288, w_eco26289, w_eco26290, w_eco26291, w_eco26292, w_eco26293, w_eco26294, w_eco26295, w_eco26296, w_eco26297, w_eco26298, w_eco26299, w_eco26300, w_eco26301, w_eco26302, w_eco26303, w_eco26304, w_eco26305, w_eco26306, w_eco26307, w_eco26308, w_eco26309, w_eco26310, w_eco26311, w_eco26312, w_eco26313, w_eco26314, w_eco26315, w_eco26316, w_eco26317, w_eco26318, w_eco26319, w_eco26320, w_eco26321, w_eco26322, w_eco26323, w_eco26324, w_eco26325, w_eco26326, w_eco26327, w_eco26328, w_eco26329, w_eco26330, w_eco26331, w_eco26332, w_eco26333, w_eco26334, w_eco26335, w_eco26336, w_eco26337, w_eco26338, w_eco26339, w_eco26340, w_eco26341, w_eco26342, w_eco26343, w_eco26344, w_eco26345, w_eco26346, w_eco26347, w_eco26348, w_eco26349, w_eco26350, w_eco26351, w_eco26352, w_eco26353, w_eco26354, w_eco26355, w_eco26356, w_eco26357, w_eco26358, w_eco26359, w_eco26360, w_eco26361, w_eco26362, w_eco26363, w_eco26364, w_eco26365, w_eco26366, w_eco26367, w_eco26368, w_eco26369, w_eco26370, w_eco26371, w_eco26372, w_eco26373, w_eco26374, w_eco26375, w_eco26376, w_eco26377, w_eco26378, w_eco26379, w_eco26380, w_eco26381, w_eco26382, w_eco26383, w_eco26384, w_eco26385, w_eco26386, w_eco26387, w_eco26388, w_eco26389, w_eco26390, w_eco26391, w_eco26392, w_eco26393, w_eco26394, w_eco26395, w_eco26396, w_eco26397, w_eco26398, w_eco26399, w_eco26400, w_eco26401, w_eco26402, w_eco26403, w_eco26404, w_eco26405, w_eco26406, w_eco26407, w_eco26408, w_eco26409, w_eco26410, w_eco26411, w_eco26412, w_eco26413, w_eco26414, w_eco26415, w_eco26416, w_eco26417, w_eco26418, w_eco26419, w_eco26420, w_eco26421, w_eco26422, w_eco26423, w_eco26424, w_eco26425, w_eco26426, w_eco26427, w_eco26428, w_eco26429, w_eco26430, w_eco26431, w_eco26432, w_eco26433, w_eco26434, w_eco26435, w_eco26436, w_eco26437, w_eco26438, w_eco26439, w_eco26440, w_eco26441, w_eco26442, w_eco26443, w_eco26444, w_eco26445, w_eco26446, w_eco26447, w_eco26448, w_eco26449, w_eco26450, w_eco26451, w_eco26452, w_eco26453, w_eco26454, w_eco26455, w_eco26456, w_eco26457, w_eco26458, w_eco26459, w_eco26460, w_eco26461, w_eco26462, w_eco26463, w_eco26464, w_eco26465, w_eco26466, w_eco26467, w_eco26468, w_eco26469, w_eco26470, w_eco26471, w_eco26472, w_eco26473, w_eco26474, w_eco26475, w_eco26476, w_eco26477, w_eco26478, w_eco26479, w_eco26480, w_eco26481, w_eco26482, w_eco26483, w_eco26484, w_eco26485, w_eco26486, w_eco26487, w_eco26488, w_eco26489, w_eco26490, w_eco26491, w_eco26492, w_eco26493, w_eco26494, w_eco26495, w_eco26496, w_eco26497, w_eco26498, w_eco26499, w_eco26500, w_eco26501, w_eco26502, w_eco26503, w_eco26504, w_eco26505, w_eco26506, w_eco26507, w_eco26508, w_eco26509, w_eco26510, w_eco26511, w_eco26512, w_eco26513, w_eco26514, w_eco26515, w_eco26516, w_eco26517, w_eco26518, w_eco26519, w_eco26520, w_eco26521, w_eco26522, w_eco26523, w_eco26524, w_eco26525, w_eco26526, w_eco26527, w_eco26528, w_eco26529, w_eco26530, w_eco26531, w_eco26532, w_eco26533, w_eco26534, w_eco26535, w_eco26536, w_eco26537, w_eco26538, w_eco26539, w_eco26540, w_eco26541, w_eco26542, w_eco26543, w_eco26544, w_eco26545, w_eco26546, w_eco26547, w_eco26548, w_eco26549, w_eco26550, w_eco26551, w_eco26552, w_eco26553, w_eco26554, w_eco26555, w_eco26556, w_eco26557, w_eco26558, w_eco26559, w_eco26560, w_eco26561, w_eco26562, w_eco26563, w_eco26564, w_eco26565, w_eco26566, w_eco26567, w_eco26568, w_eco26569, w_eco26570, w_eco26571, w_eco26572, w_eco26573, w_eco26574, w_eco26575, w_eco26576, w_eco26577, w_eco26578, w_eco26579, w_eco26580, w_eco26581, w_eco26582, w_eco26583, w_eco26584, w_eco26585, w_eco26586, w_eco26587, w_eco26588, w_eco26589, w_eco26590, w_eco26591, w_eco26592, w_eco26593, w_eco26594, w_eco26595, w_eco26596, w_eco26597, w_eco26598, w_eco26599, w_eco26600, w_eco26601, w_eco26602, w_eco26603, w_eco26604, w_eco26605, w_eco26606, w_eco26607, w_eco26608, w_eco26609, w_eco26610, w_eco26611, w_eco26612, w_eco26613, w_eco26614, w_eco26615, w_eco26616, w_eco26617, w_eco26618, w_eco26619, w_eco26620, w_eco26621, w_eco26622, w_eco26623, w_eco26624, w_eco26625, w_eco26626, w_eco26627, w_eco26628, w_eco26629, w_eco26630, w_eco26631, w_eco26632, w_eco26633, w_eco26634, w_eco26635, w_eco26636, w_eco26637, w_eco26638, w_eco26639, w_eco26640, w_eco26641, w_eco26642, w_eco26643, w_eco26644, w_eco26645, w_eco26646, w_eco26647, w_eco26648, w_eco26649, w_eco26650, w_eco26651, w_eco26652, w_eco26653, w_eco26654, w_eco26655, w_eco26656, w_eco26657, w_eco26658, w_eco26659, w_eco26660, w_eco26661, w_eco26662, w_eco26663, w_eco26664, w_eco26665, w_eco26666, w_eco26667, w_eco26668, w_eco26669, w_eco26670, w_eco26671, w_eco26672, w_eco26673, w_eco26674, w_eco26675, w_eco26676, w_eco26677, w_eco26678, w_eco26679, w_eco26680, w_eco26681, w_eco26682, w_eco26683, w_eco26684, w_eco26685, w_eco26686, w_eco26687, w_eco26688, w_eco26689, w_eco26690, w_eco26691, w_eco26692, w_eco26693, w_eco26694, w_eco26695, w_eco26696, w_eco26697, w_eco26698, w_eco26699, w_eco26700, w_eco26701, w_eco26702, w_eco26703, w_eco26704, w_eco26705, w_eco26706, w_eco26707, w_eco26708, w_eco26709, w_eco26710, w_eco26711, w_eco26712, w_eco26713, w_eco26714, w_eco26715, w_eco26716, w_eco26717, w_eco26718, w_eco26719, w_eco26720, w_eco26721, w_eco26722, w_eco26723, w_eco26724, w_eco26725, w_eco26726, w_eco26727, w_eco26728, w_eco26729, w_eco26730, w_eco26731, w_eco26732, w_eco26733, w_eco26734, w_eco26735, w_eco26736, w_eco26737, w_eco26738, w_eco26739, w_eco26740, w_eco26741, w_eco26742, w_eco26743, w_eco26744, w_eco26745, w_eco26746, w_eco26747, w_eco26748, w_eco26749, w_eco26750, w_eco26751, w_eco26752, w_eco26753, w_eco26754, w_eco26755, w_eco26756, w_eco26757, w_eco26758, w_eco26759, w_eco26760, w_eco26761, w_eco26762, w_eco26763, w_eco26764, w_eco26765, w_eco26766, w_eco26767, w_eco26768, w_eco26769, w_eco26770, w_eco26771, w_eco26772, w_eco26773, w_eco26774, w_eco26775, w_eco26776, w_eco26777, w_eco26778, w_eco26779, w_eco26780, w_eco26781, w_eco26782, w_eco26783, w_eco26784, w_eco26785, w_eco26786, w_eco26787, w_eco26788, w_eco26789, w_eco26790, w_eco26791, w_eco26792, w_eco26793, w_eco26794, w_eco26795, w_eco26796, w_eco26797, w_eco26798, w_eco26799, w_eco26800, w_eco26801, w_eco26802, w_eco26803, w_eco26804, w_eco26805, w_eco26806, w_eco26807, w_eco26808, w_eco26809, w_eco26810, w_eco26811, w_eco26812, w_eco26813, w_eco26814, w_eco26815, w_eco26816, w_eco26817, w_eco26818, w_eco26819, w_eco26820, w_eco26821, w_eco26822, w_eco26823, w_eco26824, w_eco26825, w_eco26826, w_eco26827, w_eco26828, w_eco26829, w_eco26830, w_eco26831, w_eco26832, w_eco26833, w_eco26834, w_eco26835, w_eco26836, w_eco26837, w_eco26838, w_eco26839, w_eco26840, w_eco26841, w_eco26842, w_eco26843, w_eco26844, w_eco26845, w_eco26846, w_eco26847, w_eco26848, w_eco26849, w_eco26850, w_eco26851, w_eco26852, w_eco26853, w_eco26854, w_eco26855, w_eco26856, w_eco26857, w_eco26858, w_eco26859, w_eco26860, w_eco26861, w_eco26862, w_eco26863, w_eco26864, w_eco26865, w_eco26866, w_eco26867, w_eco26868, w_eco26869, w_eco26870, w_eco26871, w_eco26872, w_eco26873, w_eco26874, w_eco26875, w_eco26876, w_eco26877, w_eco26878, w_eco26879, w_eco26880, w_eco26881, w_eco26882, w_eco26883, w_eco26884, w_eco26885, w_eco26886, w_eco26887, w_eco26888, w_eco26889, w_eco26890, w_eco26891, w_eco26892, w_eco26893, w_eco26894, w_eco26895, w_eco26896, w_eco26897, w_eco26898, w_eco26899, w_eco26900, w_eco26901, w_eco26902, w_eco26903, w_eco26904, w_eco26905, w_eco26906, w_eco26907, w_eco26908, w_eco26909, w_eco26910, w_eco26911, w_eco26912, w_eco26913, w_eco26914, w_eco26915, w_eco26916, w_eco26917, w_eco26918, w_eco26919, w_eco26920, w_eco26921, w_eco26922, w_eco26923, w_eco26924, w_eco26925, w_eco26926, w_eco26927, w_eco26928, w_eco26929, w_eco26930, w_eco26931, w_eco26932, w_eco26933, w_eco26934, w_eco26935, w_eco26936, w_eco26937, w_eco26938, w_eco26939, w_eco26940, w_eco26941, w_eco26942, w_eco26943, w_eco26944, w_eco26945, w_eco26946, w_eco26947, w_eco26948, w_eco26949, w_eco26950, w_eco26951, w_eco26952, w_eco26953, w_eco26954, w_eco26955, w_eco26956, w_eco26957, w_eco26958, w_eco26959, w_eco26960, w_eco26961, w_eco26962, w_eco26963, w_eco26964, w_eco26965, w_eco26966, w_eco26967, w_eco26968, w_eco26969, w_eco26970, w_eco26971, w_eco26972, w_eco26973, w_eco26974, w_eco26975, w_eco26976, w_eco26977, w_eco26978, w_eco26979, w_eco26980, w_eco26981, w_eco26982, w_eco26983, w_eco26984, w_eco26985, w_eco26986, w_eco26987, w_eco26988, w_eco26989, w_eco26990, w_eco26991, w_eco26992, w_eco26993, w_eco26994, w_eco26995, w_eco26996, w_eco26997, w_eco26998, w_eco26999, w_eco27000, w_eco27001, w_eco27002, w_eco27003, w_eco27004, w_eco27005, w_eco27006, w_eco27007, w_eco27008, w_eco27009, w_eco27010, w_eco27011, w_eco27012, w_eco27013, w_eco27014, w_eco27015, w_eco27016, w_eco27017, w_eco27018, w_eco27019, w_eco27020, w_eco27021, w_eco27022, w_eco27023, w_eco27024, w_eco27025, w_eco27026, w_eco27027, w_eco27028, w_eco27029, w_eco27030, w_eco27031, w_eco27032, w_eco27033, w_eco27034, w_eco27035, w_eco27036, w_eco27037, w_eco27038, w_eco27039, w_eco27040, w_eco27041, w_eco27042, w_eco27043, w_eco27044, w_eco27045, w_eco27046, w_eco27047, w_eco27048, w_eco27049, w_eco27050, w_eco27051, w_eco27052, w_eco27053, w_eco27054, w_eco27055, w_eco27056, w_eco27057, w_eco27058, w_eco27059, w_eco27060, w_eco27061, w_eco27062, w_eco27063, w_eco27064, w_eco27065, w_eco27066, w_eco27067, w_eco27068, w_eco27069, w_eco27070, w_eco27071, w_eco27072, w_eco27073, w_eco27074, w_eco27075, w_eco27076, w_eco27077, w_eco27078, w_eco27079, w_eco27080, w_eco27081, w_eco27082, w_eco27083, w_eco27084, w_eco27085, w_eco27086, w_eco27087, w_eco27088, w_eco27089, w_eco27090, w_eco27091, w_eco27092, w_eco27093, w_eco27094, w_eco27095, w_eco27096, w_eco27097, w_eco27098, w_eco27099, w_eco27100, w_eco27101, w_eco27102, w_eco27103, w_eco27104, w_eco27105, w_eco27106, w_eco27107, w_eco27108, w_eco27109, w_eco27110, w_eco27111, w_eco27112, w_eco27113, w_eco27114, w_eco27115, w_eco27116, w_eco27117, w_eco27118, w_eco27119, w_eco27120, w_eco27121, w_eco27122, w_eco27123, w_eco27124, w_eco27125, w_eco27126, w_eco27127, w_eco27128, w_eco27129, w_eco27130, w_eco27131, w_eco27132, w_eco27133, w_eco27134, w_eco27135, w_eco27136, w_eco27137, w_eco27138, w_eco27139, w_eco27140, w_eco27141, w_eco27142, w_eco27143, w_eco27144, w_eco27145, w_eco27146, w_eco27147, w_eco27148, w_eco27149, w_eco27150, w_eco27151, w_eco27152, w_eco27153, w_eco27154, w_eco27155, w_eco27156, w_eco27157, w_eco27158, w_eco27159, w_eco27160, w_eco27161, w_eco27162, w_eco27163, w_eco27164, w_eco27165, w_eco27166, w_eco27167, w_eco27168, w_eco27169, w_eco27170, w_eco27171, w_eco27172, w_eco27173, w_eco27174, w_eco27175, w_eco27176, w_eco27177, w_eco27178, w_eco27179, w_eco27180, w_eco27181, w_eco27182, w_eco27183, w_eco27184, w_eco27185, w_eco27186, w_eco27187, w_eco27188, w_eco27189, w_eco27190, w_eco27191, w_eco27192, w_eco27193, w_eco27194, w_eco27195, w_eco27196, w_eco27197, w_eco27198, w_eco27199, w_eco27200, w_eco27201, w_eco27202, w_eco27203, w_eco27204, w_eco27205, w_eco27206, w_eco27207, w_eco27208, w_eco27209, w_eco27210, w_eco27211, w_eco27212, w_eco27213, w_eco27214, w_eco27215, w_eco27216, w_eco27217, w_eco27218, w_eco27219, w_eco27220, w_eco27221, w_eco27222, w_eco27223, w_eco27224, w_eco27225, w_eco27226, w_eco27227, w_eco27228, w_eco27229, w_eco27230, w_eco27231, w_eco27232, w_eco27233, w_eco27234, w_eco27235, w_eco27236, w_eco27237, w_eco27238, w_eco27239, w_eco27240, w_eco27241, w_eco27242, w_eco27243, w_eco27244, w_eco27245, w_eco27246, w_eco27247, w_eco27248, w_eco27249, w_eco27250, w_eco27251, w_eco27252, w_eco27253, w_eco27254, w_eco27255, w_eco27256, w_eco27257, w_eco27258, w_eco27259, w_eco27260, w_eco27261, w_eco27262, w_eco27263, w_eco27264, w_eco27265, w_eco27266, w_eco27267, w_eco27268, w_eco27269, w_eco27270, w_eco27271, w_eco27272, w_eco27273, w_eco27274, w_eco27275, w_eco27276, w_eco27277, w_eco27278, w_eco27279, w_eco27280, w_eco27281, w_eco27282, w_eco27283, w_eco27284, w_eco27285, w_eco27286, w_eco27287, w_eco27288, w_eco27289, w_eco27290, w_eco27291, w_eco27292, w_eco27293, w_eco27294, w_eco27295, w_eco27296, w_eco27297, w_eco27298, w_eco27299, w_eco27300, w_eco27301, w_eco27302, w_eco27303, w_eco27304, w_eco27305, w_eco27306, w_eco27307, w_eco27308, w_eco27309, w_eco27310, w_eco27311, w_eco27312, w_eco27313, w_eco27314, w_eco27315, w_eco27316, w_eco27317, w_eco27318, w_eco27319, w_eco27320, w_eco27321, w_eco27322, w_eco27323, w_eco27324, w_eco27325, w_eco27326, w_eco27327, w_eco27328, w_eco27329, w_eco27330, w_eco27331, w_eco27332, w_eco27333, w_eco27334, w_eco27335, w_eco27336, w_eco27337, w_eco27338, w_eco27339, w_eco27340, w_eco27341, w_eco27342, w_eco27343, w_eco27344, w_eco27345, w_eco27346, w_eco27347, w_eco27348, w_eco27349, w_eco27350, w_eco27351, w_eco27352, w_eco27353, w_eco27354, w_eco27355, w_eco27356, w_eco27357, w_eco27358, w_eco27359, w_eco27360, w_eco27361, w_eco27362, w_eco27363, w_eco27364, w_eco27365, w_eco27366, w_eco27367, w_eco27368, w_eco27369, w_eco27370, w_eco27371, w_eco27372, w_eco27373, w_eco27374, w_eco27375, w_eco27376, w_eco27377, w_eco27378, w_eco27379, w_eco27380, w_eco27381, w_eco27382, w_eco27383, w_eco27384, w_eco27385, w_eco27386, w_eco27387, w_eco27388, w_eco27389, w_eco27390, w_eco27391, w_eco27392, w_eco27393, w_eco27394, w_eco27395, w_eco27396, w_eco27397, w_eco27398, w_eco27399, w_eco27400, w_eco27401, w_eco27402, w_eco27403, w_eco27404, w_eco27405, w_eco27406, w_eco27407, w_eco27408, w_eco27409, w_eco27410, w_eco27411, w_eco27412, w_eco27413, w_eco27414, w_eco27415, w_eco27416, w_eco27417, w_eco27418, w_eco27419, w_eco27420, w_eco27421, w_eco27422, w_eco27423, w_eco27424, w_eco27425, w_eco27426, w_eco27427, w_eco27428, w_eco27429, w_eco27430, w_eco27431, w_eco27432, w_eco27433, w_eco27434, w_eco27435, w_eco27436, w_eco27437, w_eco27438, w_eco27439, w_eco27440, w_eco27441, w_eco27442, w_eco27443, w_eco27444, w_eco27445, w_eco27446, w_eco27447, w_eco27448, w_eco27449, w_eco27450, w_eco27451, w_eco27452, w_eco27453, w_eco27454, w_eco27455, w_eco27456, w_eco27457, w_eco27458, w_eco27459, w_eco27460, w_eco27461, w_eco27462, w_eco27463, w_eco27464, w_eco27465, w_eco27466, w_eco27467, w_eco27468, w_eco27469, w_eco27470, w_eco27471, w_eco27472, w_eco27473, w_eco27474, w_eco27475, w_eco27476, w_eco27477, w_eco27478, w_eco27479, w_eco27480, w_eco27481, w_eco27482, w_eco27483, w_eco27484, w_eco27485, w_eco27486, w_eco27487, w_eco27488, w_eco27489, w_eco27490, w_eco27491, w_eco27492, w_eco27493, w_eco27494, w_eco27495, w_eco27496, w_eco27497, w_eco27498, w_eco27499, w_eco27500, w_eco27501, w_eco27502, w_eco27503, w_eco27504, w_eco27505, w_eco27506, w_eco27507, w_eco27508, w_eco27509, w_eco27510, w_eco27511, w_eco27512, w_eco27513, w_eco27514, w_eco27515, w_eco27516, w_eco27517, w_eco27518, w_eco27519, w_eco27520, w_eco27521, w_eco27522, w_eco27523, w_eco27524, w_eco27525, w_eco27526, w_eco27527, w_eco27528, w_eco27529, w_eco27530, w_eco27531, w_eco27532, w_eco27533, w_eco27534, w_eco27535, w_eco27536, w_eco27537, w_eco27538, w_eco27539, w_eco27540, w_eco27541, w_eco27542, w_eco27543, w_eco27544, w_eco27545, w_eco27546, w_eco27547, w_eco27548, w_eco27549, w_eco27550, w_eco27551, w_eco27552, w_eco27553, w_eco27554, w_eco27555, w_eco27556, w_eco27557, w_eco27558, w_eco27559, w_eco27560, w_eco27561, w_eco27562, w_eco27563, w_eco27564, w_eco27565, w_eco27566, w_eco27567, w_eco27568, w_eco27569, w_eco27570, w_eco27571, w_eco27572, w_eco27573, w_eco27574, w_eco27575, w_eco27576, w_eco27577, w_eco27578, w_eco27579, w_eco27580, w_eco27581, w_eco27582, w_eco27583, w_eco27584, w_eco27585, w_eco27586, w_eco27587, w_eco27588, w_eco27589, w_eco27590, w_eco27591, w_eco27592, w_eco27593, w_eco27594, w_eco27595, w_eco27596, w_eco27597, w_eco27598, w_eco27599, w_eco27600, w_eco27601, w_eco27602, w_eco27603, w_eco27604, w_eco27605, w_eco27606, w_eco27607, w_eco27608, w_eco27609, w_eco27610, w_eco27611, w_eco27612, w_eco27613, w_eco27614, w_eco27615, w_eco27616, w_eco27617, w_eco27618, w_eco27619, w_eco27620, w_eco27621, w_eco27622, w_eco27623, w_eco27624, w_eco27625, w_eco27626, w_eco27627, w_eco27628, w_eco27629, w_eco27630, w_eco27631, w_eco27632, w_eco27633, w_eco27634, w_eco27635, w_eco27636, w_eco27637, w_eco27638, w_eco27639, w_eco27640, w_eco27641, w_eco27642, w_eco27643, w_eco27644, w_eco27645, w_eco27646, w_eco27647, w_eco27648, w_eco27649, w_eco27650, w_eco27651, w_eco27652, w_eco27653, w_eco27654, w_eco27655, w_eco27656, w_eco27657, w_eco27658, w_eco27659, w_eco27660, w_eco27661, w_eco27662, w_eco27663, w_eco27664, w_eco27665, w_eco27666, w_eco27667, w_eco27668, w_eco27669, w_eco27670, w_eco27671, w_eco27672, w_eco27673, w_eco27674, w_eco27675, w_eco27676, w_eco27677, w_eco27678, w_eco27679, w_eco27680, w_eco27681, w_eco27682, w_eco27683, w_eco27684, w_eco27685, w_eco27686, w_eco27687, w_eco27688, w_eco27689, w_eco27690, w_eco27691, w_eco27692, w_eco27693, w_eco27694, w_eco27695, w_eco27696, w_eco27697, w_eco27698, w_eco27699, w_eco27700, w_eco27701, w_eco27702, w_eco27703, w_eco27704, w_eco27705, w_eco27706, w_eco27707, w_eco27708, w_eco27709, w_eco27710, w_eco27711, w_eco27712, w_eco27713, w_eco27714, w_eco27715, w_eco27716, w_eco27717, w_eco27718, w_eco27719, w_eco27720, w_eco27721, w_eco27722, w_eco27723, w_eco27724, w_eco27725, w_eco27726, w_eco27727, w_eco27728, w_eco27729, w_eco27730, w_eco27731, w_eco27732, w_eco27733, w_eco27734, w_eco27735, w_eco27736, w_eco27737, w_eco27738, w_eco27739, w_eco27740, w_eco27741, w_eco27742, w_eco27743, w_eco27744, w_eco27745, w_eco27746, w_eco27747, w_eco27748, w_eco27749, w_eco27750, w_eco27751, w_eco27752, w_eco27753, w_eco27754, w_eco27755, w_eco27756, w_eco27757, w_eco27758, w_eco27759, w_eco27760, w_eco27761, w_eco27762, w_eco27763, w_eco27764, w_eco27765, w_eco27766, w_eco27767, w_eco27768, w_eco27769, w_eco27770, w_eco27771, w_eco27772, w_eco27773, w_eco27774, w_eco27775, w_eco27776, w_eco27777, w_eco27778, w_eco27779, w_eco27780, w_eco27781, w_eco27782, w_eco27783, w_eco27784, w_eco27785, w_eco27786, w_eco27787, w_eco27788, w_eco27789, w_eco27790, w_eco27791, w_eco27792, w_eco27793, w_eco27794, w_eco27795, w_eco27796, w_eco27797, w_eco27798, w_eco27799, w_eco27800, w_eco27801, w_eco27802, w_eco27803, w_eco27804, w_eco27805, w_eco27806, w_eco27807, w_eco27808, w_eco27809, w_eco27810, w_eco27811, w_eco27812, w_eco27813, w_eco27814, w_eco27815, w_eco27816, w_eco27817, w_eco27818, w_eco27819, w_eco27820, w_eco27821, w_eco27822, w_eco27823, w_eco27824, w_eco27825, w_eco27826, w_eco27827, w_eco27828, w_eco27829, w_eco27830, w_eco27831, w_eco27832, w_eco27833, w_eco27834, w_eco27835, w_eco27836, w_eco27837, w_eco27838, w_eco27839, w_eco27840, w_eco27841, w_eco27842, w_eco27843, w_eco27844, w_eco27845, w_eco27846, w_eco27847, w_eco27848, w_eco27849, w_eco27850, w_eco27851, w_eco27852, w_eco27853, w_eco27854, w_eco27855, w_eco27856, w_eco27857, w_eco27858, w_eco27859, w_eco27860, w_eco27861, w_eco27862, w_eco27863, w_eco27864, w_eco27865, w_eco27866, w_eco27867, w_eco27868, w_eco27869, w_eco27870, w_eco27871, w_eco27872, w_eco27873, w_eco27874, w_eco27875, w_eco27876, w_eco27877, w_eco27878, w_eco27879, w_eco27880, w_eco27881, w_eco27882, w_eco27883, w_eco27884, w_eco27885, w_eco27886, w_eco27887, w_eco27888, w_eco27889, w_eco27890, w_eco27891, w_eco27892, w_eco27893, w_eco27894, w_eco27895, w_eco27896, w_eco27897, w_eco27898, w_eco27899, w_eco27900, w_eco27901, w_eco27902, w_eco27903, w_eco27904, w_eco27905, w_eco27906, w_eco27907, w_eco27908, w_eco27909, w_eco27910, w_eco27911, w_eco27912, w_eco27913, w_eco27914, w_eco27915, w_eco27916, w_eco27917, w_eco27918, w_eco27919, w_eco27920, w_eco27921, w_eco27922, w_eco27923, w_eco27924, w_eco27925, w_eco27926, w_eco27927, w_eco27928, w_eco27929, w_eco27930, w_eco27931, w_eco27932, w_eco27933, w_eco27934, w_eco27935, w_eco27936, w_eco27937, w_eco27938, w_eco27939, w_eco27940, w_eco27941, w_eco27942, w_eco27943, w_eco27944, w_eco27945, w_eco27946, w_eco27947, w_eco27948, w_eco27949, w_eco27950, w_eco27951, w_eco27952, w_eco27953, w_eco27954, w_eco27955, w_eco27956, w_eco27957, w_eco27958, w_eco27959, w_eco27960, w_eco27961, w_eco27962, w_eco27963, w_eco27964, w_eco27965, w_eco27966, w_eco27967, w_eco27968, w_eco27969, w_eco27970, w_eco27971, w_eco27972, w_eco27973, w_eco27974, w_eco27975, w_eco27976, w_eco27977, w_eco27978, w_eco27979, w_eco27980, w_eco27981, w_eco27982, w_eco27983, w_eco27984, w_eco27985, w_eco27986, w_eco27987, w_eco27988, w_eco27989, w_eco27990, w_eco27991, w_eco27992, w_eco27993, w_eco27994, w_eco27995, w_eco27996, w_eco27997, w_eco27998, w_eco27999, w_eco28000, w_eco28001, w_eco28002, w_eco28003, w_eco28004, w_eco28005, w_eco28006, w_eco28007, w_eco28008, w_eco28009, w_eco28010, w_eco28011, w_eco28012, w_eco28013, w_eco28014, w_eco28015, w_eco28016, w_eco28017, w_eco28018, w_eco28019, w_eco28020, w_eco28021, w_eco28022, w_eco28023, w_eco28024, w_eco28025, w_eco28026, w_eco28027, w_eco28028, w_eco28029, w_eco28030, w_eco28031, w_eco28032, w_eco28033, w_eco28034, w_eco28035, w_eco28036, w_eco28037, w_eco28038, w_eco28039, w_eco28040, w_eco28041, w_eco28042, w_eco28043, w_eco28044, w_eco28045, w_eco28046, w_eco28047, w_eco28048, w_eco28049, w_eco28050, w_eco28051, w_eco28052, w_eco28053, w_eco28054, w_eco28055, w_eco28056, w_eco28057, w_eco28058, w_eco28059, w_eco28060, w_eco28061, w_eco28062, w_eco28063, w_eco28064, w_eco28065, w_eco28066, w_eco28067, w_eco28068, w_eco28069, w_eco28070, w_eco28071, w_eco28072, w_eco28073, w_eco28074, w_eco28075, w_eco28076, w_eco28077, w_eco28078, w_eco28079, w_eco28080, w_eco28081, w_eco28082, w_eco28083, w_eco28084, w_eco28085, w_eco28086, w_eco28087, w_eco28088, w_eco28089, w_eco28090, w_eco28091, w_eco28092, w_eco28093, w_eco28094, w_eco28095, w_eco28096, w_eco28097, w_eco28098, w_eco28099, w_eco28100, w_eco28101, w_eco28102, w_eco28103, w_eco28104, w_eco28105, w_eco28106, w_eco28107, w_eco28108, w_eco28109, w_eco28110, w_eco28111, w_eco28112, w_eco28113, w_eco28114, w_eco28115, w_eco28116, w_eco28117, w_eco28118, w_eco28119, w_eco28120, w_eco28121, w_eco28122, w_eco28123, w_eco28124, w_eco28125, w_eco28126, w_eco28127, w_eco28128, w_eco28129, w_eco28130, w_eco28131, w_eco28132, w_eco28133, w_eco28134, w_eco28135, w_eco28136, w_eco28137, w_eco28138, w_eco28139, w_eco28140, w_eco28141, w_eco28142, w_eco28143, w_eco28144, w_eco28145, w_eco28146, w_eco28147, w_eco28148, w_eco28149, w_eco28150, w_eco28151, w_eco28152, w_eco28153, w_eco28154, w_eco28155, w_eco28156, w_eco28157, w_eco28158, w_eco28159, w_eco28160, w_eco28161, w_eco28162, w_eco28163, w_eco28164, w_eco28165, w_eco28166, w_eco28167, w_eco28168, w_eco28169, w_eco28170, w_eco28171, w_eco28172, w_eco28173, w_eco28174, w_eco28175, w_eco28176, w_eco28177, w_eco28178, w_eco28179, w_eco28180, w_eco28181, w_eco28182, w_eco28183, w_eco28184, w_eco28185, w_eco28186, w_eco28187, w_eco28188, w_eco28189, w_eco28190, w_eco28191, w_eco28192, w_eco28193, w_eco28194, w_eco28195, w_eco28196, w_eco28197, w_eco28198, w_eco28199, w_eco28200, w_eco28201, w_eco28202, w_eco28203, w_eco28204, w_eco28205, w_eco28206, w_eco28207, w_eco28208, w_eco28209, w_eco28210, w_eco28211, w_eco28212, w_eco28213, w_eco28214, w_eco28215, w_eco28216, w_eco28217, w_eco28218, w_eco28219, w_eco28220, w_eco28221, w_eco28222, w_eco28223, w_eco28224, w_eco28225, w_eco28226, w_eco28227, w_eco28228, w_eco28229, w_eco28230, w_eco28231, w_eco28232, w_eco28233, w_eco28234, w_eco28235, w_eco28236, w_eco28237, w_eco28238, w_eco28239, w_eco28240, w_eco28241, w_eco28242, w_eco28243, w_eco28244, w_eco28245, w_eco28246, w_eco28247, w_eco28248, w_eco28249, w_eco28250, w_eco28251, w_eco28252, w_eco28253, w_eco28254, w_eco28255, w_eco28256, w_eco28257, w_eco28258, w_eco28259, w_eco28260, w_eco28261, w_eco28262, w_eco28263, w_eco28264, w_eco28265, w_eco28266, w_eco28267, w_eco28268, w_eco28269, w_eco28270, w_eco28271, w_eco28272, w_eco28273, w_eco28274, w_eco28275, w_eco28276, w_eco28277, w_eco28278, w_eco28279, w_eco28280, w_eco28281, w_eco28282, w_eco28283, w_eco28284, w_eco28285, w_eco28286, w_eco28287, w_eco28288, w_eco28289, w_eco28290, w_eco28291, w_eco28292, w_eco28293, w_eco28294, w_eco28295, w_eco28296, w_eco28297, w_eco28298, w_eco28299, w_eco28300, w_eco28301, w_eco28302, w_eco28303, w_eco28304, w_eco28305, w_eco28306, w_eco28307, w_eco28308, w_eco28309, w_eco28310, w_eco28311, w_eco28312, w_eco28313, w_eco28314, w_eco28315, w_eco28316, w_eco28317, w_eco28318, w_eco28319, w_eco28320, w_eco28321, w_eco28322, w_eco28323, w_eco28324, w_eco28325, w_eco28326, w_eco28327, w_eco28328, w_eco28329, w_eco28330, w_eco28331, w_eco28332, w_eco28333, w_eco28334, w_eco28335, w_eco28336, w_eco28337, w_eco28338, w_eco28339, w_eco28340, w_eco28341, w_eco28342, w_eco28343, w_eco28344, w_eco28345, w_eco28346, w_eco28347, w_eco28348, w_eco28349, w_eco28350, w_eco28351, w_eco28352, w_eco28353, w_eco28354, w_eco28355, w_eco28356, w_eco28357, w_eco28358, w_eco28359, w_eco28360, w_eco28361, w_eco28362, w_eco28363, w_eco28364, w_eco28365, w_eco28366, w_eco28367, w_eco28368, w_eco28369, w_eco28370, w_eco28371, w_eco28372, w_eco28373, w_eco28374, w_eco28375, w_eco28376, w_eco28377, w_eco28378, w_eco28379, w_eco28380, w_eco28381, w_eco28382, w_eco28383, w_eco28384, w_eco28385, w_eco28386, w_eco28387, w_eco28388, w_eco28389, w_eco28390, w_eco28391, w_eco28392, w_eco28393, w_eco28394, w_eco28395, w_eco28396, w_eco28397, w_eco28398, w_eco28399, w_eco28400, w_eco28401, w_eco28402, w_eco28403, w_eco28404, w_eco28405, w_eco28406, w_eco28407, w_eco28408, w_eco28409, w_eco28410, w_eco28411, w_eco28412, w_eco28413, w_eco28414, w_eco28415, w_eco28416, w_eco28417, w_eco28418, w_eco28419, w_eco28420, w_eco28421, w_eco28422, w_eco28423, w_eco28424, w_eco28425, w_eco28426, w_eco28427, w_eco28428, w_eco28429, w_eco28430, w_eco28431, w_eco28432, w_eco28433, w_eco28434, w_eco28435, w_eco28436, w_eco28437, w_eco28438, w_eco28439, w_eco28440, w_eco28441, w_eco28442, w_eco28443, w_eco28444, w_eco28445, w_eco28446, w_eco28447, w_eco28448, w_eco28449, w_eco28450, w_eco28451, w_eco28452, w_eco28453, w_eco28454, w_eco28455, w_eco28456, w_eco28457, w_eco28458, w_eco28459, w_eco28460, w_eco28461, w_eco28462, w_eco28463, w_eco28464, w_eco28465, w_eco28466, w_eco28467, w_eco28468, w_eco28469, w_eco28470, w_eco28471, w_eco28472, w_eco28473, w_eco28474, w_eco28475, w_eco28476, w_eco28477, w_eco28478, w_eco28479, w_eco28480, w_eco28481, w_eco28482, w_eco28483, w_eco28484, w_eco28485, w_eco28486, w_eco28487, w_eco28488, w_eco28489, w_eco28490, w_eco28491, w_eco28492, w_eco28493, w_eco28494, w_eco28495, w_eco28496, w_eco28497, w_eco28498, w_eco28499, w_eco28500, w_eco28501, w_eco28502, w_eco28503, w_eco28504, w_eco28505, w_eco28506, w_eco28507, w_eco28508, w_eco28509, w_eco28510, w_eco28511, w_eco28512, w_eco28513, w_eco28514, w_eco28515, w_eco28516, w_eco28517, w_eco28518, w_eco28519, w_eco28520, w_eco28521, w_eco28522, w_eco28523, w_eco28524, w_eco28525, w_eco28526, w_eco28527, w_eco28528, w_eco28529, w_eco28530, w_eco28531, w_eco28532, w_eco28533, w_eco28534, w_eco28535, w_eco28536, w_eco28537, w_eco28538, w_eco28539, w_eco28540, w_eco28541, w_eco28542, w_eco28543, w_eco28544, w_eco28545, w_eco28546, w_eco28547, w_eco28548, w_eco28549, w_eco28550, w_eco28551, w_eco28552, w_eco28553, w_eco28554, w_eco28555, w_eco28556, w_eco28557, w_eco28558, w_eco28559, w_eco28560, w_eco28561, w_eco28562, w_eco28563, w_eco28564, w_eco28565, w_eco28566, w_eco28567, w_eco28568, w_eco28569, w_eco28570, w_eco28571, w_eco28572, w_eco28573, w_eco28574, w_eco28575, w_eco28576, w_eco28577, w_eco28578, w_eco28579, w_eco28580, w_eco28581, w_eco28582, w_eco28583, w_eco28584, w_eco28585, w_eco28586, w_eco28587, w_eco28588, w_eco28589, w_eco28590, w_eco28591, w_eco28592, w_eco28593, w_eco28594, w_eco28595, w_eco28596, w_eco28597, w_eco28598, w_eco28599, w_eco28600, w_eco28601, w_eco28602, w_eco28603, w_eco28604, w_eco28605, w_eco28606, w_eco28607, w_eco28608, w_eco28609, w_eco28610, w_eco28611, w_eco28612, w_eco28613, w_eco28614, w_eco28615, w_eco28616, w_eco28617, w_eco28618, w_eco28619, w_eco28620, w_eco28621, w_eco28622, w_eco28623, w_eco28624, w_eco28625, w_eco28626, w_eco28627, w_eco28628, w_eco28629, w_eco28630, w_eco28631, w_eco28632, w_eco28633, w_eco28634, w_eco28635, w_eco28636, w_eco28637, w_eco28638, w_eco28639, w_eco28640, w_eco28641, w_eco28642, w_eco28643, w_eco28644, w_eco28645, w_eco28646, w_eco28647, w_eco28648, w_eco28649, w_eco28650, w_eco28651, w_eco28652, w_eco28653, w_eco28654, w_eco28655, w_eco28656, w_eco28657, w_eco28658, w_eco28659, w_eco28660, w_eco28661, w_eco28662, w_eco28663, w_eco28664, w_eco28665, w_eco28666, w_eco28667, w_eco28668, w_eco28669, w_eco28670, w_eco28671, w_eco28672, w_eco28673, w_eco28674, w_eco28675, w_eco28676, w_eco28677, w_eco28678, w_eco28679, w_eco28680, w_eco28681, w_eco28682, w_eco28683, w_eco28684, w_eco28685, w_eco28686, w_eco28687, w_eco28688, w_eco28689, w_eco28690, w_eco28691, w_eco28692, w_eco28693, w_eco28694, w_eco28695, w_eco28696, w_eco28697, w_eco28698, w_eco28699, w_eco28700, w_eco28701, w_eco28702, w_eco28703, w_eco28704, w_eco28705, w_eco28706, w_eco28707, w_eco28708, w_eco28709, w_eco28710, w_eco28711, w_eco28712, w_eco28713, w_eco28714, w_eco28715, w_eco28716, w_eco28717, w_eco28718, w_eco28719, w_eco28720, w_eco28721, w_eco28722, w_eco28723, w_eco28724, w_eco28725, w_eco28726, w_eco28727, w_eco28728, w_eco28729, w_eco28730, w_eco28731, w_eco28732, w_eco28733, w_eco28734, w_eco28735, w_eco28736, w_eco28737, w_eco28738, w_eco28739, w_eco28740, w_eco28741, w_eco28742, w_eco28743, w_eco28744, w_eco28745, w_eco28746, w_eco28747, w_eco28748, w_eco28749, w_eco28750, w_eco28751, w_eco28752, w_eco28753, w_eco28754, w_eco28755, w_eco28756, w_eco28757, w_eco28758, w_eco28759, w_eco28760, w_eco28761, w_eco28762, w_eco28763, w_eco28764, w_eco28765, w_eco28766, w_eco28767, w_eco28768, w_eco28769, w_eco28770, w_eco28771, w_eco28772, w_eco28773, w_eco28774, w_eco28775, w_eco28776, w_eco28777, w_eco28778, w_eco28779, w_eco28780, w_eco28781, w_eco28782, w_eco28783, w_eco28784, w_eco28785, w_eco28786, w_eco28787, w_eco28788, w_eco28789, w_eco28790, w_eco28791, w_eco28792, w_eco28793, w_eco28794, w_eco28795, w_eco28796, w_eco28797, w_eco28798, w_eco28799, w_eco28800, w_eco28801, w_eco28802, w_eco28803, w_eco28804, w_eco28805, w_eco28806, w_eco28807, w_eco28808, w_eco28809, w_eco28810, w_eco28811, w_eco28812, w_eco28813, w_eco28814, w_eco28815, w_eco28816, w_eco28817, w_eco28818, w_eco28819, w_eco28820, w_eco28821, w_eco28822, w_eco28823, w_eco28824, w_eco28825, w_eco28826, w_eco28827, w_eco28828, w_eco28829, w_eco28830, w_eco28831, w_eco28832, w_eco28833, w_eco28834, w_eco28835, w_eco28836, w_eco28837, w_eco28838, w_eco28839, w_eco28840, w_eco28841, w_eco28842, w_eco28843, w_eco28844, w_eco28845, w_eco28846, w_eco28847, w_eco28848, w_eco28849, w_eco28850, w_eco28851, w_eco28852, w_eco28853, w_eco28854, w_eco28855, w_eco28856, w_eco28857, w_eco28858, w_eco28859, w_eco28860, w_eco28861, w_eco28862, w_eco28863, w_eco28864, w_eco28865, w_eco28866, w_eco28867, w_eco28868, w_eco28869, w_eco28870, w_eco28871, w_eco28872, w_eco28873, w_eco28874, w_eco28875, w_eco28876, w_eco28877, w_eco28878, w_eco28879, w_eco28880, w_eco28881, w_eco28882, w_eco28883, w_eco28884, w_eco28885, w_eco28886, w_eco28887, w_eco28888, w_eco28889, w_eco28890, w_eco28891, w_eco28892, w_eco28893, w_eco28894, w_eco28895, w_eco28896, w_eco28897, w_eco28898, w_eco28899, w_eco28900, w_eco28901, w_eco28902, w_eco28903, w_eco28904, w_eco28905, w_eco28906, w_eco28907, w_eco28908, w_eco28909, w_eco28910, w_eco28911, w_eco28912, w_eco28913, w_eco28914, w_eco28915, w_eco28916, w_eco28917, w_eco28918, w_eco28919, w_eco28920, w_eco28921, w_eco28922, w_eco28923, w_eco28924, w_eco28925, w_eco28926, w_eco28927, w_eco28928, w_eco28929, w_eco28930, w_eco28931, w_eco28932, w_eco28933, w_eco28934, w_eco28935, w_eco28936, w_eco28937, w_eco28938, w_eco28939, w_eco28940, w_eco28941, w_eco28942, w_eco28943, w_eco28944, w_eco28945, w_eco28946, w_eco28947, w_eco28948, w_eco28949, w_eco28950, w_eco28951, w_eco28952, w_eco28953, w_eco28954, w_eco28955, w_eco28956, w_eco28957, w_eco28958, w_eco28959, w_eco28960, w_eco28961, w_eco28962, w_eco28963, w_eco28964, w_eco28965, w_eco28966, w_eco28967, w_eco28968, w_eco28969, w_eco28970, w_eco28971, w_eco28972, w_eco28973, w_eco28974, w_eco28975, w_eco28976, w_eco28977, w_eco28978, w_eco28979, w_eco28980, w_eco28981, w_eco28982, w_eco28983, w_eco28984, w_eco28985, w_eco28986, w_eco28987, w_eco28988, w_eco28989, w_eco28990, w_eco28991, w_eco28992, w_eco28993, w_eco28994, w_eco28995, w_eco28996, w_eco28997, w_eco28998, w_eco28999, w_eco29000, w_eco29001, w_eco29002, w_eco29003, w_eco29004, w_eco29005, w_eco29006, w_eco29007, w_eco29008, w_eco29009, w_eco29010, w_eco29011, w_eco29012, w_eco29013, w_eco29014, w_eco29015, w_eco29016, w_eco29017, w_eco29018, w_eco29019, w_eco29020, w_eco29021, w_eco29022, w_eco29023, w_eco29024, w_eco29025, w_eco29026, w_eco29027, w_eco29028, w_eco29029, w_eco29030, w_eco29031, w_eco29032, w_eco29033, w_eco29034, w_eco29035, w_eco29036, w_eco29037, w_eco29038, w_eco29039, w_eco29040, w_eco29041, w_eco29042, w_eco29043, w_eco29044, w_eco29045, w_eco29046, w_eco29047, w_eco29048, w_eco29049, w_eco29050, w_eco29051, w_eco29052, w_eco29053, w_eco29054, w_eco29055, w_eco29056, w_eco29057, w_eco29058, w_eco29059, w_eco29060, w_eco29061, w_eco29062, w_eco29063, w_eco29064, w_eco29065, w_eco29066, w_eco29067, w_eco29068, w_eco29069, w_eco29070, w_eco29071, w_eco29072, w_eco29073, w_eco29074, w_eco29075, w_eco29076, w_eco29077, w_eco29078, w_eco29079, w_eco29080, w_eco29081, w_eco29082, w_eco29083, w_eco29084, w_eco29085, w_eco29086, w_eco29087, w_eco29088, w_eco29089, w_eco29090, w_eco29091, w_eco29092, w_eco29093, w_eco29094, w_eco29095, w_eco29096, w_eco29097, w_eco29098, w_eco29099, w_eco29100, w_eco29101, w_eco29102, w_eco29103, w_eco29104, w_eco29105, w_eco29106, w_eco29107, w_eco29108, w_eco29109, w_eco29110, w_eco29111, w_eco29112, w_eco29113, w_eco29114, w_eco29115, w_eco29116, w_eco29117, w_eco29118, w_eco29119, w_eco29120, w_eco29121, w_eco29122, w_eco29123, w_eco29124, w_eco29125, w_eco29126, w_eco29127, w_eco29128, w_eco29129, w_eco29130, w_eco29131, w_eco29132, w_eco29133, w_eco29134, w_eco29135, w_eco29136, w_eco29137, w_eco29138, w_eco29139, w_eco29140, w_eco29141, w_eco29142, w_eco29143, w_eco29144, w_eco29145, w_eco29146, w_eco29147, w_eco29148, w_eco29149, w_eco29150, w_eco29151, w_eco29152, w_eco29153, w_eco29154, w_eco29155, w_eco29156, w_eco29157, w_eco29158, w_eco29159, w_eco29160, w_eco29161, w_eco29162, w_eco29163, w_eco29164, w_eco29165, w_eco29166, w_eco29167, w_eco29168, w_eco29169, w_eco29170, w_eco29171, w_eco29172, w_eco29173, w_eco29174, w_eco29175, w_eco29176, w_eco29177, w_eco29178, w_eco29179, w_eco29180, w_eco29181, w_eco29182, w_eco29183, w_eco29184, w_eco29185, w_eco29186, w_eco29187, w_eco29188, w_eco29189, w_eco29190, w_eco29191, w_eco29192, w_eco29193, w_eco29194, w_eco29195, w_eco29196, w_eco29197, w_eco29198, w_eco29199, w_eco29200, w_eco29201, w_eco29202, w_eco29203, w_eco29204, w_eco29205, w_eco29206, w_eco29207, w_eco29208, w_eco29209, w_eco29210, w_eco29211, w_eco29212, w_eco29213, w_eco29214, w_eco29215, w_eco29216, w_eco29217, w_eco29218, w_eco29219, w_eco29220, w_eco29221, w_eco29222, w_eco29223, w_eco29224, w_eco29225, w_eco29226, w_eco29227, w_eco29228, w_eco29229, w_eco29230, w_eco29231, w_eco29232, w_eco29233, w_eco29234, w_eco29235, w_eco29236, w_eco29237, w_eco29238, w_eco29239, w_eco29240, w_eco29241, w_eco29242, w_eco29243, w_eco29244, w_eco29245, w_eco29246, w_eco29247, w_eco29248, w_eco29249, w_eco29250, w_eco29251, w_eco29252, w_eco29253, w_eco29254, w_eco29255, w_eco29256, w_eco29257, w_eco29258, w_eco29259, w_eco29260, w_eco29261, w_eco29262, w_eco29263, w_eco29264, w_eco29265, w_eco29266, w_eco29267, w_eco29268, w_eco29269, w_eco29270, w_eco29271, w_eco29272, w_eco29273, w_eco29274, w_eco29275, w_eco29276, w_eco29277, w_eco29278, w_eco29279, w_eco29280, w_eco29281, w_eco29282, w_eco29283, w_eco29284, w_eco29285, w_eco29286, w_eco29287, w_eco29288, w_eco29289, w_eco29290, w_eco29291, w_eco29292, w_eco29293, w_eco29294, w_eco29295, w_eco29296, w_eco29297, w_eco29298, w_eco29299, w_eco29300, w_eco29301, w_eco29302, w_eco29303, w_eco29304, w_eco29305, w_eco29306, w_eco29307, w_eco29308, w_eco29309, w_eco29310, w_eco29311, w_eco29312, w_eco29313, w_eco29314, w_eco29315, w_eco29316, w_eco29317, w_eco29318, w_eco29319, w_eco29320, w_eco29321, w_eco29322, w_eco29323, w_eco29324, w_eco29325, w_eco29326, w_eco29327, w_eco29328, w_eco29329, w_eco29330, w_eco29331, w_eco29332, w_eco29333, w_eco29334, w_eco29335, w_eco29336, w_eco29337, w_eco29338, w_eco29339, w_eco29340, w_eco29341, w_eco29342, w_eco29343, w_eco29344, w_eco29345, w_eco29346, w_eco29347, w_eco29348, w_eco29349, w_eco29350, w_eco29351, w_eco29352, w_eco29353, w_eco29354, w_eco29355, w_eco29356, w_eco29357, w_eco29358, w_eco29359, w_eco29360, w_eco29361, w_eco29362, w_eco29363, w_eco29364, w_eco29365, w_eco29366, w_eco29367, w_eco29368, w_eco29369, w_eco29370, w_eco29371, w_eco29372, w_eco29373, w_eco29374, w_eco29375, w_eco29376, w_eco29377, w_eco29378, w_eco29379, w_eco29380, w_eco29381, w_eco29382, w_eco29383, w_eco29384, w_eco29385, w_eco29386, w_eco29387, w_eco29388, w_eco29389, w_eco29390, w_eco29391, w_eco29392, w_eco29393, w_eco29394, w_eco29395, w_eco29396, w_eco29397, w_eco29398, w_eco29399, w_eco29400, w_eco29401, w_eco29402, w_eco29403, w_eco29404, w_eco29405, w_eco29406, w_eco29407, w_eco29408, w_eco29409, w_eco29410, w_eco29411, w_eco29412, w_eco29413, w_eco29414, w_eco29415, w_eco29416, w_eco29417, w_eco29418, w_eco29419, w_eco29420, w_eco29421, w_eco29422, w_eco29423, w_eco29424, w_eco29425, w_eco29426, w_eco29427, w_eco29428, w_eco29429, w_eco29430, w_eco29431, w_eco29432, w_eco29433, w_eco29434, w_eco29435, w_eco29436, w_eco29437, w_eco29438, w_eco29439, w_eco29440, w_eco29441, w_eco29442, w_eco29443, w_eco29444, w_eco29445, w_eco29446, w_eco29447, w_eco29448, w_eco29449, w_eco29450, w_eco29451, w_eco29452, w_eco29453, w_eco29454, w_eco29455, w_eco29456, w_eco29457, w_eco29458, w_eco29459, w_eco29460, w_eco29461, w_eco29462, w_eco29463, w_eco29464, w_eco29465, w_eco29466, w_eco29467, w_eco29468, w_eco29469, w_eco29470, w_eco29471, w_eco29472, w_eco29473, w_eco29474, w_eco29475, w_eco29476, w_eco29477, w_eco29478, w_eco29479, w_eco29480, w_eco29481, w_eco29482, w_eco29483, w_eco29484, w_eco29485, w_eco29486, w_eco29487, w_eco29488, w_eco29489, w_eco29490, w_eco29491, w_eco29492, w_eco29493, w_eco29494, w_eco29495, w_eco29496, w_eco29497, w_eco29498, w_eco29499, w_eco29500, w_eco29501, w_eco29502, w_eco29503, w_eco29504, w_eco29505, w_eco29506, w_eco29507, w_eco29508, w_eco29509, w_eco29510, w_eco29511, w_eco29512, w_eco29513, w_eco29514, w_eco29515, w_eco29516, w_eco29517, w_eco29518, w_eco29519, w_eco29520, w_eco29521, w_eco29522, w_eco29523, w_eco29524, w_eco29525, w_eco29526, w_eco29527, w_eco29528, w_eco29529, w_eco29530, w_eco29531, w_eco29532, w_eco29533, w_eco29534, w_eco29535, w_eco29536, w_eco29537, w_eco29538, w_eco29539, w_eco29540, w_eco29541, w_eco29542, w_eco29543, w_eco29544, w_eco29545, w_eco29546, w_eco29547, w_eco29548, w_eco29549, w_eco29550, w_eco29551, w_eco29552, w_eco29553, w_eco29554, w_eco29555, w_eco29556, w_eco29557, w_eco29558, w_eco29559, w_eco29560, w_eco29561, w_eco29562, w_eco29563, w_eco29564, w_eco29565, w_eco29566, w_eco29567, w_eco29568, w_eco29569, w_eco29570, w_eco29571, w_eco29572, w_eco29573, w_eco29574, w_eco29575, w_eco29576, w_eco29577, w_eco29578, w_eco29579, w_eco29580, w_eco29581, w_eco29582, w_eco29583, w_eco29584, w_eco29585, w_eco29586, w_eco29587, w_eco29588, w_eco29589, w_eco29590, w_eco29591, w_eco29592, w_eco29593, w_eco29594, w_eco29595, w_eco29596, w_eco29597, w_eco29598, w_eco29599, w_eco29600, w_eco29601, w_eco29602, w_eco29603, w_eco29604, w_eco29605, w_eco29606, w_eco29607, w_eco29608, w_eco29609, w_eco29610, w_eco29611, w_eco29612, w_eco29613, w_eco29614, w_eco29615, w_eco29616, w_eco29617, w_eco29618, w_eco29619, w_eco29620, w_eco29621, w_eco29622, w_eco29623, w_eco29624, w_eco29625, w_eco29626, w_eco29627, w_eco29628, w_eco29629, w_eco29630, w_eco29631, w_eco29632, w_eco29633, w_eco29634, w_eco29635, w_eco29636, w_eco29637, w_eco29638, w_eco29639, w_eco29640, w_eco29641, w_eco29642, w_eco29643, w_eco29644, w_eco29645, w_eco29646, w_eco29647, w_eco29648, w_eco29649, w_eco29650, w_eco29651, w_eco29652, w_eco29653, w_eco29654, w_eco29655, w_eco29656, w_eco29657, w_eco29658, w_eco29659, w_eco29660, w_eco29661, w_eco29662, w_eco29663, w_eco29664, w_eco29665, w_eco29666, w_eco29667, w_eco29668, w_eco29669, w_eco29670, w_eco29671, w_eco29672, w_eco29673, w_eco29674, w_eco29675, w_eco29676, w_eco29677, w_eco29678, w_eco29679, w_eco29680, w_eco29681, w_eco29682, w_eco29683, w_eco29684, w_eco29685, w_eco29686, w_eco29687, w_eco29688, w_eco29689, w_eco29690, w_eco29691, w_eco29692, w_eco29693, w_eco29694, w_eco29695, w_eco29696, w_eco29697, w_eco29698, w_eco29699, w_eco29700, w_eco29701, w_eco29702, w_eco29703, w_eco29704, w_eco29705, w_eco29706, w_eco29707, w_eco29708, w_eco29709, w_eco29710, w_eco29711, w_eco29712, w_eco29713, w_eco29714, w_eco29715, w_eco29716, w_eco29717, w_eco29718, w_eco29719, w_eco29720, w_eco29721, w_eco29722, w_eco29723, w_eco29724, w_eco29725, w_eco29726, w_eco29727, w_eco29728, w_eco29729, w_eco29730, w_eco29731, w_eco29732, w_eco29733, w_eco29734, w_eco29735, w_eco29736, w_eco29737, w_eco29738, w_eco29739, w_eco29740, w_eco29741, w_eco29742, w_eco29743, w_eco29744, w_eco29745, w_eco29746, w_eco29747, w_eco29748, w_eco29749, w_eco29750, w_eco29751, w_eco29752, w_eco29753, w_eco29754, w_eco29755, w_eco29756, w_eco29757, w_eco29758, w_eco29759, w_eco29760, w_eco29761, w_eco29762, w_eco29763, w_eco29764, w_eco29765, w_eco29766, w_eco29767, w_eco29768, w_eco29769, w_eco29770, w_eco29771, w_eco29772, w_eco29773, w_eco29774, w_eco29775, w_eco29776, w_eco29777, w_eco29778, w_eco29779, w_eco29780, w_eco29781, w_eco29782, w_eco29783, w_eco29784, w_eco29785, w_eco29786, w_eco29787, w_eco29788, w_eco29789, w_eco29790, w_eco29791, w_eco29792, w_eco29793, w_eco29794, w_eco29795, w_eco29796, w_eco29797, w_eco29798, w_eco29799, w_eco29800, w_eco29801, w_eco29802, w_eco29803, w_eco29804, w_eco29805, w_eco29806, w_eco29807, w_eco29808, w_eco29809, w_eco29810, w_eco29811, w_eco29812, w_eco29813, w_eco29814, w_eco29815, w_eco29816, w_eco29817, w_eco29818, w_eco29819, w_eco29820, w_eco29821, w_eco29822, w_eco29823, w_eco29824, w_eco29825, w_eco29826, w_eco29827, w_eco29828, w_eco29829, w_eco29830, w_eco29831, w_eco29832, w_eco29833, w_eco29834, w_eco29835, w_eco29836, w_eco29837, w_eco29838, w_eco29839, w_eco29840, w_eco29841, w_eco29842, w_eco29843, w_eco29844, w_eco29845, w_eco29846, w_eco29847, w_eco29848, w_eco29849, w_eco29850, w_eco29851, w_eco29852, w_eco29853, w_eco29854, w_eco29855, w_eco29856, w_eco29857, w_eco29858, w_eco29859, w_eco29860, w_eco29861, w_eco29862, w_eco29863, w_eco29864, w_eco29865, w_eco29866, w_eco29867, w_eco29868, w_eco29869, w_eco29870, w_eco29871, w_eco29872, w_eco29873, w_eco29874, w_eco29875, w_eco29876, w_eco29877, w_eco29878, w_eco29879, w_eco29880, w_eco29881, w_eco29882, w_eco29883, w_eco29884, w_eco29885, w_eco29886, w_eco29887, w_eco29888, w_eco29889, w_eco29890, w_eco29891, w_eco29892, w_eco29893, w_eco29894, w_eco29895, w_eco29896, w_eco29897, w_eco29898, w_eco29899, w_eco29900, w_eco29901, w_eco29902, w_eco29903, w_eco29904, w_eco29905, w_eco29906, w_eco29907, w_eco29908, w_eco29909, w_eco29910, w_eco29911, w_eco29912, w_eco29913, w_eco29914, w_eco29915, w_eco29916, w_eco29917, w_eco29918, w_eco29919, w_eco29920, w_eco29921, w_eco29922, w_eco29923, w_eco29924, w_eco29925, w_eco29926, w_eco29927, w_eco29928, w_eco29929, w_eco29930, w_eco29931, w_eco29932, w_eco29933, w_eco29934, w_eco29935, w_eco29936, w_eco29937, w_eco29938, w_eco29939, w_eco29940, w_eco29941, w_eco29942, w_eco29943, w_eco29944, w_eco29945, w_eco29946, w_eco29947, w_eco29948, w_eco29949, w_eco29950, w_eco29951, w_eco29952, w_eco29953, w_eco29954, w_eco29955, w_eco29956, w_eco29957, w_eco29958, w_eco29959, w_eco29960, w_eco29961, w_eco29962, w_eco29963, w_eco29964, w_eco29965, w_eco29966, w_eco29967, w_eco29968, w_eco29969, w_eco29970, w_eco29971, w_eco29972, w_eco29973, w_eco29974, w_eco29975, w_eco29976, w_eco29977, w_eco29978, w_eco29979, w_eco29980, w_eco29981, w_eco29982, w_eco29983, w_eco29984, w_eco29985, w_eco29986, w_eco29987, w_eco29988, w_eco29989, w_eco29990, w_eco29991, w_eco29992, w_eco29993, w_eco29994, w_eco29995, w_eco29996, w_eco29997, w_eco29998, w_eco29999, w_eco30000, w_eco30001, w_eco30002, w_eco30003, w_eco30004, w_eco30005, w_eco30006, w_eco30007, w_eco30008, w_eco30009, w_eco30010, w_eco30011, w_eco30012, w_eco30013, w_eco30014, w_eco30015, w_eco30016, w_eco30017, w_eco30018, w_eco30019, w_eco30020, w_eco30021, w_eco30022, w_eco30023, w_eco30024, w_eco30025, w_eco30026, w_eco30027, w_eco30028, w_eco30029, w_eco30030, w_eco30031, w_eco30032, w_eco30033, w_eco30034, w_eco30035, w_eco30036, w_eco30037, w_eco30038, w_eco30039, w_eco30040, w_eco30041, w_eco30042, w_eco30043, w_eco30044, w_eco30045, w_eco30046, w_eco30047, w_eco30048, w_eco30049, w_eco30050, w_eco30051, w_eco30052, w_eco30053, w_eco30054, w_eco30055, w_eco30056, w_eco30057, w_eco30058, w_eco30059, w_eco30060, w_eco30061, w_eco30062, w_eco30063, w_eco30064, w_eco30065, w_eco30066, w_eco30067, w_eco30068, w_eco30069, w_eco30070, w_eco30071, w_eco30072, w_eco30073, w_eco30074, w_eco30075, w_eco30076, w_eco30077, w_eco30078, w_eco30079, w_eco30080, w_eco30081, w_eco30082, w_eco30083, w_eco30084, w_eco30085, w_eco30086, w_eco30087, w_eco30088, w_eco30089, w_eco30090, w_eco30091, w_eco30092, w_eco30093, w_eco30094, w_eco30095, w_eco30096, w_eco30097, w_eco30098, w_eco30099, w_eco30100, w_eco30101, w_eco30102, w_eco30103, w_eco30104, w_eco30105, w_eco30106, w_eco30107, w_eco30108, w_eco30109, w_eco30110, w_eco30111, w_eco30112, w_eco30113, w_eco30114, w_eco30115, w_eco30116, w_eco30117, w_eco30118, w_eco30119, w_eco30120, w_eco30121, w_eco30122, w_eco30123, w_eco30124, w_eco30125, w_eco30126, w_eco30127, w_eco30128, w_eco30129, w_eco30130, w_eco30131, w_eco30132, w_eco30133, w_eco30134, w_eco30135, w_eco30136, w_eco30137, w_eco30138, w_eco30139, w_eco30140, w_eco30141, w_eco30142, w_eco30143, w_eco30144, w_eco30145, w_eco30146, w_eco30147, w_eco30148, w_eco30149, w_eco30150, w_eco30151, w_eco30152, w_eco30153, w_eco30154, w_eco30155, w_eco30156, w_eco30157, w_eco30158, w_eco30159, w_eco30160, w_eco30161, w_eco30162, w_eco30163, w_eco30164, w_eco30165, w_eco30166, w_eco30167, w_eco30168, w_eco30169, w_eco30170, w_eco30171, w_eco30172, w_eco30173, w_eco30174, w_eco30175, w_eco30176, w_eco30177, w_eco30178, w_eco30179, w_eco30180, w_eco30181, w_eco30182, w_eco30183, w_eco30184, w_eco30185, w_eco30186, w_eco30187, w_eco30188, w_eco30189, w_eco30190, w_eco30191, w_eco30192, w_eco30193, w_eco30194, w_eco30195, w_eco30196, w_eco30197, w_eco30198, w_eco30199, w_eco30200, w_eco30201, w_eco30202, w_eco30203, w_eco30204, w_eco30205, w_eco30206, w_eco30207, w_eco30208, w_eco30209, w_eco30210, w_eco30211, w_eco30212, w_eco30213, w_eco30214, w_eco30215, w_eco30216, w_eco30217, w_eco30218, w_eco30219, w_eco30220, w_eco30221, w_eco30222, w_eco30223, w_eco30224, w_eco30225, w_eco30226, w_eco30227, w_eco30228, w_eco30229, w_eco30230, w_eco30231, w_eco30232, w_eco30233, w_eco30234, w_eco30235, w_eco30236, w_eco30237, w_eco30238, w_eco30239, w_eco30240, w_eco30241, w_eco30242, w_eco30243, w_eco30244, w_eco30245, w_eco30246, w_eco30247, w_eco30248, w_eco30249, w_eco30250, w_eco30251, w_eco30252, w_eco30253, w_eco30254, w_eco30255, w_eco30256, w_eco30257, w_eco30258, w_eco30259, w_eco30260, w_eco30261, w_eco30262, w_eco30263, w_eco30264, w_eco30265, w_eco30266, w_eco30267, w_eco30268, w_eco30269, w_eco30270, w_eco30271, w_eco30272, w_eco30273, w_eco30274, w_eco30275, w_eco30276, w_eco30277, w_eco30278, w_eco30279, w_eco30280, w_eco30281, w_eco30282, w_eco30283, w_eco30284, w_eco30285, w_eco30286, w_eco30287, w_eco30288, w_eco30289, w_eco30290, w_eco30291, w_eco30292, w_eco30293, w_eco30294, w_eco30295, w_eco30296, w_eco30297, w_eco30298, w_eco30299, w_eco30300, w_eco30301, w_eco30302, w_eco30303, w_eco30304, w_eco30305, w_eco30306, w_eco30307, w_eco30308, w_eco30309, w_eco30310, w_eco30311, w_eco30312, w_eco30313, w_eco30314, w_eco30315, w_eco30316, w_eco30317, w_eco30318, w_eco30319, w_eco30320, w_eco30321, w_eco30322, w_eco30323, w_eco30324, w_eco30325, w_eco30326, w_eco30327, w_eco30328, w_eco30329, w_eco30330, w_eco30331, w_eco30332, w_eco30333, w_eco30334, w_eco30335, w_eco30336, w_eco30337, w_eco30338, w_eco30339, w_eco30340, w_eco30341, w_eco30342, w_eco30343, w_eco30344, w_eco30345, w_eco30346, w_eco30347, w_eco30348, w_eco30349, w_eco30350, w_eco30351, w_eco30352, w_eco30353, w_eco30354, w_eco30355, w_eco30356, w_eco30357, w_eco30358, w_eco30359, w_eco30360, w_eco30361, w_eco30362, w_eco30363, w_eco30364, w_eco30365, w_eco30366, w_eco30367, w_eco30368, w_eco30369, w_eco30370, w_eco30371, w_eco30372, w_eco30373, w_eco30374, w_eco30375, w_eco30376, w_eco30377, w_eco30378, w_eco30379, w_eco30380, w_eco30381, w_eco30382, w_eco30383, w_eco30384, w_eco30385, w_eco30386, w_eco30387, w_eco30388, w_eco30389, w_eco30390, w_eco30391, w_eco30392, w_eco30393, w_eco30394, w_eco30395, w_eco30396, w_eco30397, w_eco30398, w_eco30399, w_eco30400, w_eco30401, w_eco30402, w_eco30403, w_eco30404, w_eco30405, w_eco30406, w_eco30407, w_eco30408, w_eco30409, w_eco30410, w_eco30411, w_eco30412, w_eco30413, w_eco30414, w_eco30415, w_eco30416, w_eco30417, w_eco30418, w_eco30419, w_eco30420, w_eco30421, w_eco30422, w_eco30423, w_eco30424, w_eco30425, w_eco30426, w_eco30427, w_eco30428, w_eco30429, w_eco30430, w_eco30431, w_eco30432, w_eco30433, w_eco30434, w_eco30435, w_eco30436, w_eco30437, w_eco30438, w_eco30439, w_eco30440, w_eco30441, w_eco30442, w_eco30443, w_eco30444, w_eco30445, w_eco30446, w_eco30447, w_eco30448, w_eco30449, w_eco30450, w_eco30451, w_eco30452, w_eco30453, w_eco30454, w_eco30455, w_eco30456, w_eco30457, w_eco30458, w_eco30459, w_eco30460, w_eco30461, w_eco30462, w_eco30463, w_eco30464, w_eco30465, w_eco30466, w_eco30467, w_eco30468, w_eco30469, w_eco30470, w_eco30471, w_eco30472, w_eco30473, w_eco30474, w_eco30475, w_eco30476, w_eco30477, w_eco30478, w_eco30479, w_eco30480, w_eco30481, w_eco30482, w_eco30483, w_eco30484, w_eco30485, w_eco30486, w_eco30487, w_eco30488, w_eco30489, w_eco30490, w_eco30491, w_eco30492, w_eco30493, w_eco30494, w_eco30495, w_eco30496, w_eco30497, w_eco30498, w_eco30499, w_eco30500, w_eco30501, w_eco30502, w_eco30503, w_eco30504, w_eco30505, w_eco30506, w_eco30507, w_eco30508, w_eco30509, w_eco30510, w_eco30511, w_eco30512, w_eco30513, w_eco30514, w_eco30515, w_eco30516, w_eco30517, w_eco30518, w_eco30519, w_eco30520, w_eco30521, w_eco30522, w_eco30523, w_eco30524, w_eco30525, w_eco30526, w_eco30527, w_eco30528, w_eco30529, w_eco30530, w_eco30531, w_eco30532, w_eco30533, w_eco30534, w_eco30535, w_eco30536, w_eco30537, w_eco30538, w_eco30539, w_eco30540, w_eco30541, w_eco30542, w_eco30543, w_eco30544, w_eco30545, w_eco30546, w_eco30547, w_eco30548, w_eco30549, w_eco30550, w_eco30551, w_eco30552, w_eco30553, w_eco30554, w_eco30555, w_eco30556, w_eco30557, w_eco30558, w_eco30559, w_eco30560, w_eco30561, w_eco30562, w_eco30563, w_eco30564, w_eco30565, w_eco30566, w_eco30567, w_eco30568, w_eco30569, w_eco30570, w_eco30571, w_eco30572, w_eco30573, w_eco30574, w_eco30575, w_eco30576, w_eco30577, w_eco30578, w_eco30579, w_eco30580, w_eco30581, w_eco30582, w_eco30583, w_eco30584, w_eco30585, w_eco30586, w_eco30587, w_eco30588, w_eco30589, w_eco30590, w_eco30591, w_eco30592, w_eco30593, w_eco30594, w_eco30595, w_eco30596, w_eco30597, w_eco30598, w_eco30599, w_eco30600, w_eco30601, w_eco30602, w_eco30603, w_eco30604, w_eco30605, w_eco30606, w_eco30607, w_eco30608, w_eco30609, w_eco30610, w_eco30611, w_eco30612, w_eco30613, w_eco30614, w_eco30615, w_eco30616, w_eco30617, w_eco30618, w_eco30619, w_eco30620, w_eco30621, w_eco30622, w_eco30623, w_eco30624, w_eco30625, w_eco30626, w_eco30627, w_eco30628, w_eco30629, w_eco30630, w_eco30631, w_eco30632, w_eco30633, w_eco30634, w_eco30635, w_eco30636, w_eco30637, w_eco30638, w_eco30639, w_eco30640, w_eco30641, w_eco30642, w_eco30643, w_eco30644, w_eco30645, w_eco30646, w_eco30647, w_eco30648, w_eco30649, w_eco30650, w_eco30651, w_eco30652, w_eco30653, w_eco30654, w_eco30655, w_eco30656, w_eco30657, w_eco30658, w_eco30659, w_eco30660, w_eco30661, w_eco30662, w_eco30663, w_eco30664, w_eco30665, w_eco30666, w_eco30667, w_eco30668, w_eco30669, w_eco30670, w_eco30671, w_eco30672, w_eco30673, w_eco30674, w_eco30675, w_eco30676, w_eco30677, w_eco30678, w_eco30679, w_eco30680, w_eco30681, w_eco30682, w_eco30683, w_eco30684, w_eco30685, w_eco30686, w_eco30687, w_eco30688, w_eco30689, w_eco30690, w_eco30691, w_eco30692, w_eco30693, w_eco30694, w_eco30695, w_eco30696, w_eco30697, w_eco30698, w_eco30699, w_eco30700, w_eco30701, w_eco30702, w_eco30703, w_eco30704, w_eco30705, w_eco30706, w_eco30707, w_eco30708, w_eco30709, w_eco30710, w_eco30711, w_eco30712, w_eco30713, w_eco30714, w_eco30715, w_eco30716, w_eco30717, w_eco30718, w_eco30719, w_eco30720, w_eco30721, w_eco30722, w_eco30723, w_eco30724, w_eco30725, w_eco30726, w_eco30727, w_eco30728, w_eco30729, w_eco30730, w_eco30731, w_eco30732, w_eco30733, w_eco30734, w_eco30735, w_eco30736, w_eco30737, w_eco30738, w_eco30739, w_eco30740, w_eco30741, w_eco30742, w_eco30743, w_eco30744, w_eco30745, w_eco30746, w_eco30747, w_eco30748, w_eco30749, w_eco30750, w_eco30751, w_eco30752, w_eco30753, w_eco30754, w_eco30755, w_eco30756, w_eco30757, w_eco30758, w_eco30759, w_eco30760, w_eco30761, w_eco30762, w_eco30763, w_eco30764, w_eco30765, w_eco30766, w_eco30767, w_eco30768, w_eco30769, w_eco30770, w_eco30771, w_eco30772, w_eco30773, w_eco30774, w_eco30775, w_eco30776, w_eco30777, w_eco30778, w_eco30779, w_eco30780, w_eco30781, w_eco30782, w_eco30783, w_eco30784, w_eco30785, w_eco30786, w_eco30787, w_eco30788, w_eco30789, w_eco30790, w_eco30791, w_eco30792, w_eco30793, w_eco30794, w_eco30795, w_eco30796, w_eco30797, w_eco30798, w_eco30799, w_eco30800, w_eco30801, w_eco30802, w_eco30803, w_eco30804, w_eco30805, w_eco30806, w_eco30807, w_eco30808, w_eco30809, w_eco30810, w_eco30811, w_eco30812, w_eco30813, w_eco30814, w_eco30815, w_eco30816, w_eco30817, w_eco30818, w_eco30819, w_eco30820, w_eco30821, w_eco30822, w_eco30823, w_eco30824, w_eco30825, w_eco30826, w_eco30827, w_eco30828, w_eco30829, w_eco30830, w_eco30831, w_eco30832, w_eco30833, w_eco30834, w_eco30835, w_eco30836, w_eco30837, w_eco30838, w_eco30839, w_eco30840, w_eco30841, w_eco30842, w_eco30843, w_eco30844, w_eco30845, w_eco30846, w_eco30847, w_eco30848, w_eco30849, w_eco30850, w_eco30851, w_eco30852, w_eco30853, w_eco30854, w_eco30855, w_eco30856, w_eco30857, w_eco30858, w_eco30859, w_eco30860, w_eco30861, w_eco30862, w_eco30863, w_eco30864, w_eco30865, w_eco30866, w_eco30867, w_eco30868, w_eco30869, w_eco30870, w_eco30871, w_eco30872, w_eco30873, w_eco30874, w_eco30875, w_eco30876, w_eco30877, w_eco30878, w_eco30879, w_eco30880, w_eco30881, w_eco30882, w_eco30883, w_eco30884, w_eco30885, w_eco30886, w_eco30887, w_eco30888, w_eco30889, w_eco30890, w_eco30891, w_eco30892, w_eco30893, w_eco30894, w_eco30895, w_eco30896, w_eco30897, w_eco30898, w_eco30899, w_eco30900, w_eco30901, w_eco30902, w_eco30903, w_eco30904, w_eco30905, w_eco30906, w_eco30907, w_eco30908, w_eco30909, w_eco30910, w_eco30911, w_eco30912, w_eco30913, w_eco30914, w_eco30915, w_eco30916, w_eco30917, w_eco30918, w_eco30919, w_eco30920, w_eco30921, w_eco30922, w_eco30923, w_eco30924, w_eco30925, w_eco30926, w_eco30927, w_eco30928, w_eco30929, w_eco30930, w_eco30931, w_eco30932, w_eco30933, w_eco30934, w_eco30935, w_eco30936, w_eco30937, w_eco30938, w_eco30939, w_eco30940, w_eco30941, w_eco30942, w_eco30943, w_eco30944, w_eco30945, w_eco30946, w_eco30947, w_eco30948, w_eco30949, w_eco30950, w_eco30951, w_eco30952, w_eco30953, w_eco30954, w_eco30955, w_eco30956, w_eco30957, w_eco30958, w_eco30959, w_eco30960, w_eco30961, w_eco30962, w_eco30963, w_eco30964, w_eco30965, w_eco30966, w_eco30967, w_eco30968, w_eco30969, w_eco30970, w_eco30971, w_eco30972, w_eco30973, w_eco30974, w_eco30975, w_eco30976, w_eco30977, w_eco30978, w_eco30979, w_eco30980, w_eco30981, w_eco30982, w_eco30983, w_eco30984, w_eco30985, w_eco30986, w_eco30987, w_eco30988, w_eco30989, w_eco30990, w_eco30991, w_eco30992, w_eco30993, w_eco30994, w_eco30995, w_eco30996, w_eco30997, w_eco30998, w_eco30999, w_eco31000, w_eco31001, w_eco31002, w_eco31003, w_eco31004, w_eco31005, w_eco31006, w_eco31007, w_eco31008, w_eco31009, w_eco31010, w_eco31011, w_eco31012, w_eco31013, w_eco31014, w_eco31015, w_eco31016, w_eco31017, w_eco31018, w_eco31019, w_eco31020, w_eco31021, w_eco31022, w_eco31023, w_eco31024, w_eco31025, w_eco31026, w_eco31027, w_eco31028, w_eco31029, w_eco31030, w_eco31031, w_eco31032, w_eco31033, w_eco31034, w_eco31035, w_eco31036, w_eco31037, w_eco31038, w_eco31039, w_eco31040, w_eco31041, w_eco31042, w_eco31043, w_eco31044, w_eco31045, w_eco31046, w_eco31047, w_eco31048, w_eco31049, w_eco31050, w_eco31051, w_eco31052, w_eco31053, w_eco31054, w_eco31055, w_eco31056, w_eco31057, w_eco31058, w_eco31059, w_eco31060, w_eco31061, w_eco31062, w_eco31063, w_eco31064, w_eco31065, w_eco31066, w_eco31067, w_eco31068, w_eco31069, w_eco31070, w_eco31071, w_eco31072, w_eco31073, w_eco31074, w_eco31075, w_eco31076, w_eco31077, w_eco31078, w_eco31079, w_eco31080, w_eco31081, w_eco31082, w_eco31083, w_eco31084, w_eco31085, w_eco31086, w_eco31087, w_eco31088, w_eco31089, w_eco31090, w_eco31091, w_eco31092, w_eco31093, w_eco31094, w_eco31095, w_eco31096, w_eco31097, w_eco31098, w_eco31099, w_eco31100, w_eco31101, w_eco31102, w_eco31103, w_eco31104, w_eco31105, w_eco31106, w_eco31107, w_eco31108, w_eco31109, w_eco31110, w_eco31111, w_eco31112, w_eco31113, w_eco31114, w_eco31115, w_eco31116, w_eco31117, w_eco31118, w_eco31119, w_eco31120, w_eco31121, w_eco31122, w_eco31123, w_eco31124, w_eco31125, w_eco31126, w_eco31127, w_eco31128, w_eco31129, w_eco31130, w_eco31131, w_eco31132, w_eco31133, w_eco31134, w_eco31135, w_eco31136, w_eco31137, w_eco31138, w_eco31139, w_eco31140, w_eco31141, w_eco31142, w_eco31143, w_eco31144, w_eco31145, w_eco31146, w_eco31147, w_eco31148, w_eco31149, w_eco31150, w_eco31151, w_eco31152, w_eco31153, w_eco31154, w_eco31155, w_eco31156, w_eco31157, w_eco31158, w_eco31159, w_eco31160, w_eco31161, w_eco31162, w_eco31163, w_eco31164, w_eco31165, w_eco31166, w_eco31167, w_eco31168, w_eco31169, w_eco31170, w_eco31171, w_eco31172, w_eco31173, w_eco31174, w_eco31175, w_eco31176, w_eco31177, w_eco31178, w_eco31179, w_eco31180, w_eco31181, w_eco31182, w_eco31183, w_eco31184, w_eco31185, w_eco31186, w_eco31187, w_eco31188, w_eco31189, w_eco31190, w_eco31191, w_eco31192, w_eco31193, w_eco31194, w_eco31195, w_eco31196, w_eco31197, w_eco31198, w_eco31199, w_eco31200, w_eco31201, w_eco31202, w_eco31203, w_eco31204, w_eco31205, w_eco31206, w_eco31207, w_eco31208, w_eco31209, w_eco31210, w_eco31211, w_eco31212, w_eco31213, w_eco31214, w_eco31215, w_eco31216, w_eco31217, w_eco31218, w_eco31219, w_eco31220, w_eco31221, w_eco31222, w_eco31223, w_eco31224, w_eco31225, w_eco31226, w_eco31227, w_eco31228, w_eco31229, w_eco31230, w_eco31231, w_eco31232, w_eco31233, w_eco31234, w_eco31235, w_eco31236, w_eco31237, w_eco31238, w_eco31239, w_eco31240, w_eco31241, w_eco31242, w_eco31243, w_eco31244, w_eco31245, w_eco31246, w_eco31247, w_eco31248, w_eco31249, w_eco31250, w_eco31251, w_eco31252, w_eco31253, w_eco31254, w_eco31255, w_eco31256, w_eco31257, w_eco31258, w_eco31259, w_eco31260, w_eco31261, w_eco31262, w_eco31263, w_eco31264, w_eco31265, w_eco31266, w_eco31267, w_eco31268, w_eco31269, w_eco31270, w_eco31271, w_eco31272, w_eco31273, w_eco31274, w_eco31275, w_eco31276, w_eco31277, w_eco31278, w_eco31279, w_eco31280, w_eco31281, w_eco31282, w_eco31283, w_eco31284, w_eco31285, w_eco31286, w_eco31287, w_eco31288, w_eco31289, w_eco31290, w_eco31291, w_eco31292, w_eco31293, w_eco31294, w_eco31295, w_eco31296, w_eco31297, w_eco31298, w_eco31299, w_eco31300, w_eco31301, w_eco31302, w_eco31303, w_eco31304, w_eco31305, w_eco31306, w_eco31307, w_eco31308, w_eco31309, w_eco31310, w_eco31311, w_eco31312, w_eco31313, w_eco31314, w_eco31315, w_eco31316, w_eco31317, w_eco31318, w_eco31319, w_eco31320, w_eco31321, w_eco31322, w_eco31323, w_eco31324, w_eco31325, w_eco31326, w_eco31327, w_eco31328, w_eco31329, w_eco31330, w_eco31331, w_eco31332, w_eco31333, w_eco31334, w_eco31335, w_eco31336, w_eco31337, w_eco31338, w_eco31339, w_eco31340, w_eco31341, w_eco31342, w_eco31343, w_eco31344, w_eco31345, w_eco31346, w_eco31347, w_eco31348, w_eco31349, w_eco31350, w_eco31351, w_eco31352, w_eco31353, w_eco31354, w_eco31355, w_eco31356, w_eco31357, w_eco31358, w_eco31359, w_eco31360, w_eco31361, w_eco31362, w_eco31363, w_eco31364, w_eco31365, w_eco31366, w_eco31367, w_eco31368, w_eco31369, w_eco31370, w_eco31371, w_eco31372, w_eco31373, w_eco31374, w_eco31375, w_eco31376, w_eco31377, w_eco31378, w_eco31379, w_eco31380, w_eco31381, w_eco31382, w_eco31383, w_eco31384, w_eco31385, w_eco31386, w_eco31387, w_eco31388, w_eco31389, w_eco31390, w_eco31391, w_eco31392, w_eco31393, w_eco31394, w_eco31395, w_eco31396, w_eco31397, w_eco31398, w_eco31399, w_eco31400, w_eco31401, w_eco31402, w_eco31403, w_eco31404, w_eco31405, w_eco31406, w_eco31407, w_eco31408, w_eco31409, w_eco31410, w_eco31411, w_eco31412, w_eco31413, w_eco31414, w_eco31415, w_eco31416, w_eco31417, w_eco31418, w_eco31419, w_eco31420, w_eco31421, w_eco31422, w_eco31423, w_eco31424, w_eco31425, w_eco31426, w_eco31427, w_eco31428, w_eco31429, w_eco31430, w_eco31431, w_eco31432, w_eco31433, w_eco31434, w_eco31435, w_eco31436, w_eco31437, w_eco31438, w_eco31439, w_eco31440, w_eco31441, w_eco31442, w_eco31443, w_eco31444, w_eco31445, w_eco31446, w_eco31447, w_eco31448, w_eco31449, w_eco31450, w_eco31451, w_eco31452, w_eco31453, w_eco31454, w_eco31455, w_eco31456, w_eco31457, w_eco31458, w_eco31459, w_eco31460, w_eco31461, w_eco31462, w_eco31463, w_eco31464, w_eco31465, w_eco31466, w_eco31467, w_eco31468, w_eco31469, w_eco31470, w_eco31471, w_eco31472, w_eco31473, w_eco31474, w_eco31475, w_eco31476, w_eco31477, w_eco31478, w_eco31479, w_eco31480, w_eco31481, w_eco31482, w_eco31483, w_eco31484, w_eco31485, w_eco31486, w_eco31487, w_eco31488, w_eco31489, w_eco31490, w_eco31491, w_eco31492, w_eco31493, w_eco31494, w_eco31495, w_eco31496, w_eco31497, w_eco31498, w_eco31499, w_eco31500, w_eco31501, w_eco31502, w_eco31503, w_eco31504, w_eco31505, w_eco31506, w_eco31507, w_eco31508, w_eco31509, w_eco31510, w_eco31511, w_eco31512, w_eco31513, w_eco31514, w_eco31515, w_eco31516, w_eco31517, w_eco31518, w_eco31519, w_eco31520, w_eco31521, w_eco31522, w_eco31523, w_eco31524, w_eco31525, w_eco31526, w_eco31527, w_eco31528, w_eco31529, w_eco31530, w_eco31531, w_eco31532, w_eco31533, w_eco31534, w_eco31535, w_eco31536, w_eco31537, w_eco31538, w_eco31539, w_eco31540, w_eco31541, w_eco31542, w_eco31543, w_eco31544, w_eco31545, w_eco31546, w_eco31547, w_eco31548, w_eco31549, w_eco31550, w_eco31551, w_eco31552, w_eco31553, w_eco31554, w_eco31555, w_eco31556, w_eco31557, w_eco31558, w_eco31559, w_eco31560, w_eco31561, w_eco31562, w_eco31563, w_eco31564, w_eco31565, w_eco31566, w_eco31567, w_eco31568, w_eco31569, w_eco31570, w_eco31571, w_eco31572, w_eco31573, w_eco31574, w_eco31575, w_eco31576, w_eco31577, w_eco31578, w_eco31579, w_eco31580, w_eco31581, w_eco31582, w_eco31583, w_eco31584, w_eco31585, w_eco31586, w_eco31587, w_eco31588, w_eco31589, w_eco31590, w_eco31591, w_eco31592, w_eco31593, w_eco31594, w_eco31595, w_eco31596, w_eco31597, w_eco31598, w_eco31599, w_eco31600, w_eco31601, w_eco31602, w_eco31603, w_eco31604, w_eco31605, w_eco31606, w_eco31607, w_eco31608, w_eco31609, w_eco31610, w_eco31611, w_eco31612, w_eco31613, w_eco31614, w_eco31615, w_eco31616, w_eco31617, w_eco31618, w_eco31619, w_eco31620, w_eco31621, w_eco31622, w_eco31623, w_eco31624, w_eco31625, w_eco31626, w_eco31627, w_eco31628, w_eco31629, w_eco31630, w_eco31631, w_eco31632, w_eco31633, w_eco31634, w_eco31635, w_eco31636, w_eco31637, w_eco31638, w_eco31639, w_eco31640, w_eco31641, w_eco31642, w_eco31643, w_eco31644, w_eco31645, w_eco31646, w_eco31647, w_eco31648, w_eco31649, w_eco31650, w_eco31651, w_eco31652, w_eco31653, w_eco31654, w_eco31655, w_eco31656, w_eco31657, w_eco31658, w_eco31659, w_eco31660, w_eco31661, w_eco31662, w_eco31663, w_eco31664, w_eco31665, w_eco31666, w_eco31667, w_eco31668, w_eco31669, w_eco31670, w_eco31671, w_eco31672, w_eco31673, w_eco31674, w_eco31675, w_eco31676, w_eco31677, w_eco31678, w_eco31679, w_eco31680, w_eco31681, w_eco31682, w_eco31683, w_eco31684, w_eco31685, w_eco31686, w_eco31687, w_eco31688, w_eco31689, w_eco31690, w_eco31691, w_eco31692, w_eco31693, w_eco31694, w_eco31695, w_eco31696, w_eco31697, w_eco31698, w_eco31699, w_eco31700, w_eco31701, w_eco31702, w_eco31703, w_eco31704, w_eco31705, w_eco31706, w_eco31707, w_eco31708, w_eco31709, w_eco31710, w_eco31711, w_eco31712, w_eco31713, w_eco31714, w_eco31715, w_eco31716, w_eco31717, w_eco31718, w_eco31719, w_eco31720, w_eco31721, w_eco31722, w_eco31723, w_eco31724, w_eco31725, w_eco31726, w_eco31727, w_eco31728, w_eco31729, w_eco31730, w_eco31731, w_eco31732, w_eco31733, w_eco31734, w_eco31735, w_eco31736, w_eco31737, w_eco31738, w_eco31739, w_eco31740, w_eco31741, w_eco31742, w_eco31743, w_eco31744, w_eco31745, w_eco31746, w_eco31747, w_eco31748, w_eco31749, w_eco31750, w_eco31751, w_eco31752, w_eco31753, w_eco31754, w_eco31755, w_eco31756, w_eco31757, w_eco31758, w_eco31759, w_eco31760, w_eco31761, w_eco31762, w_eco31763, w_eco31764, w_eco31765, w_eco31766, w_eco31767, w_eco31768, w_eco31769, w_eco31770, w_eco31771, w_eco31772, w_eco31773, w_eco31774, w_eco31775, w_eco31776, w_eco31777, w_eco31778, w_eco31779, w_eco31780, w_eco31781, w_eco31782, w_eco31783, w_eco31784, w_eco31785, w_eco31786, w_eco31787, w_eco31788, w_eco31789, w_eco31790, w_eco31791, w_eco31792, w_eco31793, w_eco31794, w_eco31795, w_eco31796, w_eco31797, w_eco31798, w_eco31799, w_eco31800, w_eco31801, w_eco31802, w_eco31803, w_eco31804, w_eco31805, w_eco31806, w_eco31807, w_eco31808, w_eco31809, w_eco31810, w_eco31811, w_eco31812, w_eco31813, w_eco31814, w_eco31815, w_eco31816, w_eco31817, w_eco31818, w_eco31819, w_eco31820, w_eco31821, w_eco31822, w_eco31823, w_eco31824, w_eco31825, w_eco31826, w_eco31827, w_eco31828, w_eco31829, w_eco31830, w_eco31831, w_eco31832, w_eco31833, w_eco31834, w_eco31835, w_eco31836, w_eco31837, w_eco31838, w_eco31839, w_eco31840, w_eco31841, w_eco31842, w_eco31843, w_eco31844, w_eco31845, w_eco31846, w_eco31847, w_eco31848, w_eco31849, w_eco31850, w_eco31851, w_eco31852, w_eco31853, w_eco31854, w_eco31855, w_eco31856, w_eco31857, w_eco31858, w_eco31859, w_eco31860, w_eco31861, w_eco31862, w_eco31863, w_eco31864, w_eco31865, w_eco31866, w_eco31867, w_eco31868, w_eco31869, w_eco31870, w_eco31871, w_eco31872, w_eco31873, w_eco31874, w_eco31875, w_eco31876, w_eco31877, w_eco31878, w_eco31879, w_eco31880, w_eco31881, w_eco31882, w_eco31883, w_eco31884, w_eco31885, w_eco31886, w_eco31887, w_eco31888, w_eco31889, w_eco31890, w_eco31891, w_eco31892, w_eco31893, w_eco31894, w_eco31895, w_eco31896, w_eco31897, w_eco31898, w_eco31899, w_eco31900, w_eco31901, w_eco31902, w_eco31903, w_eco31904, w_eco31905, w_eco31906, w_eco31907, w_eco31908, w_eco31909, w_eco31910, w_eco31911, w_eco31912, w_eco31913, w_eco31914, w_eco31915, w_eco31916, w_eco31917, w_eco31918, w_eco31919, w_eco31920, w_eco31921, w_eco31922, w_eco31923, w_eco31924, w_eco31925, w_eco31926, w_eco31927, w_eco31928, w_eco31929, w_eco31930, w_eco31931, w_eco31932, w_eco31933, w_eco31934, w_eco31935, w_eco31936, w_eco31937, w_eco31938, w_eco31939, w_eco31940, w_eco31941, w_eco31942, w_eco31943, w_eco31944, w_eco31945, w_eco31946, w_eco31947, w_eco31948, w_eco31949, w_eco31950, w_eco31951, w_eco31952, w_eco31953, w_eco31954, w_eco31955, w_eco31956, w_eco31957, w_eco31958, w_eco31959, w_eco31960, w_eco31961, w_eco31962, w_eco31963, w_eco31964, w_eco31965, w_eco31966, w_eco31967, w_eco31968, w_eco31969, w_eco31970, w_eco31971, w_eco31972, w_eco31973, w_eco31974, w_eco31975, w_eco31976, w_eco31977, w_eco31978, w_eco31979, w_eco31980, w_eco31981, w_eco31982, w_eco31983, w_eco31984, w_eco31985, w_eco31986, w_eco31987, w_eco31988, w_eco31989, w_eco31990, w_eco31991, w_eco31992, w_eco31993, w_eco31994, w_eco31995, w_eco31996, w_eco31997, w_eco31998, w_eco31999, w_eco32000, w_eco32001, w_eco32002, w_eco32003, w_eco32004, w_eco32005, w_eco32006, w_eco32007, w_eco32008, w_eco32009, w_eco32010, w_eco32011, w_eco32012, w_eco32013, w_eco32014, w_eco32015, w_eco32016, w_eco32017, w_eco32018, w_eco32019, w_eco32020, w_eco32021, w_eco32022, w_eco32023, w_eco32024, w_eco32025, w_eco32026, w_eco32027, w_eco32028, w_eco32029, w_eco32030, w_eco32031, w_eco32032, w_eco32033, w_eco32034, w_eco32035, w_eco32036, w_eco32037, w_eco32038, w_eco32039, w_eco32040, w_eco32041, w_eco32042, w_eco32043, w_eco32044, w_eco32045, w_eco32046, w_eco32047, w_eco32048, w_eco32049, w_eco32050, w_eco32051, w_eco32052, w_eco32053, w_eco32054, w_eco32055, w_eco32056, w_eco32057, w_eco32058, w_eco32059, w_eco32060, w_eco32061, w_eco32062, w_eco32063, w_eco32064, w_eco32065, w_eco32066, w_eco32067, w_eco32068, w_eco32069, w_eco32070, w_eco32071, w_eco32072, w_eco32073, w_eco32074, w_eco32075, w_eco32076, w_eco32077, w_eco32078, w_eco32079, w_eco32080, w_eco32081, w_eco32082, w_eco32083, w_eco32084, w_eco32085, w_eco32086, w_eco32087, w_eco32088, w_eco32089, w_eco32090, w_eco32091, w_eco32092, w_eco32093, w_eco32094, w_eco32095, w_eco32096, w_eco32097, w_eco32098, w_eco32099, w_eco32100, w_eco32101, w_eco32102, w_eco32103, w_eco32104, w_eco32105, w_eco32106, w_eco32107, w_eco32108, w_eco32109, w_eco32110, w_eco32111, w_eco32112, w_eco32113, w_eco32114, w_eco32115, w_eco32116, w_eco32117, w_eco32118, w_eco32119, w_eco32120, w_eco32121, w_eco32122, w_eco32123, w_eco32124, w_eco32125, w_eco32126, w_eco32127, w_eco32128, w_eco32129, w_eco32130, w_eco32131, w_eco32132, w_eco32133, w_eco32134, w_eco32135, w_eco32136, w_eco32137, w_eco32138, w_eco32139, w_eco32140, w_eco32141, w_eco32142, w_eco32143, w_eco32144, w_eco32145, w_eco32146, w_eco32147, w_eco32148, w_eco32149, w_eco32150, w_eco32151, w_eco32152, w_eco32153, w_eco32154, w_eco32155, w_eco32156, w_eco32157, w_eco32158, w_eco32159, w_eco32160, w_eco32161, w_eco32162, w_eco32163, w_eco32164, w_eco32165, w_eco32166, w_eco32167, w_eco32168, w_eco32169, w_eco32170, w_eco32171, w_eco32172, w_eco32173, w_eco32174, w_eco32175, w_eco32176, w_eco32177, w_eco32178, w_eco32179, w_eco32180, w_eco32181, w_eco32182, w_eco32183, w_eco32184, w_eco32185, w_eco32186, w_eco32187, w_eco32188, w_eco32189, w_eco32190, w_eco32191, w_eco32192, w_eco32193, w_eco32194, w_eco32195, w_eco32196, w_eco32197, w_eco32198, w_eco32199, w_eco32200, w_eco32201, w_eco32202, w_eco32203, w_eco32204, w_eco32205, w_eco32206, w_eco32207, w_eco32208, w_eco32209, w_eco32210, w_eco32211, w_eco32212, w_eco32213, w_eco32214, w_eco32215, w_eco32216, w_eco32217, w_eco32218, w_eco32219, w_eco32220, w_eco32221, w_eco32222, w_eco32223, w_eco32224, w_eco32225, w_eco32226, w_eco32227, w_eco32228, w_eco32229, w_eco32230, w_eco32231, w_eco32232, w_eco32233, w_eco32234, w_eco32235, w_eco32236, w_eco32237, w_eco32238, w_eco32239, w_eco32240, w_eco32241, w_eco32242, w_eco32243, w_eco32244, w_eco32245, w_eco32246, w_eco32247, w_eco32248, w_eco32249, w_eco32250, w_eco32251, w_eco32252, w_eco32253, w_eco32254, w_eco32255, w_eco32256, w_eco32257, w_eco32258, w_eco32259, w_eco32260, w_eco32261, w_eco32262, w_eco32263, w_eco32264, w_eco32265, w_eco32266, w_eco32267, w_eco32268, w_eco32269, w_eco32270, w_eco32271, w_eco32272, w_eco32273, w_eco32274, w_eco32275, w_eco32276, w_eco32277, w_eco32278, w_eco32279, w_eco32280, w_eco32281, w_eco32282, w_eco32283, w_eco32284, w_eco32285, w_eco32286, w_eco32287, w_eco32288, w_eco32289, w_eco32290, w_eco32291, w_eco32292, w_eco32293, w_eco32294, w_eco32295, w_eco32296, w_eco32297, w_eco32298, w_eco32299, w_eco32300, w_eco32301, w_eco32302, w_eco32303, w_eco32304, w_eco32305, w_eco32306, w_eco32307, w_eco32308, w_eco32309, w_eco32310, w_eco32311, w_eco32312, w_eco32313, w_eco32314, w_eco32315, w_eco32316, w_eco32317, w_eco32318, w_eco32319, w_eco32320, w_eco32321, w_eco32322, w_eco32323, w_eco32324, w_eco32325, w_eco32326, w_eco32327, w_eco32328, w_eco32329, w_eco32330, w_eco32331, w_eco32332, w_eco32333, w_eco32334, w_eco32335, w_eco32336, w_eco32337, w_eco32338, w_eco32339, w_eco32340, w_eco32341, w_eco32342, w_eco32343, w_eco32344, w_eco32345, w_eco32346, w_eco32347, w_eco32348, w_eco32349, w_eco32350, w_eco32351, w_eco32352, w_eco32353, w_eco32354, w_eco32355, w_eco32356, w_eco32357, w_eco32358, w_eco32359, w_eco32360, w_eco32361, w_eco32362, w_eco32363, w_eco32364, w_eco32365, w_eco32366, w_eco32367, w_eco32368, w_eco32369, w_eco32370, w_eco32371, w_eco32372, w_eco32373, w_eco32374, w_eco32375, w_eco32376, w_eco32377, w_eco32378, w_eco32379, w_eco32380, w_eco32381, w_eco32382, w_eco32383, w_eco32384, w_eco32385, w_eco32386, w_eco32387, w_eco32388, w_eco32389, w_eco32390, w_eco32391, w_eco32392, w_eco32393, w_eco32394, w_eco32395, w_eco32396, w_eco32397, w_eco32398, w_eco32399, w_eco32400, w_eco32401, w_eco32402, w_eco32403, w_eco32404, w_eco32405, w_eco32406, w_eco32407, w_eco32408, w_eco32409, w_eco32410, w_eco32411, w_eco32412, w_eco32413, w_eco32414, w_eco32415, w_eco32416, w_eco32417, w_eco32418, w_eco32419, w_eco32420, w_eco32421, w_eco32422, w_eco32423, w_eco32424, w_eco32425, w_eco32426, w_eco32427, w_eco32428, w_eco32429, w_eco32430, w_eco32431, w_eco32432, w_eco32433, w_eco32434, w_eco32435, w_eco32436, w_eco32437, w_eco32438, w_eco32439, w_eco32440, w_eco32441, w_eco32442, w_eco32443, w_eco32444, w_eco32445, w_eco32446, w_eco32447, w_eco32448, w_eco32449, w_eco32450, w_eco32451, w_eco32452, w_eco32453, w_eco32454, w_eco32455, w_eco32456, w_eco32457, w_eco32458, w_eco32459, w_eco32460, w_eco32461, w_eco32462, w_eco32463, w_eco32464, w_eco32465, w_eco32466, w_eco32467, w_eco32468, w_eco32469, w_eco32470, w_eco32471, w_eco32472, w_eco32473, w_eco32474, w_eco32475, w_eco32476, w_eco32477, w_eco32478, w_eco32479, w_eco32480, w_eco32481, w_eco32482, w_eco32483, w_eco32484, w_eco32485, w_eco32486, w_eco32487, w_eco32488, w_eco32489, w_eco32490, w_eco32491, w_eco32492, w_eco32493, w_eco32494, w_eco32495, w_eco32496, w_eco32497, w_eco32498, w_eco32499, w_eco32500, w_eco32501, w_eco32502, w_eco32503, w_eco32504, w_eco32505, w_eco32506, w_eco32507, w_eco32508, w_eco32509, w_eco32510, w_eco32511, w_eco32512, w_eco32513, w_eco32514, w_eco32515, w_eco32516, w_eco32517, w_eco32518, w_eco32519, w_eco32520, w_eco32521, w_eco32522, w_eco32523, w_eco32524, w_eco32525, w_eco32526, w_eco32527, w_eco32528, w_eco32529, w_eco32530, w_eco32531, w_eco32532, w_eco32533, w_eco32534, w_eco32535, w_eco32536, w_eco32537, w_eco32538, w_eco32539, w_eco32540, w_eco32541, w_eco32542, w_eco32543, w_eco32544, w_eco32545, w_eco32546, w_eco32547, w_eco32548, w_eco32549, w_eco32550, w_eco32551, w_eco32552, w_eco32553, w_eco32554, w_eco32555, w_eco32556, w_eco32557, w_eco32558, w_eco32559, w_eco32560, w_eco32561, w_eco32562, w_eco32563, w_eco32564, w_eco32565, w_eco32566, w_eco32567, w_eco32568, w_eco32569, w_eco32570, w_eco32571, w_eco32572, w_eco32573, w_eco32574, w_eco32575, w_eco32576, w_eco32577, w_eco32578, w_eco32579, w_eco32580, w_eco32581, w_eco32582, w_eco32583, w_eco32584, w_eco32585, w_eco32586, w_eco32587, w_eco32588, w_eco32589, w_eco32590, w_eco32591, w_eco32592, w_eco32593, w_eco32594, w_eco32595, w_eco32596, w_eco32597, w_eco32598, w_eco32599, w_eco32600, w_eco32601, w_eco32602, w_eco32603, w_eco32604, w_eco32605, w_eco32606, w_eco32607, w_eco32608, w_eco32609, w_eco32610, w_eco32611, w_eco32612, w_eco32613, w_eco32614, w_eco32615, w_eco32616, w_eco32617, w_eco32618, w_eco32619, w_eco32620, w_eco32621, w_eco32622, w_eco32623, w_eco32624, w_eco32625, w_eco32626, w_eco32627, w_eco32628, w_eco32629, w_eco32630, w_eco32631, w_eco32632, w_eco32633, w_eco32634, w_eco32635, w_eco32636, w_eco32637, w_eco32638, w_eco32639, w_eco32640, w_eco32641, w_eco32642, w_eco32643, w_eco32644, w_eco32645, w_eco32646, w_eco32647, w_eco32648, w_eco32649, w_eco32650, w_eco32651, w_eco32652, w_eco32653, w_eco32654, w_eco32655, w_eco32656, w_eco32657, w_eco32658, w_eco32659, w_eco32660, w_eco32661, w_eco32662, w_eco32663, w_eco32664, w_eco32665, w_eco32666, w_eco32667, w_eco32668, w_eco32669, w_eco32670, w_eco32671, w_eco32672, w_eco32673, w_eco32674, w_eco32675, w_eco32676, w_eco32677, w_eco32678, w_eco32679, w_eco32680, w_eco32681, w_eco32682, w_eco32683, w_eco32684, w_eco32685, w_eco32686, w_eco32687, w_eco32688, w_eco32689, w_eco32690, w_eco32691, w_eco32692, w_eco32693, w_eco32694, w_eco32695, w_eco32696, w_eco32697, w_eco32698, w_eco32699, w_eco32700, w_eco32701, w_eco32702, w_eco32703, w_eco32704, w_eco32705, w_eco32706, w_eco32707, w_eco32708, w_eco32709, w_eco32710, w_eco32711, w_eco32712, w_eco32713, w_eco32714, w_eco32715, w_eco32716, w_eco32717, w_eco32718, w_eco32719, w_eco32720, w_eco32721, w_eco32722, w_eco32723, w_eco32724, w_eco32725, w_eco32726, w_eco32727, w_eco32728, w_eco32729, w_eco32730, w_eco32731, w_eco32732, w_eco32733, w_eco32734, w_eco32735, w_eco32736, w_eco32737, w_eco32738, w_eco32739, w_eco32740, w_eco32741, w_eco32742, w_eco32743, w_eco32744, w_eco32745, w_eco32746, w_eco32747, w_eco32748, w_eco32749, w_eco32750, w_eco32751, w_eco32752, w_eco32753, w_eco32754, w_eco32755, w_eco32756, w_eco32757, w_eco32758, w_eco32759, w_eco32760, w_eco32761, w_eco32762, w_eco32763, w_eco32764, w_eco32765, w_eco32766, w_eco32767, w_eco32768, w_eco32769, w_eco32770, w_eco32771, w_eco32772, w_eco32773, w_eco32774, w_eco32775, w_eco32776, w_eco32777, w_eco32778, w_eco32779, w_eco32780, w_eco32781, w_eco32782, w_eco32783, w_eco32784, w_eco32785, w_eco32786, w_eco32787, w_eco32788, w_eco32789, w_eco32790, w_eco32791, w_eco32792, w_eco32793, w_eco32794, w_eco32795, w_eco32796, w_eco32797, w_eco32798, w_eco32799, w_eco32800, w_eco32801, w_eco32802, w_eco32803, w_eco32804, w_eco32805, w_eco32806, w_eco32807, w_eco32808, w_eco32809, w_eco32810, w_eco32811, w_eco32812, w_eco32813, w_eco32814, w_eco32815, w_eco32816, w_eco32817, w_eco32818, w_eco32819, w_eco32820, w_eco32821, w_eco32822, w_eco32823, w_eco32824, w_eco32825, w_eco32826, w_eco32827, w_eco32828, w_eco32829, w_eco32830, w_eco32831, w_eco32832, w_eco32833, w_eco32834, w_eco32835, w_eco32836, w_eco32837, w_eco32838, w_eco32839, w_eco32840, w_eco32841, w_eco32842, w_eco32843, w_eco32844, w_eco32845, w_eco32846, w_eco32847, w_eco32848, w_eco32849, w_eco32850, w_eco32851, w_eco32852, w_eco32853, w_eco32854, w_eco32855, w_eco32856, w_eco32857, w_eco32858, w_eco32859, w_eco32860, w_eco32861, w_eco32862, w_eco32863, w_eco32864, w_eco32865, w_eco32866, w_eco32867, w_eco32868, w_eco32869, w_eco32870, w_eco32871, w_eco32872, w_eco32873, w_eco32874, w_eco32875, w_eco32876, w_eco32877, w_eco32878, w_eco32879, w_eco32880, w_eco32881, w_eco32882, w_eco32883, w_eco32884, w_eco32885, w_eco32886, w_eco32887, w_eco32888, w_eco32889, w_eco32890, w_eco32891, w_eco32892, w_eco32893, w_eco32894, w_eco32895, w_eco32896, w_eco32897, w_eco32898, w_eco32899, w_eco32900, w_eco32901, w_eco32902, w_eco32903, w_eco32904, w_eco32905, w_eco32906, w_eco32907, w_eco32908, w_eco32909, w_eco32910, w_eco32911, w_eco32912, w_eco32913, w_eco32914, w_eco32915, w_eco32916, w_eco32917, w_eco32918, w_eco32919, w_eco32920, w_eco32921, w_eco32922, w_eco32923, w_eco32924, w_eco32925, w_eco32926, w_eco32927, w_eco32928, w_eco32929, w_eco32930, w_eco32931, w_eco32932, w_eco32933, w_eco32934, w_eco32935, w_eco32936, w_eco32937, w_eco32938, w_eco32939, w_eco32940, w_eco32941, w_eco32942, w_eco32943, w_eco32944, w_eco32945, w_eco32946, w_eco32947, w_eco32948, w_eco32949, w_eco32950, w_eco32951, w_eco32952, w_eco32953, w_eco32954, w_eco32955, w_eco32956, w_eco32957, w_eco32958, w_eco32959, w_eco32960, w_eco32961, w_eco32962, w_eco32963, w_eco32964, w_eco32965, w_eco32966, w_eco32967, w_eco32968, w_eco32969, w_eco32970, w_eco32971, w_eco32972, w_eco32973, w_eco32974, w_eco32975, w_eco32976, w_eco32977, w_eco32978, w_eco32979, w_eco32980, w_eco32981, w_eco32982, w_eco32983, w_eco32984, w_eco32985, w_eco32986, w_eco32987, w_eco32988, w_eco32989, w_eco32990, w_eco32991, w_eco32992, w_eco32993, w_eco32994, w_eco32995, w_eco32996, w_eco32997, w_eco32998, w_eco32999, w_eco33000, w_eco33001, w_eco33002, w_eco33003, w_eco33004, w_eco33005, w_eco33006, w_eco33007, w_eco33008, w_eco33009, w_eco33010, w_eco33011, w_eco33012, w_eco33013, w_eco33014, w_eco33015, w_eco33016, w_eco33017, w_eco33018, w_eco33019, w_eco33020, w_eco33021, w_eco33022, w_eco33023, w_eco33024, w_eco33025, w_eco33026, w_eco33027, w_eco33028, w_eco33029, w_eco33030, w_eco33031, w_eco33032, w_eco33033, w_eco33034, w_eco33035, w_eco33036, w_eco33037, w_eco33038, w_eco33039, w_eco33040, w_eco33041, w_eco33042, w_eco33043, w_eco33044, w_eco33045, w_eco33046, w_eco33047, w_eco33048, w_eco33049, w_eco33050, w_eco33051, w_eco33052, w_eco33053, w_eco33054, w_eco33055, w_eco33056, w_eco33057, w_eco33058, w_eco33059, w_eco33060, w_eco33061, w_eco33062, w_eco33063, w_eco33064, w_eco33065, w_eco33066, w_eco33067, w_eco33068, w_eco33069, w_eco33070, w_eco33071, w_eco33072, w_eco33073, w_eco33074, w_eco33075, w_eco33076, w_eco33077, w_eco33078, w_eco33079, w_eco33080, w_eco33081, w_eco33082, w_eco33083, w_eco33084, w_eco33085, w_eco33086, w_eco33087, w_eco33088, w_eco33089, w_eco33090, w_eco33091, w_eco33092, w_eco33093, w_eco33094, w_eco33095, w_eco33096, w_eco33097, w_eco33098, w_eco33099, w_eco33100, w_eco33101, w_eco33102, w_eco33103, w_eco33104, w_eco33105, w_eco33106, w_eco33107, w_eco33108, w_eco33109, w_eco33110, w_eco33111, w_eco33112, w_eco33113, w_eco33114, w_eco33115, w_eco33116, w_eco33117, w_eco33118, w_eco33119, w_eco33120, w_eco33121, w_eco33122, w_eco33123, w_eco33124, w_eco33125, w_eco33126, w_eco33127, w_eco33128, w_eco33129, w_eco33130, w_eco33131, w_eco33132, w_eco33133, w_eco33134, w_eco33135, w_eco33136, w_eco33137, w_eco33138, w_eco33139, w_eco33140, w_eco33141, w_eco33142, w_eco33143, w_eco33144, w_eco33145, w_eco33146, w_eco33147, w_eco33148, w_eco33149, w_eco33150, w_eco33151, w_eco33152, w_eco33153, w_eco33154, w_eco33155, w_eco33156, w_eco33157, w_eco33158, w_eco33159, w_eco33160, w_eco33161, w_eco33162, w_eco33163, w_eco33164, w_eco33165, w_eco33166, w_eco33167, w_eco33168, w_eco33169, w_eco33170, w_eco33171, w_eco33172, w_eco33173, w_eco33174, w_eco33175, w_eco33176, w_eco33177, w_eco33178, w_eco33179, w_eco33180, w_eco33181, w_eco33182, w_eco33183, w_eco33184, w_eco33185, w_eco33186, w_eco33187, w_eco33188, w_eco33189, w_eco33190, w_eco33191, w_eco33192, w_eco33193, w_eco33194, w_eco33195, w_eco33196, w_eco33197, w_eco33198, w_eco33199, w_eco33200, w_eco33201, w_eco33202, w_eco33203, w_eco33204, w_eco33205, w_eco33206, w_eco33207, w_eco33208, w_eco33209, w_eco33210, w_eco33211, w_eco33212, w_eco33213, w_eco33214, w_eco33215, w_eco33216, w_eco33217, w_eco33218, w_eco33219, w_eco33220, w_eco33221, w_eco33222, w_eco33223, w_eco33224, w_eco33225, w_eco33226, w_eco33227, w_eco33228, w_eco33229, w_eco33230, w_eco33231, w_eco33232, w_eco33233, w_eco33234, w_eco33235, w_eco33236, w_eco33237, w_eco33238, w_eco33239, w_eco33240, w_eco33241, w_eco33242, w_eco33243, w_eco33244, w_eco33245, w_eco33246, w_eco33247, w_eco33248, w_eco33249, w_eco33250, w_eco33251, w_eco33252, w_eco33253, w_eco33254, w_eco33255, w_eco33256, w_eco33257, w_eco33258, w_eco33259, w_eco33260, w_eco33261, w_eco33262, w_eco33263, w_eco33264, w_eco33265, w_eco33266, w_eco33267, w_eco33268, w_eco33269, w_eco33270, w_eco33271, w_eco33272, w_eco33273, w_eco33274, w_eco33275, w_eco33276, w_eco33277, w_eco33278, w_eco33279, w_eco33280, w_eco33281, w_eco33282, w_eco33283, w_eco33284, w_eco33285, w_eco33286, w_eco33287, w_eco33288, w_eco33289, w_eco33290, w_eco33291, w_eco33292, w_eco33293, w_eco33294, w_eco33295, w_eco33296, w_eco33297, w_eco33298, w_eco33299, w_eco33300, w_eco33301, w_eco33302, w_eco33303, w_eco33304, w_eco33305, w_eco33306, w_eco33307, w_eco33308, w_eco33309, w_eco33310, w_eco33311, w_eco33312, w_eco33313, w_eco33314, w_eco33315, w_eco33316, w_eco33317, w_eco33318, w_eco33319, w_eco33320, w_eco33321, w_eco33322, w_eco33323, w_eco33324, w_eco33325, w_eco33326, w_eco33327, w_eco33328, w_eco33329, w_eco33330, w_eco33331, w_eco33332, w_eco33333, w_eco33334, w_eco33335, w_eco33336, w_eco33337, w_eco33338, w_eco33339, w_eco33340, w_eco33341, w_eco33342, w_eco33343, w_eco33344, w_eco33345, w_eco33346, w_eco33347, w_eco33348, w_eco33349, w_eco33350, w_eco33351, w_eco33352, w_eco33353, w_eco33354, w_eco33355, w_eco33356, w_eco33357, w_eco33358, w_eco33359, w_eco33360, w_eco33361, w_eco33362, w_eco33363, w_eco33364, w_eco33365, w_eco33366, w_eco33367, w_eco33368, w_eco33369, w_eco33370, w_eco33371, w_eco33372, w_eco33373, w_eco33374, w_eco33375, w_eco33376, w_eco33377, w_eco33378, w_eco33379, w_eco33380, w_eco33381, w_eco33382, w_eco33383, w_eco33384, w_eco33385, w_eco33386, w_eco33387, w_eco33388, w_eco33389, w_eco33390, w_eco33391, w_eco33392, w_eco33393, w_eco33394, w_eco33395, w_eco33396, w_eco33397, w_eco33398, w_eco33399, w_eco33400, w_eco33401, w_eco33402, w_eco33403, w_eco33404, w_eco33405, w_eco33406, w_eco33407, w_eco33408, w_eco33409, w_eco33410, w_eco33411, w_eco33412, w_eco33413, w_eco33414, w_eco33415, w_eco33416, w_eco33417, w_eco33418, w_eco33419, w_eco33420, w_eco33421, w_eco33422, w_eco33423, w_eco33424, w_eco33425, w_eco33426, w_eco33427, w_eco33428, w_eco33429, w_eco33430, w_eco33431, w_eco33432, w_eco33433, w_eco33434, w_eco33435, w_eco33436, w_eco33437, w_eco33438, w_eco33439, w_eco33440, w_eco33441, w_eco33442, w_eco33443, w_eco33444, w_eco33445, w_eco33446, w_eco33447, w_eco33448, w_eco33449, w_eco33450, w_eco33451, w_eco33452, w_eco33453, w_eco33454, w_eco33455, w_eco33456, w_eco33457, w_eco33458, w_eco33459, w_eco33460, w_eco33461, w_eco33462, w_eco33463, w_eco33464, w_eco33465, w_eco33466, w_eco33467, w_eco33468, w_eco33469, w_eco33470, w_eco33471, w_eco33472, w_eco33473, w_eco33474, w_eco33475, w_eco33476, w_eco33477, w_eco33478, w_eco33479, w_eco33480, w_eco33481, w_eco33482, w_eco33483, w_eco33484, w_eco33485, w_eco33486, w_eco33487, w_eco33488, w_eco33489, w_eco33490, w_eco33491, w_eco33492, w_eco33493, w_eco33494, w_eco33495, w_eco33496, w_eco33497, w_eco33498, w_eco33499, w_eco33500, w_eco33501, w_eco33502, w_eco33503, w_eco33504, w_eco33505, w_eco33506, w_eco33507, w_eco33508, w_eco33509, w_eco33510, w_eco33511, w_eco33512, w_eco33513, w_eco33514, w_eco33515, w_eco33516, w_eco33517, w_eco33518, w_eco33519, w_eco33520, w_eco33521, w_eco33522, w_eco33523, w_eco33524, w_eco33525, w_eco33526, w_eco33527, w_eco33528, w_eco33529, w_eco33530, w_eco33531, w_eco33532, w_eco33533, w_eco33534, w_eco33535, w_eco33536, w_eco33537, w_eco33538, w_eco33539, w_eco33540, w_eco33541, w_eco33542, w_eco33543, w_eco33544, w_eco33545, w_eco33546, w_eco33547, w_eco33548, w_eco33549, w_eco33550, w_eco33551, w_eco33552, w_eco33553, w_eco33554, w_eco33555, w_eco33556, w_eco33557, w_eco33558, w_eco33559, w_eco33560, w_eco33561, w_eco33562, w_eco33563, w_eco33564, w_eco33565, w_eco33566, w_eco33567, w_eco33568, w_eco33569, w_eco33570, w_eco33571, w_eco33572, w_eco33573, w_eco33574, w_eco33575, w_eco33576, w_eco33577, w_eco33578, w_eco33579, w_eco33580, w_eco33581, w_eco33582, w_eco33583, w_eco33584, w_eco33585, w_eco33586, w_eco33587, w_eco33588, w_eco33589, w_eco33590, w_eco33591, w_eco33592, w_eco33593, w_eco33594, w_eco33595, w_eco33596, w_eco33597, w_eco33598, w_eco33599, w_eco33600, w_eco33601, w_eco33602, w_eco33603, w_eco33604, w_eco33605, w_eco33606, w_eco33607, w_eco33608, w_eco33609, w_eco33610, w_eco33611, w_eco33612, w_eco33613, w_eco33614, w_eco33615, w_eco33616, w_eco33617, w_eco33618, w_eco33619, w_eco33620, w_eco33621, w_eco33622, w_eco33623, w_eco33624, w_eco33625, w_eco33626, w_eco33627, w_eco33628, w_eco33629, w_eco33630, w_eco33631, w_eco33632, w_eco33633, w_eco33634, w_eco33635, w_eco33636, w_eco33637, w_eco33638, w_eco33639, w_eco33640, w_eco33641, w_eco33642, w_eco33643, w_eco33644, w_eco33645, w_eco33646, w_eco33647, w_eco33648, w_eco33649, w_eco33650, w_eco33651, w_eco33652, w_eco33653, w_eco33654, w_eco33655, w_eco33656, w_eco33657, w_eco33658, w_eco33659, w_eco33660, w_eco33661, w_eco33662, w_eco33663, w_eco33664, w_eco33665, w_eco33666, w_eco33667, w_eco33668, w_eco33669, w_eco33670, w_eco33671, w_eco33672, w_eco33673, w_eco33674, w_eco33675, w_eco33676, w_eco33677, w_eco33678, w_eco33679, w_eco33680, w_eco33681, w_eco33682, w_eco33683, w_eco33684, w_eco33685, w_eco33686, w_eco33687, w_eco33688, w_eco33689, w_eco33690, w_eco33691, w_eco33692, w_eco33693, w_eco33694, w_eco33695, w_eco33696, w_eco33697, w_eco33698, w_eco33699, w_eco33700, w_eco33701, w_eco33702, w_eco33703, w_eco33704, w_eco33705, w_eco33706, w_eco33707, w_eco33708, w_eco33709, w_eco33710, w_eco33711, w_eco33712, w_eco33713, w_eco33714, w_eco33715, w_eco33716, w_eco33717, w_eco33718, w_eco33719, w_eco33720, w_eco33721, w_eco33722, w_eco33723, w_eco33724, w_eco33725, w_eco33726, w_eco33727, w_eco33728, w_eco33729, w_eco33730, w_eco33731, w_eco33732, w_eco33733, w_eco33734, w_eco33735, w_eco33736, w_eco33737, w_eco33738, w_eco33739, w_eco33740, w_eco33741, w_eco33742, w_eco33743, w_eco33744, w_eco33745, w_eco33746, w_eco33747, w_eco33748, w_eco33749, w_eco33750, w_eco33751, w_eco33752, w_eco33753, w_eco33754, w_eco33755, w_eco33756, w_eco33757, w_eco33758, w_eco33759, w_eco33760, w_eco33761, w_eco33762, w_eco33763, w_eco33764, w_eco33765, w_eco33766, w_eco33767, w_eco33768, w_eco33769, w_eco33770, w_eco33771, w_eco33772, w_eco33773, w_eco33774, w_eco33775, w_eco33776, w_eco33777, w_eco33778, w_eco33779, w_eco33780, w_eco33781, w_eco33782, w_eco33783, w_eco33784, w_eco33785, w_eco33786, w_eco33787, w_eco33788, w_eco33789, w_eco33790, w_eco33791, w_eco33792, w_eco33793, w_eco33794, w_eco33795, w_eco33796, w_eco33797, w_eco33798, w_eco33799, w_eco33800, w_eco33801, w_eco33802, w_eco33803, w_eco33804, w_eco33805, w_eco33806, w_eco33807, w_eco33808, w_eco33809, w_eco33810, w_eco33811, w_eco33812, w_eco33813, w_eco33814, w_eco33815, w_eco33816, w_eco33817, w_eco33818, w_eco33819, w_eco33820, w_eco33821, w_eco33822, w_eco33823, w_eco33824, w_eco33825, w_eco33826, w_eco33827, w_eco33828, w_eco33829, w_eco33830, w_eco33831, w_eco33832, w_eco33833, w_eco33834, w_eco33835, w_eco33836, w_eco33837, w_eco33838, w_eco33839, w_eco33840, w_eco33841, w_eco33842, w_eco33843, w_eco33844, w_eco33845, w_eco33846, w_eco33847, w_eco33848, w_eco33849, w_eco33850, w_eco33851, w_eco33852, w_eco33853, w_eco33854, w_eco33855, w_eco33856, w_eco33857, w_eco33858, w_eco33859, w_eco33860, w_eco33861, w_eco33862, w_eco33863, w_eco33864, w_eco33865, w_eco33866, w_eco33867, w_eco33868, w_eco33869, w_eco33870, w_eco33871, w_eco33872, w_eco33873, w_eco33874, w_eco33875, w_eco33876, w_eco33877, w_eco33878, w_eco33879, w_eco33880, w_eco33881, w_eco33882, w_eco33883, w_eco33884, w_eco33885, w_eco33886, w_eco33887, w_eco33888, w_eco33889, w_eco33890, w_eco33891, w_eco33892, w_eco33893, w_eco33894, w_eco33895, w_eco33896, w_eco33897, w_eco33898, w_eco33899, w_eco33900, w_eco33901, w_eco33902, w_eco33903, w_eco33904, w_eco33905, w_eco33906, w_eco33907, w_eco33908, w_eco33909, w_eco33910, w_eco33911, w_eco33912, w_eco33913, w_eco33914, w_eco33915, w_eco33916, w_eco33917, w_eco33918, w_eco33919, w_eco33920, w_eco33921, w_eco33922, w_eco33923, w_eco33924, w_eco33925, w_eco33926, w_eco33927, w_eco33928, w_eco33929, w_eco33930, w_eco33931, w_eco33932, w_eco33933, w_eco33934, w_eco33935, w_eco33936, w_eco33937, w_eco33938, w_eco33939, w_eco33940, w_eco33941, w_eco33942, w_eco33943, w_eco33944, w_eco33945, w_eco33946, w_eco33947, w_eco33948, w_eco33949, w_eco33950, w_eco33951, w_eco33952, w_eco33953, w_eco33954, w_eco33955, w_eco33956, w_eco33957, w_eco33958, w_eco33959, w_eco33960, w_eco33961, w_eco33962, w_eco33963, w_eco33964, w_eco33965, w_eco33966, w_eco33967, w_eco33968, w_eco33969, w_eco33970, w_eco33971, w_eco33972, w_eco33973, w_eco33974, w_eco33975, w_eco33976, w_eco33977, w_eco33978, w_eco33979, w_eco33980, w_eco33981, w_eco33982, w_eco33983, w_eco33984, w_eco33985, w_eco33986, w_eco33987, w_eco33988, w_eco33989, w_eco33990, w_eco33991, w_eco33992, w_eco33993, w_eco33994, w_eco33995, w_eco33996, w_eco33997, w_eco33998, w_eco33999, w_eco34000, w_eco34001, w_eco34002, w_eco34003, w_eco34004, w_eco34005, w_eco34006, w_eco34007, w_eco34008, w_eco34009, w_eco34010, w_eco34011, w_eco34012, w_eco34013, w_eco34014, w_eco34015, w_eco34016, w_eco34017, w_eco34018, w_eco34019, w_eco34020, w_eco34021, w_eco34022, w_eco34023, w_eco34024, w_eco34025, w_eco34026, w_eco34027, w_eco34028, w_eco34029, w_eco34030, w_eco34031, w_eco34032, w_eco34033, w_eco34034, w_eco34035, w_eco34036, w_eco34037, w_eco34038, w_eco34039, w_eco34040, w_eco34041, w_eco34042, w_eco34043, w_eco34044, w_eco34045, w_eco34046, w_eco34047, w_eco34048, w_eco34049, w_eco34050, w_eco34051, w_eco34052, w_eco34053, w_eco34054, w_eco34055, w_eco34056, w_eco34057, w_eco34058, w_eco34059, w_eco34060, w_eco34061, w_eco34062, w_eco34063, w_eco34064, w_eco34065, w_eco34066, w_eco34067, w_eco34068, w_eco34069, w_eco34070, w_eco34071, w_eco34072, w_eco34073, w_eco34074, w_eco34075, w_eco34076, w_eco34077, w_eco34078, w_eco34079, w_eco34080, w_eco34081, w_eco34082, w_eco34083, w_eco34084, w_eco34085, w_eco34086, w_eco34087, w_eco34088, w_eco34089, w_eco34090, w_eco34091, w_eco34092, w_eco34093, w_eco34094, w_eco34095, w_eco34096, w_eco34097, w_eco34098, w_eco34099, w_eco34100, w_eco34101, w_eco34102, w_eco34103, w_eco34104, w_eco34105, w_eco34106, w_eco34107, w_eco34108, w_eco34109, w_eco34110, w_eco34111, w_eco34112, w_eco34113, w_eco34114, w_eco34115, w_eco34116, w_eco34117, w_eco34118, w_eco34119, w_eco34120, w_eco34121, w_eco34122, w_eco34123, w_eco34124, w_eco34125, w_eco34126, w_eco34127, w_eco34128, w_eco34129, w_eco34130, w_eco34131, w_eco34132, w_eco34133, w_eco34134, w_eco34135, w_eco34136, w_eco34137, w_eco34138, w_eco34139, w_eco34140, w_eco34141, w_eco34142, w_eco34143, w_eco34144, w_eco34145, w_eco34146, w_eco34147, w_eco34148, w_eco34149, w_eco34150, w_eco34151, w_eco34152, w_eco34153, w_eco34154, w_eco34155, w_eco34156, w_eco34157, w_eco34158, w_eco34159, w_eco34160, w_eco34161, w_eco34162, w_eco34163, w_eco34164, w_eco34165, w_eco34166, w_eco34167, w_eco34168, w_eco34169, w_eco34170, w_eco34171, w_eco34172, w_eco34173, w_eco34174, w_eco34175, w_eco34176, w_eco34177, w_eco34178, w_eco34179, w_eco34180, w_eco34181, w_eco34182, w_eco34183, w_eco34184, w_eco34185, w_eco34186, w_eco34187, w_eco34188, w_eco34189, w_eco34190, w_eco34191, w_eco34192, w_eco34193, w_eco34194, w_eco34195, w_eco34196, w_eco34197, w_eco34198, w_eco34199, w_eco34200, w_eco34201, w_eco34202, w_eco34203, w_eco34204, w_eco34205, w_eco34206, w_eco34207, w_eco34208, w_eco34209, w_eco34210, w_eco34211, w_eco34212, w_eco34213, w_eco34214, w_eco34215, w_eco34216, w_eco34217, w_eco34218, w_eco34219, w_eco34220, w_eco34221, w_eco34222, w_eco34223, w_eco34224, w_eco34225, w_eco34226, w_eco34227, w_eco34228, w_eco34229, w_eco34230, w_eco34231, w_eco34232, w_eco34233, w_eco34234, w_eco34235, w_eco34236, w_eco34237, w_eco34238, w_eco34239, w_eco34240, w_eco34241, w_eco34242, w_eco34243, w_eco34244, w_eco34245, w_eco34246, w_eco34247, w_eco34248, w_eco34249, w_eco34250, w_eco34251, w_eco34252, w_eco34253, w_eco34254, w_eco34255, w_eco34256, w_eco34257, w_eco34258, w_eco34259, w_eco34260, w_eco34261, w_eco34262, w_eco34263, w_eco34264, w_eco34265, w_eco34266, w_eco34267, w_eco34268, w_eco34269, w_eco34270, w_eco34271, w_eco34272, w_eco34273, w_eco34274, w_eco34275, w_eco34276, w_eco34277, w_eco34278, w_eco34279, w_eco34280, w_eco34281, w_eco34282, w_eco34283, w_eco34284, w_eco34285, w_eco34286, w_eco34287, w_eco34288, w_eco34289, w_eco34290, w_eco34291, w_eco34292, w_eco34293, w_eco34294, w_eco34295, w_eco34296, w_eco34297, w_eco34298, w_eco34299, w_eco34300, w_eco34301, w_eco34302, w_eco34303, w_eco34304, w_eco34305, w_eco34306, w_eco34307, w_eco34308, w_eco34309, w_eco34310, w_eco34311, w_eco34312, w_eco34313, w_eco34314, w_eco34315, w_eco34316, w_eco34317, w_eco34318, w_eco34319, w_eco34320, w_eco34321, w_eco34322, w_eco34323, w_eco34324, w_eco34325, w_eco34326, w_eco34327, w_eco34328, w_eco34329, w_eco34330, w_eco34331, w_eco34332, w_eco34333, w_eco34334, w_eco34335, w_eco34336, w_eco34337, w_eco34338, w_eco34339, w_eco34340, w_eco34341, w_eco34342, w_eco34343, w_eco34344, w_eco34345, w_eco34346, w_eco34347, w_eco34348, w_eco34349, w_eco34350, w_eco34351, w_eco34352, w_eco34353, w_eco34354, w_eco34355, w_eco34356, w_eco34357, w_eco34358, w_eco34359, w_eco34360, w_eco34361, w_eco34362, w_eco34363, w_eco34364, w_eco34365, w_eco34366, w_eco34367, w_eco34368, w_eco34369, w_eco34370, w_eco34371, w_eco34372, w_eco34373, w_eco34374, w_eco34375, w_eco34376, w_eco34377, w_eco34378, w_eco34379, w_eco34380, w_eco34381, w_eco34382, w_eco34383, w_eco34384, w_eco34385, w_eco34386, w_eco34387, w_eco34388, w_eco34389, w_eco34390, w_eco34391, w_eco34392, w_eco34393, w_eco34394, w_eco34395, w_eco34396, w_eco34397, w_eco34398, w_eco34399, w_eco34400, w_eco34401, w_eco34402, w_eco34403, w_eco34404, w_eco34405, w_eco34406, w_eco34407, w_eco34408, w_eco34409, w_eco34410, w_eco34411, w_eco34412, w_eco34413, w_eco34414, w_eco34415, w_eco34416, w_eco34417, w_eco34418, w_eco34419, w_eco34420, w_eco34421, w_eco34422, w_eco34423, w_eco34424, w_eco34425, w_eco34426, w_eco34427, w_eco34428, w_eco34429, w_eco34430, w_eco34431, w_eco34432, w_eco34433, w_eco34434, w_eco34435, w_eco34436, w_eco34437, w_eco34438, w_eco34439, w_eco34440, w_eco34441, w_eco34442, w_eco34443, w_eco34444, w_eco34445, w_eco34446, w_eco34447, w_eco34448, w_eco34449, w_eco34450, w_eco34451, w_eco34452, w_eco34453, w_eco34454, w_eco34455, w_eco34456, w_eco34457, w_eco34458, w_eco34459, w_eco34460, w_eco34461, w_eco34462, w_eco34463, w_eco34464, w_eco34465, w_eco34466, w_eco34467, w_eco34468, w_eco34469, w_eco34470, w_eco34471, w_eco34472, w_eco34473, w_eco34474, w_eco34475, w_eco34476, w_eco34477, w_eco34478, w_eco34479, w_eco34480, w_eco34481, w_eco34482, w_eco34483, w_eco34484, w_eco34485, w_eco34486, w_eco34487, w_eco34488, w_eco34489, w_eco34490, w_eco34491, w_eco34492, w_eco34493, w_eco34494, w_eco34495, w_eco34496, w_eco34497, w_eco34498, w_eco34499, w_eco34500, w_eco34501, w_eco34502, w_eco34503, w_eco34504, w_eco34505, w_eco34506, w_eco34507, w_eco34508, w_eco34509, w_eco34510, w_eco34511, w_eco34512, w_eco34513, w_eco34514, w_eco34515, w_eco34516, w_eco34517, w_eco34518, w_eco34519, w_eco34520, w_eco34521, w_eco34522, w_eco34523, w_eco34524, w_eco34525, w_eco34526, w_eco34527, w_eco34528, w_eco34529, w_eco34530, w_eco34531, w_eco34532, w_eco34533, w_eco34534, w_eco34535, w_eco34536, w_eco34537, w_eco34538, w_eco34539, w_eco34540, w_eco34541, w_eco34542, w_eco34543, w_eco34544, w_eco34545, w_eco34546, w_eco34547, w_eco34548, w_eco34549, w_eco34550, w_eco34551, w_eco34552, w_eco34553, w_eco34554, w_eco34555, w_eco34556, w_eco34557, w_eco34558, w_eco34559, w_eco34560, w_eco34561, w_eco34562, w_eco34563, w_eco34564, w_eco34565, w_eco34566, w_eco34567, w_eco34568, w_eco34569, w_eco34570, w_eco34571, w_eco34572, w_eco34573, w_eco34574, w_eco34575, w_eco34576, w_eco34577, w_eco34578, w_eco34579, w_eco34580, w_eco34581, w_eco34582, w_eco34583, w_eco34584, w_eco34585, w_eco34586, w_eco34587, w_eco34588, w_eco34589, w_eco34590, w_eco34591, w_eco34592, w_eco34593, w_eco34594, w_eco34595, w_eco34596, w_eco34597, w_eco34598, w_eco34599, w_eco34600, w_eco34601, w_eco34602, w_eco34603, w_eco34604, w_eco34605, w_eco34606, w_eco34607, w_eco34608, w_eco34609, w_eco34610, w_eco34611, w_eco34612, w_eco34613, w_eco34614, w_eco34615, w_eco34616, w_eco34617, w_eco34618, w_eco34619, w_eco34620, w_eco34621, w_eco34622, w_eco34623, w_eco34624, w_eco34625, w_eco34626, w_eco34627, w_eco34628, w_eco34629, w_eco34630, w_eco34631, w_eco34632, w_eco34633, w_eco34634, w_eco34635, w_eco34636, w_eco34637, w_eco34638, w_eco34639, w_eco34640, w_eco34641, w_eco34642, w_eco34643, w_eco34644, w_eco34645, w_eco34646, w_eco34647, w_eco34648, w_eco34649, w_eco34650, w_eco34651, w_eco34652, w_eco34653, w_eco34654, w_eco34655, w_eco34656, w_eco34657, w_eco34658, w_eco34659, w_eco34660, w_eco34661, w_eco34662, w_eco34663, w_eco34664, w_eco34665, w_eco34666, w_eco34667, w_eco34668, w_eco34669, w_eco34670, w_eco34671, w_eco34672, w_eco34673, w_eco34674, w_eco34675, w_eco34676, w_eco34677, w_eco34678, w_eco34679, w_eco34680, w_eco34681, w_eco34682, w_eco34683, w_eco34684, w_eco34685, w_eco34686, w_eco34687, w_eco34688, w_eco34689, w_eco34690, w_eco34691, w_eco34692, w_eco34693, w_eco34694, w_eco34695, w_eco34696, w_eco34697, w_eco34698, w_eco34699, w_eco34700, w_eco34701, w_eco34702, w_eco34703, w_eco34704, w_eco34705, w_eco34706, w_eco34707, w_eco34708, w_eco34709, w_eco34710, w_eco34711, w_eco34712, w_eco34713, w_eco34714, w_eco34715, w_eco34716, w_eco34717, w_eco34718, w_eco34719, w_eco34720, w_eco34721, w_eco34722, w_eco34723, w_eco34724, w_eco34725, w_eco34726, w_eco34727, w_eco34728, w_eco34729, w_eco34730, w_eco34731, w_eco34732, w_eco34733, w_eco34734, w_eco34735, w_eco34736, w_eco34737, w_eco34738, w_eco34739, w_eco34740, w_eco34741, w_eco34742, w_eco34743, w_eco34744, w_eco34745, w_eco34746, w_eco34747, w_eco34748, w_eco34749, w_eco34750, w_eco34751, w_eco34752, w_eco34753, w_eco34754, w_eco34755, w_eco34756, w_eco34757, w_eco34758, w_eco34759, w_eco34760, w_eco34761, w_eco34762, w_eco34763, w_eco34764, w_eco34765, w_eco34766, w_eco34767, w_eco34768, w_eco34769, w_eco34770, w_eco34771, w_eco34772, w_eco34773, w_eco34774, w_eco34775, w_eco34776, w_eco34777, w_eco34778, w_eco34779, w_eco34780, w_eco34781, w_eco34782, w_eco34783, w_eco34784, w_eco34785, w_eco34786, w_eco34787, w_eco34788, w_eco34789, w_eco34790, w_eco34791, w_eco34792, w_eco34793, w_eco34794, w_eco34795, w_eco34796, w_eco34797, w_eco34798, w_eco34799, w_eco34800, w_eco34801, w_eco34802, w_eco34803, w_eco34804, w_eco34805, w_eco34806, w_eco34807, w_eco34808, w_eco34809, w_eco34810, w_eco34811, w_eco34812, w_eco34813, w_eco34814, w_eco34815, w_eco34816, w_eco34817, w_eco34818, w_eco34819, w_eco34820, w_eco34821, w_eco34822, w_eco34823, w_eco34824, w_eco34825, w_eco34826, w_eco34827, w_eco34828, w_eco34829, w_eco34830, w_eco34831, w_eco34832, w_eco34833, w_eco34834, w_eco34835, w_eco34836, w_eco34837, w_eco34838, w_eco34839, w_eco34840, w_eco34841, w_eco34842, w_eco34843, w_eco34844, w_eco34845, w_eco34846, w_eco34847, w_eco34848, w_eco34849, w_eco34850, w_eco34851, w_eco34852, w_eco34853, w_eco34854, w_eco34855, w_eco34856, w_eco34857, w_eco34858, w_eco34859, w_eco34860, w_eco34861, w_eco34862, w_eco34863, w_eco34864, w_eco34865, w_eco34866, w_eco34867, w_eco34868, w_eco34869, w_eco34870, w_eco34871, w_eco34872, w_eco34873, w_eco34874, w_eco34875, w_eco34876, w_eco34877, w_eco34878, w_eco34879, w_eco34880, w_eco34881, w_eco34882, w_eco34883, w_eco34884, w_eco34885, w_eco34886, w_eco34887, w_eco34888, w_eco34889, w_eco34890, w_eco34891, w_eco34892, w_eco34893, w_eco34894, w_eco34895, w_eco34896, w_eco34897, w_eco34898, w_eco34899, w_eco34900, w_eco34901, w_eco34902, w_eco34903, w_eco34904, w_eco34905, w_eco34906, w_eco34907, w_eco34908, w_eco34909, w_eco34910, w_eco34911, w_eco34912, w_eco34913, w_eco34914, w_eco34915, w_eco34916, w_eco34917, w_eco34918, w_eco34919, w_eco34920, w_eco34921, w_eco34922, w_eco34923, w_eco34924, w_eco34925, w_eco34926, w_eco34927, w_eco34928, w_eco34929, w_eco34930, w_eco34931, w_eco34932, w_eco34933, w_eco34934, w_eco34935, w_eco34936, w_eco34937, w_eco34938, w_eco34939, w_eco34940, w_eco34941, w_eco34942, w_eco34943, w_eco34944, w_eco34945, w_eco34946, w_eco34947, w_eco34948, w_eco34949, w_eco34950, w_eco34951, w_eco34952, w_eco34953, w_eco34954, w_eco34955, w_eco34956, w_eco34957, w_eco34958, w_eco34959, w_eco34960, w_eco34961, w_eco34962, w_eco34963, w_eco34964, w_eco34965, w_eco34966, w_eco34967, w_eco34968, w_eco34969, w_eco34970, w_eco34971, w_eco34972, w_eco34973, w_eco34974, w_eco34975, w_eco34976, w_eco34977, w_eco34978, w_eco34979, w_eco34980, w_eco34981, w_eco34982, w_eco34983, w_eco34984, w_eco34985, w_eco34986, w_eco34987, w_eco34988, w_eco34989, w_eco34990, w_eco34991, w_eco34992, w_eco34993, w_eco34994, w_eco34995, w_eco34996, w_eco34997, w_eco34998, w_eco34999, w_eco35000, w_eco35001, w_eco35002, w_eco35003, w_eco35004, w_eco35005, w_eco35006, w_eco35007, w_eco35008, w_eco35009, w_eco35010, w_eco35011, w_eco35012, w_eco35013, w_eco35014, w_eco35015, w_eco35016, w_eco35017, w_eco35018, w_eco35019, w_eco35020, w_eco35021, w_eco35022, w_eco35023, w_eco35024, w_eco35025, w_eco35026, w_eco35027, w_eco35028, w_eco35029, w_eco35030, w_eco35031, w_eco35032, w_eco35033, w_eco35034, w_eco35035, w_eco35036, w_eco35037, w_eco35038, w_eco35039, w_eco35040, w_eco35041, w_eco35042, w_eco35043, w_eco35044, w_eco35045, w_eco35046, w_eco35047, w_eco35048, w_eco35049, w_eco35050, w_eco35051, w_eco35052, w_eco35053, w_eco35054, w_eco35055, w_eco35056, w_eco35057, w_eco35058, w_eco35059, w_eco35060, w_eco35061, w_eco35062, w_eco35063, w_eco35064, w_eco35065, w_eco35066, w_eco35067, w_eco35068, w_eco35069, w_eco35070, w_eco35071, w_eco35072, w_eco35073, w_eco35074, w_eco35075, w_eco35076, w_eco35077, w_eco35078, w_eco35079, w_eco35080, w_eco35081, w_eco35082, w_eco35083, w_eco35084, w_eco35085, w_eco35086, w_eco35087, w_eco35088, w_eco35089, w_eco35090, w_eco35091, w_eco35092, w_eco35093, w_eco35094, w_eco35095, w_eco35096, w_eco35097, w_eco35098, w_eco35099, w_eco35100, w_eco35101, w_eco35102, w_eco35103, w_eco35104, w_eco35105, w_eco35106, w_eco35107, w_eco35108, w_eco35109, w_eco35110, w_eco35111, w_eco35112, w_eco35113, w_eco35114, w_eco35115, w_eco35116, w_eco35117, w_eco35118, w_eco35119, w_eco35120, w_eco35121, w_eco35122, w_eco35123, w_eco35124, w_eco35125, w_eco35126, w_eco35127, w_eco35128, w_eco35129, w_eco35130, w_eco35131, w_eco35132, w_eco35133, w_eco35134, w_eco35135, w_eco35136, w_eco35137, w_eco35138, w_eco35139, w_eco35140, w_eco35141, w_eco35142, w_eco35143, w_eco35144, w_eco35145, w_eco35146, w_eco35147, w_eco35148, w_eco35149, w_eco35150, w_eco35151, w_eco35152, w_eco35153, w_eco35154, w_eco35155, w_eco35156, w_eco35157, w_eco35158, w_eco35159, w_eco35160, w_eco35161, w_eco35162, w_eco35163, w_eco35164, w_eco35165, w_eco35166, w_eco35167, w_eco35168, w_eco35169, w_eco35170, w_eco35171, w_eco35172, w_eco35173, w_eco35174, w_eco35175, w_eco35176, w_eco35177, w_eco35178, w_eco35179, w_eco35180, w_eco35181, w_eco35182, w_eco35183, w_eco35184, w_eco35185, w_eco35186, w_eco35187, w_eco35188, w_eco35189, w_eco35190, w_eco35191, w_eco35192, w_eco35193, w_eco35194, w_eco35195, w_eco35196, w_eco35197, w_eco35198, w_eco35199, w_eco35200, w_eco35201, w_eco35202, w_eco35203, w_eco35204, w_eco35205, w_eco35206, w_eco35207, w_eco35208, w_eco35209, w_eco35210, w_eco35211, w_eco35212, w_eco35213, w_eco35214, w_eco35215, w_eco35216, w_eco35217, w_eco35218, w_eco35219, w_eco35220, w_eco35221, w_eco35222, w_eco35223, w_eco35224, w_eco35225, w_eco35226, w_eco35227, w_eco35228, w_eco35229, w_eco35230, w_eco35231, w_eco35232, w_eco35233, w_eco35234, w_eco35235, w_eco35236, w_eco35237, w_eco35238, w_eco35239, w_eco35240, w_eco35241, w_eco35242, w_eco35243, w_eco35244, w_eco35245, w_eco35246, w_eco35247, w_eco35248, w_eco35249, w_eco35250, w_eco35251, w_eco35252, w_eco35253, w_eco35254, w_eco35255, w_eco35256, w_eco35257, w_eco35258, w_eco35259, w_eco35260, w_eco35261, w_eco35262, w_eco35263, w_eco35264, w_eco35265, w_eco35266, w_eco35267, w_eco35268, w_eco35269, w_eco35270, w_eco35271, w_eco35272, w_eco35273, w_eco35274, w_eco35275, w_eco35276, w_eco35277, w_eco35278, w_eco35279, w_eco35280, w_eco35281, w_eco35282, w_eco35283, w_eco35284, w_eco35285, w_eco35286, w_eco35287, w_eco35288, w_eco35289, w_eco35290, w_eco35291, w_eco35292, w_eco35293, w_eco35294, w_eco35295, w_eco35296, w_eco35297, w_eco35298, w_eco35299, w_eco35300, w_eco35301, w_eco35302, w_eco35303, w_eco35304, w_eco35305, w_eco35306, w_eco35307, w_eco35308, w_eco35309, w_eco35310, w_eco35311, w_eco35312, w_eco35313, w_eco35314, w_eco35315, w_eco35316, w_eco35317, w_eco35318, w_eco35319, w_eco35320, w_eco35321, w_eco35322, w_eco35323, w_eco35324, w_eco35325, w_eco35326, w_eco35327, w_eco35328, w_eco35329, w_eco35330, w_eco35331, w_eco35332, w_eco35333, w_eco35334, w_eco35335, w_eco35336, w_eco35337, w_eco35338, w_eco35339, w_eco35340, w_eco35341, w_eco35342, w_eco35343, w_eco35344, w_eco35345, w_eco35346, w_eco35347, w_eco35348, w_eco35349, w_eco35350, w_eco35351, w_eco35352, w_eco35353, w_eco35354, w_eco35355, w_eco35356, w_eco35357, w_eco35358, w_eco35359, w_eco35360, w_eco35361, w_eco35362, w_eco35363, w_eco35364, w_eco35365, w_eco35366, w_eco35367, w_eco35368, w_eco35369, w_eco35370, w_eco35371, w_eco35372, w_eco35373, w_eco35374, w_eco35375, w_eco35376, w_eco35377, w_eco35378, w_eco35379, w_eco35380, w_eco35381, w_eco35382, w_eco35383, w_eco35384, w_eco35385, w_eco35386, w_eco35387, w_eco35388, w_eco35389, w_eco35390, w_eco35391, w_eco35392, w_eco35393, w_eco35394, w_eco35395, w_eco35396, w_eco35397, w_eco35398, w_eco35399, w_eco35400, w_eco35401, w_eco35402, w_eco35403, w_eco35404, w_eco35405, w_eco35406, w_eco35407, w_eco35408, w_eco35409, w_eco35410, w_eco35411, w_eco35412, w_eco35413, w_eco35414, w_eco35415, w_eco35416, w_eco35417, w_eco35418, w_eco35419, w_eco35420, w_eco35421, w_eco35422, w_eco35423, w_eco35424, w_eco35425, w_eco35426, w_eco35427, w_eco35428, w_eco35429, w_eco35430, w_eco35431, w_eco35432, w_eco35433, w_eco35434, w_eco35435, w_eco35436, w_eco35437, w_eco35438, w_eco35439, w_eco35440, w_eco35441, w_eco35442, w_eco35443, w_eco35444, w_eco35445, w_eco35446, w_eco35447, w_eco35448, w_eco35449, w_eco35450, w_eco35451, w_eco35452, w_eco35453, w_eco35454, w_eco35455, w_eco35456, w_eco35457, w_eco35458, w_eco35459, w_eco35460, w_eco35461, w_eco35462, w_eco35463, w_eco35464, w_eco35465, w_eco35466, w_eco35467, w_eco35468, w_eco35469, w_eco35470, w_eco35471, w_eco35472, w_eco35473, w_eco35474, w_eco35475, w_eco35476, w_eco35477, w_eco35478, w_eco35479, w_eco35480, w_eco35481, w_eco35482, w_eco35483, w_eco35484, w_eco35485, w_eco35486, w_eco35487, w_eco35488, w_eco35489, w_eco35490, w_eco35491, w_eco35492, w_eco35493, w_eco35494, w_eco35495, w_eco35496, w_eco35497, w_eco35498, w_eco35499, w_eco35500, w_eco35501, w_eco35502, w_eco35503, w_eco35504, w_eco35505, w_eco35506, w_eco35507, w_eco35508, w_eco35509, w_eco35510, w_eco35511, w_eco35512, w_eco35513, w_eco35514, w_eco35515, w_eco35516, w_eco35517, w_eco35518, w_eco35519, w_eco35520, w_eco35521, w_eco35522, w_eco35523, w_eco35524, w_eco35525, w_eco35526, w_eco35527, w_eco35528, w_eco35529, w_eco35530, w_eco35531, w_eco35532, w_eco35533, w_eco35534, w_eco35535, w_eco35536, w_eco35537, w_eco35538, w_eco35539, w_eco35540, w_eco35541, w_eco35542, w_eco35543, w_eco35544, w_eco35545, w_eco35546, w_eco35547, w_eco35548, w_eco35549, w_eco35550, w_eco35551, w_eco35552, w_eco35553, w_eco35554, w_eco35555, w_eco35556, w_eco35557, w_eco35558, w_eco35559, w_eco35560, w_eco35561, w_eco35562, w_eco35563, w_eco35564, w_eco35565, w_eco35566, w_eco35567, w_eco35568, w_eco35569, w_eco35570, w_eco35571, w_eco35572, w_eco35573, w_eco35574, w_eco35575, w_eco35576, w_eco35577, w_eco35578, w_eco35579, w_eco35580, w_eco35581, w_eco35582, w_eco35583, w_eco35584, w_eco35585, w_eco35586, w_eco35587, w_eco35588, w_eco35589, w_eco35590, w_eco35591, w_eco35592, w_eco35593, w_eco35594, w_eco35595, w_eco35596, w_eco35597, w_eco35598, w_eco35599, w_eco35600, w_eco35601, w_eco35602, w_eco35603, w_eco35604, w_eco35605, w_eco35606, w_eco35607, w_eco35608, w_eco35609, w_eco35610, w_eco35611, w_eco35612, w_eco35613, w_eco35614, w_eco35615, w_eco35616, w_eco35617, w_eco35618, w_eco35619, w_eco35620, w_eco35621, w_eco35622, w_eco35623, w_eco35624, w_eco35625, w_eco35626, w_eco35627, w_eco35628, w_eco35629, w_eco35630, w_eco35631, w_eco35632, w_eco35633, w_eco35634, w_eco35635, w_eco35636, w_eco35637, w_eco35638, w_eco35639, w_eco35640, w_eco35641, w_eco35642, w_eco35643, w_eco35644, w_eco35645, w_eco35646, w_eco35647, w_eco35648, w_eco35649, w_eco35650, w_eco35651, w_eco35652, w_eco35653, w_eco35654, w_eco35655, w_eco35656, w_eco35657, w_eco35658, w_eco35659, w_eco35660, w_eco35661, w_eco35662, w_eco35663, w_eco35664, w_eco35665, w_eco35666, w_eco35667, w_eco35668, w_eco35669, w_eco35670, w_eco35671, w_eco35672, w_eco35673, w_eco35674, w_eco35675, w_eco35676, w_eco35677, w_eco35678, w_eco35679, w_eco35680, w_eco35681, w_eco35682, w_eco35683, w_eco35684, w_eco35685, w_eco35686, w_eco35687, w_eco35688, w_eco35689, w_eco35690, w_eco35691, w_eco35692, w_eco35693, w_eco35694, w_eco35695, w_eco35696, w_eco35697, w_eco35698, w_eco35699, w_eco35700, w_eco35701, w_eco35702, w_eco35703, w_eco35704, w_eco35705, w_eco35706, w_eco35707, w_eco35708, w_eco35709, w_eco35710, w_eco35711, w_eco35712, w_eco35713, w_eco35714, w_eco35715, w_eco35716, w_eco35717, w_eco35718, w_eco35719, w_eco35720, w_eco35721, w_eco35722, w_eco35723, w_eco35724, w_eco35725, w_eco35726, w_eco35727, w_eco35728, w_eco35729, w_eco35730, w_eco35731, w_eco35732, w_eco35733, w_eco35734, w_eco35735, w_eco35736, w_eco35737, w_eco35738, w_eco35739, w_eco35740, w_eco35741, w_eco35742, w_eco35743, w_eco35744, w_eco35745, w_eco35746, w_eco35747, w_eco35748, w_eco35749, w_eco35750, w_eco35751, w_eco35752, w_eco35753, w_eco35754, w_eco35755, w_eco35756, w_eco35757, w_eco35758, w_eco35759, w_eco35760, w_eco35761, w_eco35762, w_eco35763, w_eco35764, w_eco35765, w_eco35766, w_eco35767, w_eco35768, w_eco35769, w_eco35770, w_eco35771, w_eco35772, w_eco35773, w_eco35774, w_eco35775, w_eco35776, w_eco35777, w_eco35778, w_eco35779, w_eco35780, w_eco35781, w_eco35782, w_eco35783, w_eco35784, w_eco35785, w_eco35786, w_eco35787, w_eco35788, w_eco35789, w_eco35790, w_eco35791, w_eco35792, w_eco35793, w_eco35794, w_eco35795, w_eco35796, w_eco35797, w_eco35798, w_eco35799, w_eco35800, w_eco35801, w_eco35802, w_eco35803, w_eco35804, w_eco35805, w_eco35806, w_eco35807, w_eco35808, w_eco35809, w_eco35810, w_eco35811, w_eco35812, w_eco35813, w_eco35814, w_eco35815, w_eco35816, w_eco35817, w_eco35818, w_eco35819, w_eco35820, w_eco35821, w_eco35822, w_eco35823, w_eco35824, w_eco35825, w_eco35826, w_eco35827, w_eco35828, w_eco35829, w_eco35830, w_eco35831, w_eco35832, w_eco35833, w_eco35834, w_eco35835, w_eco35836, w_eco35837, w_eco35838, w_eco35839, w_eco35840, w_eco35841, w_eco35842, w_eco35843, w_eco35844, w_eco35845, w_eco35846, w_eco35847, w_eco35848, w_eco35849, w_eco35850, w_eco35851, w_eco35852, w_eco35853, w_eco35854, w_eco35855, w_eco35856, w_eco35857, w_eco35858, w_eco35859, w_eco35860, w_eco35861, w_eco35862, w_eco35863, w_eco35864, w_eco35865, w_eco35866, w_eco35867, w_eco35868, w_eco35869, w_eco35870, w_eco35871, w_eco35872, w_eco35873, w_eco35874, w_eco35875, w_eco35876, w_eco35877, w_eco35878, w_eco35879, w_eco35880, w_eco35881, w_eco35882, w_eco35883, w_eco35884, w_eco35885, w_eco35886, w_eco35887, w_eco35888, w_eco35889, w_eco35890, w_eco35891, w_eco35892, w_eco35893, w_eco35894, w_eco35895, w_eco35896, w_eco35897, w_eco35898, w_eco35899, w_eco35900, w_eco35901, w_eco35902, w_eco35903, w_eco35904, w_eco35905, w_eco35906, w_eco35907, w_eco35908, w_eco35909, w_eco35910, w_eco35911, w_eco35912, w_eco35913, w_eco35914, w_eco35915, w_eco35916, w_eco35917, w_eco35918, w_eco35919, w_eco35920, w_eco35921, w_eco35922, w_eco35923, w_eco35924, w_eco35925, w_eco35926, w_eco35927, w_eco35928, w_eco35929, w_eco35930, w_eco35931, w_eco35932, w_eco35933, w_eco35934, w_eco35935, w_eco35936, w_eco35937, w_eco35938, w_eco35939, w_eco35940, w_eco35941, w_eco35942, w_eco35943, w_eco35944, w_eco35945, w_eco35946, w_eco35947, w_eco35948, w_eco35949, w_eco35950, w_eco35951, w_eco35952, w_eco35953, w_eco35954, w_eco35955, w_eco35956, w_eco35957, w_eco35958, w_eco35959, w_eco35960, w_eco35961, w_eco35962, w_eco35963, w_eco35964, w_eco35965, w_eco35966, w_eco35967, w_eco35968, w_eco35969, w_eco35970, w_eco35971, w_eco35972, w_eco35973, w_eco35974, w_eco35975, w_eco35976, w_eco35977, w_eco35978, w_eco35979, w_eco35980, w_eco35981, w_eco35982, w_eco35983, w_eco35984, w_eco35985, w_eco35986, w_eco35987, w_eco35988, w_eco35989, w_eco35990, w_eco35991, w_eco35992, w_eco35993, w_eco35994, w_eco35995, w_eco35996, w_eco35997, w_eco35998, w_eco35999, w_eco36000, w_eco36001, w_eco36002, w_eco36003, w_eco36004, w_eco36005, w_eco36006, w_eco36007, w_eco36008, w_eco36009, w_eco36010, w_eco36011, w_eco36012, w_eco36013, w_eco36014, w_eco36015, w_eco36016, w_eco36017, w_eco36018, w_eco36019, w_eco36020, w_eco36021, w_eco36022, w_eco36023, w_eco36024, w_eco36025, w_eco36026, w_eco36027, w_eco36028, w_eco36029, w_eco36030, w_eco36031, w_eco36032, w_eco36033, w_eco36034, w_eco36035, w_eco36036, w_eco36037, w_eco36038, w_eco36039, w_eco36040, w_eco36041, w_eco36042, w_eco36043, w_eco36044, w_eco36045, w_eco36046, w_eco36047, w_eco36048, w_eco36049, w_eco36050, w_eco36051, w_eco36052, w_eco36053, w_eco36054, w_eco36055, w_eco36056, w_eco36057, w_eco36058, w_eco36059, w_eco36060, w_eco36061, w_eco36062, w_eco36063, w_eco36064, w_eco36065, w_eco36066, w_eco36067, w_eco36068, w_eco36069, w_eco36070, w_eco36071, w_eco36072, w_eco36073, w_eco36074, w_eco36075, w_eco36076, w_eco36077, w_eco36078, w_eco36079, w_eco36080, w_eco36081, w_eco36082, w_eco36083, w_eco36084, w_eco36085, w_eco36086, w_eco36087, w_eco36088, w_eco36089, w_eco36090, w_eco36091, w_eco36092, w_eco36093, w_eco36094, w_eco36095, w_eco36096, w_eco36097, w_eco36098, w_eco36099, w_eco36100, w_eco36101, w_eco36102, w_eco36103, w_eco36104, w_eco36105, w_eco36106, w_eco36107, w_eco36108, w_eco36109, w_eco36110, w_eco36111, w_eco36112, w_eco36113, w_eco36114, w_eco36115, w_eco36116, w_eco36117, w_eco36118, w_eco36119, w_eco36120, w_eco36121, w_eco36122, w_eco36123, w_eco36124, w_eco36125, w_eco36126, w_eco36127, w_eco36128, w_eco36129, w_eco36130, w_eco36131, w_eco36132, w_eco36133, w_eco36134, w_eco36135, w_eco36136, w_eco36137, w_eco36138, w_eco36139, w_eco36140, w_eco36141, w_eco36142, w_eco36143, w_eco36144, w_eco36145, w_eco36146, w_eco36147, w_eco36148, w_eco36149, w_eco36150, w_eco36151, w_eco36152, w_eco36153, w_eco36154, w_eco36155, w_eco36156, w_eco36157, w_eco36158, w_eco36159, w_eco36160, w_eco36161, w_eco36162, w_eco36163, w_eco36164, w_eco36165, w_eco36166, w_eco36167, w_eco36168, w_eco36169, w_eco36170, w_eco36171, w_eco36172, w_eco36173, w_eco36174, w_eco36175, w_eco36176, w_eco36177, w_eco36178, w_eco36179, w_eco36180, w_eco36181, w_eco36182, w_eco36183, w_eco36184, w_eco36185, w_eco36186, w_eco36187, w_eco36188, w_eco36189, w_eco36190, w_eco36191, w_eco36192, w_eco36193, w_eco36194, w_eco36195, w_eco36196, w_eco36197, w_eco36198, w_eco36199, w_eco36200, w_eco36201, w_eco36202, w_eco36203, w_eco36204, w_eco36205, w_eco36206, w_eco36207, w_eco36208, w_eco36209, w_eco36210, w_eco36211, w_eco36212, w_eco36213, w_eco36214, w_eco36215, w_eco36216, w_eco36217, w_eco36218, w_eco36219, w_eco36220, w_eco36221, w_eco36222, w_eco36223, w_eco36224, w_eco36225, w_eco36226, w_eco36227, w_eco36228, w_eco36229, w_eco36230, w_eco36231, w_eco36232, w_eco36233, w_eco36234, w_eco36235, w_eco36236, w_eco36237, w_eco36238, w_eco36239, w_eco36240, w_eco36241, w_eco36242, w_eco36243, w_eco36244, w_eco36245, w_eco36246, w_eco36247, w_eco36248, w_eco36249, w_eco36250, w_eco36251, w_eco36252, w_eco36253, w_eco36254, w_eco36255, w_eco36256, w_eco36257, w_eco36258, w_eco36259, w_eco36260, w_eco36261, w_eco36262, w_eco36263, w_eco36264, w_eco36265, w_eco36266, w_eco36267, w_eco36268, w_eco36269, w_eco36270, w_eco36271, w_eco36272, w_eco36273, w_eco36274, w_eco36275, w_eco36276, w_eco36277, w_eco36278, w_eco36279, w_eco36280, w_eco36281, w_eco36282, w_eco36283, w_eco36284, w_eco36285, w_eco36286, w_eco36287, w_eco36288, w_eco36289, w_eco36290, w_eco36291, w_eco36292, w_eco36293, w_eco36294, w_eco36295, w_eco36296, w_eco36297, w_eco36298, w_eco36299, w_eco36300, w_eco36301, w_eco36302, w_eco36303, w_eco36304, w_eco36305, w_eco36306, w_eco36307, w_eco36308, w_eco36309, w_eco36310, w_eco36311, w_eco36312, w_eco36313, w_eco36314, w_eco36315, w_eco36316, w_eco36317, w_eco36318, w_eco36319, w_eco36320, w_eco36321, w_eco36322, w_eco36323, w_eco36324, w_eco36325, w_eco36326, w_eco36327, w_eco36328, w_eco36329, w_eco36330, w_eco36331, w_eco36332, w_eco36333, w_eco36334, w_eco36335, w_eco36336, w_eco36337, w_eco36338, w_eco36339, w_eco36340, w_eco36341, w_eco36342, w_eco36343, w_eco36344, w_eco36345, w_eco36346, w_eco36347, w_eco36348, w_eco36349, w_eco36350, w_eco36351, w_eco36352, w_eco36353, w_eco36354, w_eco36355, w_eco36356, w_eco36357, w_eco36358, w_eco36359, w_eco36360, w_eco36361, w_eco36362, w_eco36363, w_eco36364, w_eco36365, w_eco36366, w_eco36367, w_eco36368, w_eco36369, w_eco36370, w_eco36371, w_eco36372, w_eco36373, w_eco36374, w_eco36375, w_eco36376, w_eco36377, w_eco36378, w_eco36379, w_eco36380, w_eco36381, w_eco36382, w_eco36383, w_eco36384, w_eco36385, w_eco36386, w_eco36387, w_eco36388, w_eco36389, w_eco36390, w_eco36391, w_eco36392, w_eco36393, w_eco36394, w_eco36395, w_eco36396, w_eco36397, w_eco36398, w_eco36399, w_eco36400, w_eco36401, w_eco36402, w_eco36403, w_eco36404, w_eco36405, w_eco36406, w_eco36407, w_eco36408, w_eco36409, w_eco36410, w_eco36411, w_eco36412, w_eco36413, w_eco36414, w_eco36415, w_eco36416, w_eco36417, w_eco36418, w_eco36419, w_eco36420, w_eco36421, w_eco36422, w_eco36423, w_eco36424, w_eco36425, w_eco36426, w_eco36427, w_eco36428, w_eco36429, w_eco36430, w_eco36431, w_eco36432, w_eco36433, w_eco36434, w_eco36435, w_eco36436, w_eco36437, w_eco36438, w_eco36439, w_eco36440, w_eco36441, w_eco36442, w_eco36443, w_eco36444, w_eco36445, w_eco36446, w_eco36447, w_eco36448, w_eco36449, w_eco36450, w_eco36451, w_eco36452, w_eco36453, w_eco36454, w_eco36455, w_eco36456, w_eco36457, w_eco36458, w_eco36459, w_eco36460, w_eco36461, w_eco36462, w_eco36463, w_eco36464, w_eco36465, w_eco36466, w_eco36467, w_eco36468, w_eco36469, w_eco36470, w_eco36471, w_eco36472, w_eco36473, w_eco36474, w_eco36475, w_eco36476, w_eco36477, w_eco36478, w_eco36479, w_eco36480, w_eco36481, w_eco36482, w_eco36483, w_eco36484, w_eco36485, w_eco36486, w_eco36487, w_eco36488, w_eco36489, w_eco36490, w_eco36491, w_eco36492, w_eco36493, w_eco36494, w_eco36495, w_eco36496, w_eco36497, w_eco36498, w_eco36499, w_eco36500, w_eco36501, w_eco36502, w_eco36503, w_eco36504, w_eco36505, w_eco36506, w_eco36507, w_eco36508, w_eco36509, w_eco36510, w_eco36511, w_eco36512, w_eco36513, w_eco36514, w_eco36515, w_eco36516, w_eco36517, w_eco36518, w_eco36519, w_eco36520, w_eco36521, w_eco36522, w_eco36523, w_eco36524, w_eco36525, w_eco36526, w_eco36527, w_eco36528, w_eco36529, w_eco36530, w_eco36531, w_eco36532, w_eco36533, w_eco36534, w_eco36535, w_eco36536, w_eco36537, w_eco36538, w_eco36539, w_eco36540, w_eco36541, w_eco36542, w_eco36543, w_eco36544, w_eco36545, w_eco36546, w_eco36547, w_eco36548, w_eco36549, w_eco36550, w_eco36551, w_eco36552, w_eco36553, w_eco36554, w_eco36555, w_eco36556, w_eco36557, w_eco36558, w_eco36559, w_eco36560, w_eco36561, w_eco36562, w_eco36563, w_eco36564, w_eco36565, w_eco36566, w_eco36567, w_eco36568, w_eco36569, w_eco36570, w_eco36571, w_eco36572, w_eco36573, w_eco36574, w_eco36575, w_eco36576, w_eco36577, w_eco36578, w_eco36579, w_eco36580, w_eco36581, w_eco36582, w_eco36583, w_eco36584, w_eco36585, w_eco36586, w_eco36587, w_eco36588, w_eco36589, w_eco36590, w_eco36591, w_eco36592, w_eco36593, w_eco36594, w_eco36595, w_eco36596, w_eco36597, w_eco36598, w_eco36599, w_eco36600, w_eco36601, w_eco36602, w_eco36603, w_eco36604, w_eco36605, w_eco36606, w_eco36607, w_eco36608, w_eco36609, w_eco36610, w_eco36611, w_eco36612, w_eco36613, w_eco36614, w_eco36615, w_eco36616, w_eco36617, w_eco36618, w_eco36619, w_eco36620, w_eco36621, w_eco36622, w_eco36623, w_eco36624, w_eco36625, w_eco36626, w_eco36627, w_eco36628, w_eco36629, w_eco36630, w_eco36631, w_eco36632, w_eco36633, w_eco36634, w_eco36635, w_eco36636, w_eco36637, w_eco36638, w_eco36639, w_eco36640, w_eco36641, w_eco36642, w_eco36643, w_eco36644, w_eco36645, w_eco36646, w_eco36647, w_eco36648, w_eco36649, w_eco36650, w_eco36651, w_eco36652, w_eco36653, w_eco36654, w_eco36655, w_eco36656, w_eco36657, w_eco36658, w_eco36659, w_eco36660, w_eco36661, w_eco36662, w_eco36663, w_eco36664, w_eco36665, w_eco36666, w_eco36667, w_eco36668, w_eco36669, w_eco36670, w_eco36671, w_eco36672, w_eco36673, w_eco36674, w_eco36675, w_eco36676, w_eco36677, w_eco36678, w_eco36679, w_eco36680, w_eco36681, w_eco36682, w_eco36683, w_eco36684, w_eco36685, w_eco36686, w_eco36687, w_eco36688, w_eco36689, w_eco36690, w_eco36691, w_eco36692, w_eco36693, w_eco36694, w_eco36695, w_eco36696, w_eco36697, w_eco36698, w_eco36699, w_eco36700, w_eco36701, w_eco36702, w_eco36703, w_eco36704, w_eco36705, w_eco36706, w_eco36707, w_eco36708, w_eco36709, w_eco36710, w_eco36711, w_eco36712, w_eco36713, w_eco36714, w_eco36715, w_eco36716, w_eco36717, w_eco36718, w_eco36719, w_eco36720, w_eco36721, w_eco36722, w_eco36723, w_eco36724, w_eco36725, w_eco36726, w_eco36727, w_eco36728, w_eco36729, w_eco36730, w_eco36731, w_eco36732, w_eco36733, w_eco36734, w_eco36735, w_eco36736, w_eco36737, w_eco36738, w_eco36739, w_eco36740, w_eco36741, w_eco36742, w_eco36743, w_eco36744, w_eco36745, w_eco36746, w_eco36747, w_eco36748, w_eco36749, w_eco36750, w_eco36751, w_eco36752, w_eco36753, w_eco36754, w_eco36755, w_eco36756, w_eco36757, w_eco36758, w_eco36759, w_eco36760, w_eco36761, w_eco36762, w_eco36763, w_eco36764, w_eco36765, w_eco36766, w_eco36767, w_eco36768, w_eco36769, w_eco36770, w_eco36771, w_eco36772, w_eco36773, w_eco36774, w_eco36775, w_eco36776, w_eco36777, w_eco36778, w_eco36779, w_eco36780, w_eco36781, w_eco36782, w_eco36783, w_eco36784, w_eco36785, w_eco36786, w_eco36787, w_eco36788, w_eco36789, w_eco36790, w_eco36791, w_eco36792, w_eco36793, w_eco36794, w_eco36795, w_eco36796, w_eco36797, w_eco36798, w_eco36799, w_eco36800, w_eco36801, w_eco36802, w_eco36803, w_eco36804, w_eco36805, w_eco36806, w_eco36807, w_eco36808, w_eco36809, w_eco36810, w_eco36811, w_eco36812, w_eco36813, w_eco36814, w_eco36815, w_eco36816, w_eco36817, w_eco36818, w_eco36819, w_eco36820, w_eco36821, w_eco36822, w_eco36823, w_eco36824, w_eco36825, w_eco36826, w_eco36827, w_eco36828, w_eco36829, w_eco36830, w_eco36831, w_eco36832, w_eco36833, w_eco36834, w_eco36835, w_eco36836, w_eco36837, w_eco36838, w_eco36839, w_eco36840, w_eco36841, w_eco36842, w_eco36843, w_eco36844, w_eco36845, w_eco36846, w_eco36847, w_eco36848, w_eco36849, w_eco36850, w_eco36851, w_eco36852, w_eco36853, w_eco36854, w_eco36855, w_eco36856, w_eco36857, w_eco36858, w_eco36859, w_eco36860, w_eco36861, w_eco36862, w_eco36863, w_eco36864, w_eco36865, w_eco36866, w_eco36867, w_eco36868, w_eco36869, w_eco36870, w_eco36871, w_eco36872, w_eco36873, w_eco36874, w_eco36875, w_eco36876, w_eco36877, w_eco36878, w_eco36879, w_eco36880, w_eco36881, w_eco36882, w_eco36883, w_eco36884, w_eco36885, w_eco36886, w_eco36887, w_eco36888, w_eco36889, w_eco36890, w_eco36891, w_eco36892, w_eco36893, w_eco36894, w_eco36895, w_eco36896, w_eco36897, w_eco36898, w_eco36899, w_eco36900, w_eco36901, w_eco36902, w_eco36903, w_eco36904, w_eco36905, w_eco36906, w_eco36907, w_eco36908, w_eco36909, w_eco36910, w_eco36911, w_eco36912, w_eco36913, w_eco36914, w_eco36915, w_eco36916, w_eco36917, w_eco36918, w_eco36919, w_eco36920, w_eco36921, w_eco36922, w_eco36923, w_eco36924, w_eco36925, w_eco36926, w_eco36927, w_eco36928, w_eco36929, w_eco36930, w_eco36931, w_eco36932, w_eco36933, w_eco36934, w_eco36935, w_eco36936, w_eco36937, w_eco36938, w_eco36939, w_eco36940, w_eco36941, w_eco36942, w_eco36943, w_eco36944, w_eco36945, w_eco36946, w_eco36947, w_eco36948, w_eco36949, w_eco36950, w_eco36951, w_eco36952, w_eco36953, w_eco36954, w_eco36955, w_eco36956, w_eco36957, w_eco36958, w_eco36959, w_eco36960, w_eco36961, w_eco36962, w_eco36963, w_eco36964, w_eco36965, w_eco36966, w_eco36967, w_eco36968, w_eco36969, w_eco36970, w_eco36971, w_eco36972, w_eco36973, w_eco36974, w_eco36975, w_eco36976, w_eco36977, w_eco36978, w_eco36979, w_eco36980, w_eco36981, w_eco36982, w_eco36983, w_eco36984, w_eco36985, w_eco36986, w_eco36987, w_eco36988, w_eco36989, w_eco36990, w_eco36991, w_eco36992, w_eco36993, w_eco36994, w_eco36995, w_eco36996, w_eco36997, w_eco36998, w_eco36999, w_eco37000, w_eco37001, w_eco37002, w_eco37003, w_eco37004, w_eco37005, w_eco37006, w_eco37007, w_eco37008, w_eco37009, w_eco37010, w_eco37011, w_eco37012, w_eco37013, w_eco37014, w_eco37015, w_eco37016, w_eco37017, w_eco37018, w_eco37019, w_eco37020, w_eco37021, w_eco37022, w_eco37023, w_eco37024, w_eco37025, w_eco37026, w_eco37027, w_eco37028, w_eco37029, w_eco37030, w_eco37031, w_eco37032, w_eco37033, w_eco37034, w_eco37035, w_eco37036, w_eco37037, w_eco37038, w_eco37039, w_eco37040, w_eco37041, w_eco37042, w_eco37043, w_eco37044, w_eco37045, w_eco37046, w_eco37047, w_eco37048, w_eco37049, w_eco37050, w_eco37051, w_eco37052, w_eco37053, w_eco37054, w_eco37055, w_eco37056, w_eco37057, w_eco37058, w_eco37059, w_eco37060, w_eco37061, w_eco37062, w_eco37063, w_eco37064, w_eco37065, w_eco37066, w_eco37067, w_eco37068, w_eco37069, w_eco37070, w_eco37071, w_eco37072, w_eco37073, w_eco37074, w_eco37075, w_eco37076, w_eco37077, w_eco37078, w_eco37079, w_eco37080, w_eco37081, w_eco37082, w_eco37083, w_eco37084, w_eco37085, w_eco37086, w_eco37087, w_eco37088, w_eco37089, w_eco37090, w_eco37091, w_eco37092, w_eco37093, w_eco37094, w_eco37095, w_eco37096, w_eco37097, w_eco37098, w_eco37099, w_eco37100, w_eco37101, w_eco37102, w_eco37103, w_eco37104, w_eco37105, w_eco37106, w_eco37107, w_eco37108, w_eco37109, w_eco37110, w_eco37111, w_eco37112, w_eco37113, w_eco37114, w_eco37115, w_eco37116, w_eco37117, w_eco37118, w_eco37119, w_eco37120, w_eco37121, w_eco37122, w_eco37123, w_eco37124, w_eco37125, w_eco37126, w_eco37127, w_eco37128, w_eco37129, w_eco37130, w_eco37131, w_eco37132, w_eco37133, w_eco37134, w_eco37135, w_eco37136, w_eco37137, w_eco37138, w_eco37139, w_eco37140, w_eco37141, w_eco37142, w_eco37143, w_eco37144, w_eco37145, w_eco37146, w_eco37147, w_eco37148, w_eco37149, w_eco37150, w_eco37151, w_eco37152, w_eco37153, w_eco37154, w_eco37155, w_eco37156, w_eco37157, w_eco37158, w_eco37159, w_eco37160, w_eco37161, w_eco37162, w_eco37163, w_eco37164, w_eco37165, w_eco37166, w_eco37167, w_eco37168, w_eco37169, w_eco37170, w_eco37171, w_eco37172, w_eco37173, w_eco37174, w_eco37175, w_eco37176, w_eco37177, w_eco37178, w_eco37179, w_eco37180, w_eco37181, w_eco37182, w_eco37183, w_eco37184, w_eco37185, w_eco37186, w_eco37187, w_eco37188, w_eco37189, w_eco37190, w_eco37191, w_eco37192, w_eco37193, w_eco37194, w_eco37195, w_eco37196, w_eco37197, w_eco37198, w_eco37199, w_eco37200, w_eco37201, w_eco37202, w_eco37203, w_eco37204, w_eco37205, w_eco37206, w_eco37207, w_eco37208, w_eco37209, w_eco37210, w_eco37211, w_eco37212, w_eco37213, w_eco37214, w_eco37215, w_eco37216, w_eco37217, w_eco37218, w_eco37219, w_eco37220, w_eco37221, w_eco37222, w_eco37223, w_eco37224, w_eco37225, w_eco37226, w_eco37227, w_eco37228, w_eco37229, w_eco37230, w_eco37231, w_eco37232, w_eco37233, w_eco37234, w_eco37235, w_eco37236, w_eco37237, w_eco37238, w_eco37239, w_eco37240, w_eco37241, w_eco37242, w_eco37243, w_eco37244, w_eco37245, w_eco37246, w_eco37247, w_eco37248, w_eco37249, w_eco37250, w_eco37251, w_eco37252, w_eco37253, w_eco37254, w_eco37255, w_eco37256, w_eco37257, w_eco37258, w_eco37259, w_eco37260, w_eco37261, w_eco37262, w_eco37263, w_eco37264, w_eco37265, w_eco37266, w_eco37267, w_eco37268, w_eco37269, w_eco37270, w_eco37271, w_eco37272, w_eco37273, w_eco37274, w_eco37275, w_eco37276, w_eco37277, w_eco37278, w_eco37279, w_eco37280, w_eco37281, w_eco37282, w_eco37283, w_eco37284, w_eco37285, w_eco37286, w_eco37287, w_eco37288, w_eco37289, w_eco37290, w_eco37291, w_eco37292, w_eco37293, w_eco37294, w_eco37295, w_eco37296, w_eco37297, w_eco37298, w_eco37299, w_eco37300, w_eco37301, w_eco37302, w_eco37303, w_eco37304, w_eco37305, w_eco37306, w_eco37307, w_eco37308, w_eco37309, w_eco37310, w_eco37311, w_eco37312, w_eco37313, w_eco37314, w_eco37315, w_eco37316, w_eco37317, w_eco37318, w_eco37319, w_eco37320, w_eco37321, w_eco37322, w_eco37323, w_eco37324, w_eco37325, w_eco37326, w_eco37327, w_eco37328, w_eco37329, w_eco37330, w_eco37331, w_eco37332, w_eco37333, w_eco37334, w_eco37335, w_eco37336, w_eco37337, w_eco37338, w_eco37339, w_eco37340, w_eco37341, w_eco37342, w_eco37343, w_eco37344, w_eco37345, w_eco37346, w_eco37347, w_eco37348, w_eco37349, w_eco37350, w_eco37351, w_eco37352, w_eco37353, w_eco37354, w_eco37355, w_eco37356, w_eco37357, w_eco37358, w_eco37359, w_eco37360, w_eco37361, w_eco37362, w_eco37363, w_eco37364, w_eco37365, w_eco37366, w_eco37367, w_eco37368, w_eco37369, w_eco37370, w_eco37371, w_eco37372, w_eco37373, w_eco37374, w_eco37375, w_eco37376, w_eco37377, w_eco37378, w_eco37379, w_eco37380, w_eco37381, w_eco37382, w_eco37383, w_eco37384, w_eco37385, w_eco37386, w_eco37387, w_eco37388, w_eco37389, w_eco37390, w_eco37391, w_eco37392, w_eco37393, w_eco37394, w_eco37395, w_eco37396, w_eco37397, w_eco37398, w_eco37399, w_eco37400, w_eco37401, w_eco37402, w_eco37403, w_eco37404, w_eco37405, w_eco37406, w_eco37407, w_eco37408, w_eco37409, w_eco37410, w_eco37411, w_eco37412, w_eco37413, w_eco37414, w_eco37415, w_eco37416, w_eco37417, w_eco37418, w_eco37419, w_eco37420, w_eco37421, w_eco37422, w_eco37423, w_eco37424, w_eco37425, w_eco37426, w_eco37427, w_eco37428, w_eco37429, w_eco37430, w_eco37431, w_eco37432, w_eco37433, w_eco37434, w_eco37435, w_eco37436, w_eco37437, w_eco37438, w_eco37439, w_eco37440, w_eco37441, w_eco37442, w_eco37443, w_eco37444, w_eco37445, w_eco37446, w_eco37447, w_eco37448, w_eco37449, w_eco37450, w_eco37451, w_eco37452, w_eco37453, w_eco37454, w_eco37455, w_eco37456, w_eco37457, w_eco37458, w_eco37459, w_eco37460, w_eco37461, w_eco37462, w_eco37463, w_eco37464, w_eco37465, w_eco37466, w_eco37467, w_eco37468, w_eco37469, w_eco37470, w_eco37471, w_eco37472, w_eco37473, w_eco37474, w_eco37475, w_eco37476, w_eco37477, w_eco37478, w_eco37479, w_eco37480, w_eco37481, w_eco37482, w_eco37483, w_eco37484, w_eco37485, w_eco37486, w_eco37487, w_eco37488, w_eco37489, w_eco37490, w_eco37491, w_eco37492, w_eco37493, w_eco37494, w_eco37495, w_eco37496, w_eco37497, w_eco37498, w_eco37499, w_eco37500, w_eco37501, w_eco37502, w_eco37503, w_eco37504, w_eco37505, w_eco37506, w_eco37507, w_eco37508, w_eco37509, w_eco37510, w_eco37511, w_eco37512, w_eco37513, w_eco37514, w_eco37515, w_eco37516, w_eco37517, w_eco37518, w_eco37519, w_eco37520, w_eco37521, w_eco37522, w_eco37523, w_eco37524, w_eco37525, w_eco37526, w_eco37527, w_eco37528, w_eco37529, w_eco37530, w_eco37531, w_eco37532, w_eco37533, w_eco37534, w_eco37535, w_eco37536, w_eco37537, w_eco37538, w_eco37539, w_eco37540, w_eco37541, w_eco37542, w_eco37543, w_eco37544, w_eco37545, w_eco37546, w_eco37547, w_eco37548, w_eco37549, w_eco37550, w_eco37551, w_eco37552, w_eco37553, w_eco37554, w_eco37555, w_eco37556, w_eco37557, w_eco37558, w_eco37559, w_eco37560, w_eco37561, w_eco37562, w_eco37563, w_eco37564, w_eco37565, w_eco37566, w_eco37567, w_eco37568, w_eco37569, w_eco37570, w_eco37571, w_eco37572, w_eco37573, w_eco37574, w_eco37575, w_eco37576, w_eco37577, w_eco37578, w_eco37579, w_eco37580, w_eco37581, w_eco37582, w_eco37583, w_eco37584, w_eco37585, w_eco37586, w_eco37587, w_eco37588, w_eco37589, w_eco37590, w_eco37591, w_eco37592, w_eco37593, w_eco37594, w_eco37595, w_eco37596, w_eco37597, w_eco37598, w_eco37599, w_eco37600, w_eco37601, w_eco37602, w_eco37603, w_eco37604, w_eco37605, w_eco37606, w_eco37607, w_eco37608, w_eco37609, w_eco37610, w_eco37611, w_eco37612, w_eco37613, w_eco37614, w_eco37615, w_eco37616, w_eco37617, w_eco37618, w_eco37619, w_eco37620, w_eco37621, w_eco37622, w_eco37623, w_eco37624, w_eco37625, w_eco37626, w_eco37627, w_eco37628, w_eco37629, w_eco37630, w_eco37631, w_eco37632, w_eco37633, w_eco37634, w_eco37635, w_eco37636, w_eco37637, w_eco37638, w_eco37639, w_eco37640, w_eco37641, w_eco37642, w_eco37643, w_eco37644, w_eco37645, w_eco37646, w_eco37647, w_eco37648, w_eco37649, w_eco37650, w_eco37651, w_eco37652, w_eco37653, w_eco37654, w_eco37655, w_eco37656, w_eco37657, w_eco37658, w_eco37659, w_eco37660, w_eco37661, w_eco37662, w_eco37663, w_eco37664, w_eco37665, w_eco37666, w_eco37667, w_eco37668, w_eco37669, w_eco37670, w_eco37671, w_eco37672, w_eco37673, w_eco37674, w_eco37675, w_eco37676, w_eco37677, w_eco37678, w_eco37679, w_eco37680, w_eco37681, w_eco37682, w_eco37683, w_eco37684, w_eco37685, w_eco37686, w_eco37687, w_eco37688, w_eco37689, w_eco37690, w_eco37691, w_eco37692, w_eco37693, w_eco37694, w_eco37695, w_eco37696, w_eco37697, w_eco37698, w_eco37699, w_eco37700, w_eco37701, w_eco37702, w_eco37703, w_eco37704, w_eco37705, w_eco37706, w_eco37707, w_eco37708, w_eco37709, w_eco37710, w_eco37711, w_eco37712, w_eco37713, w_eco37714, w_eco37715, w_eco37716, w_eco37717, w_eco37718, w_eco37719, w_eco37720, w_eco37721, w_eco37722, w_eco37723, w_eco37724, w_eco37725, w_eco37726, w_eco37727, w_eco37728, w_eco37729, w_eco37730, w_eco37731, w_eco37732, w_eco37733, w_eco37734, w_eco37735, w_eco37736, w_eco37737, w_eco37738, w_eco37739, w_eco37740, w_eco37741, w_eco37742, w_eco37743, w_eco37744, w_eco37745, w_eco37746, w_eco37747, w_eco37748, w_eco37749, w_eco37750, w_eco37751, w_eco37752, w_eco37753, w_eco37754, w_eco37755, w_eco37756, w_eco37757, w_eco37758, w_eco37759, w_eco37760, w_eco37761, w_eco37762, w_eco37763, w_eco37764, w_eco37765, w_eco37766, w_eco37767, w_eco37768, w_eco37769, w_eco37770, w_eco37771, w_eco37772, w_eco37773, w_eco37774, w_eco37775, w_eco37776, w_eco37777, w_eco37778, w_eco37779, w_eco37780, w_eco37781, w_eco37782, w_eco37783, w_eco37784, w_eco37785, w_eco37786, w_eco37787, w_eco37788, w_eco37789, w_eco37790, w_eco37791, w_eco37792, w_eco37793, w_eco37794, w_eco37795, w_eco37796, w_eco37797, w_eco37798, w_eco37799, w_eco37800, w_eco37801, w_eco37802, w_eco37803, w_eco37804, w_eco37805, w_eco37806, w_eco37807, w_eco37808, w_eco37809, w_eco37810, w_eco37811, w_eco37812, w_eco37813, w_eco37814, w_eco37815, w_eco37816, w_eco37817, w_eco37818, w_eco37819, w_eco37820, w_eco37821, w_eco37822, w_eco37823, w_eco37824, w_eco37825, w_eco37826, w_eco37827, w_eco37828, w_eco37829, w_eco37830, w_eco37831, w_eco37832, w_eco37833, w_eco37834, w_eco37835, w_eco37836, w_eco37837, w_eco37838, w_eco37839, w_eco37840, w_eco37841, w_eco37842, w_eco37843, w_eco37844, w_eco37845, w_eco37846, w_eco37847, w_eco37848, w_eco37849, w_eco37850, w_eco37851, w_eco37852, w_eco37853, w_eco37854, w_eco37855, w_eco37856, w_eco37857, w_eco37858, w_eco37859, w_eco37860, w_eco37861, w_eco37862, w_eco37863, w_eco37864, w_eco37865, w_eco37866, w_eco37867, w_eco37868, w_eco37869, w_eco37870, w_eco37871, w_eco37872, w_eco37873, w_eco37874, w_eco37875, w_eco37876, w_eco37877, w_eco37878, w_eco37879, w_eco37880, w_eco37881, w_eco37882, w_eco37883, w_eco37884, w_eco37885, w_eco37886, w_eco37887, w_eco37888, w_eco37889, w_eco37890, w_eco37891, w_eco37892, w_eco37893, w_eco37894, w_eco37895, w_eco37896, w_eco37897, w_eco37898, w_eco37899, w_eco37900, w_eco37901, w_eco37902, w_eco37903, w_eco37904, w_eco37905, w_eco37906, w_eco37907, w_eco37908, w_eco37909, w_eco37910, w_eco37911, w_eco37912, w_eco37913, w_eco37914, w_eco37915, w_eco37916, w_eco37917, w_eco37918, w_eco37919, w_eco37920, w_eco37921, w_eco37922, w_eco37923, w_eco37924, w_eco37925, w_eco37926, w_eco37927, w_eco37928, w_eco37929, w_eco37930, w_eco37931, w_eco37932, w_eco37933, w_eco37934, w_eco37935, w_eco37936, w_eco37937, w_eco37938, w_eco37939, w_eco37940, w_eco37941, w_eco37942, w_eco37943, w_eco37944, w_eco37945, w_eco37946, w_eco37947, w_eco37948, w_eco37949, w_eco37950, w_eco37951, w_eco37952, w_eco37953, w_eco37954, w_eco37955, w_eco37956, w_eco37957, w_eco37958, w_eco37959, w_eco37960, w_eco37961, w_eco37962, w_eco37963, w_eco37964, w_eco37965, w_eco37966, w_eco37967, w_eco37968, w_eco37969, w_eco37970, w_eco37971, w_eco37972, w_eco37973, w_eco37974, w_eco37975, w_eco37976, w_eco37977, w_eco37978, w_eco37979, w_eco37980, w_eco37981, w_eco37982, w_eco37983, w_eco37984, w_eco37985, w_eco37986, w_eco37987, w_eco37988, w_eco37989, w_eco37990, w_eco37991, w_eco37992, w_eco37993, w_eco37994, w_eco37995, w_eco37996, w_eco37997, w_eco37998, w_eco37999, w_eco38000, w_eco38001, w_eco38002, w_eco38003, w_eco38004, w_eco38005, w_eco38006, w_eco38007, w_eco38008, w_eco38009, w_eco38010, w_eco38011, w_eco38012, w_eco38013, w_eco38014, w_eco38015, w_eco38016, w_eco38017, w_eco38018, w_eco38019, w_eco38020, w_eco38021, w_eco38022, w_eco38023, w_eco38024, w_eco38025, w_eco38026, w_eco38027, w_eco38028, w_eco38029, w_eco38030, w_eco38031, w_eco38032, w_eco38033, w_eco38034, w_eco38035, w_eco38036, w_eco38037, w_eco38038, w_eco38039, w_eco38040, w_eco38041, w_eco38042, w_eco38043, w_eco38044, w_eco38045, w_eco38046, w_eco38047, w_eco38048, w_eco38049, w_eco38050, w_eco38051, w_eco38052, w_eco38053, w_eco38054, w_eco38055, w_eco38056, w_eco38057, w_eco38058, w_eco38059, w_eco38060, w_eco38061, w_eco38062, w_eco38063, w_eco38064, w_eco38065, w_eco38066, w_eco38067, w_eco38068, w_eco38069, w_eco38070, w_eco38071, w_eco38072, w_eco38073, w_eco38074, w_eco38075, w_eco38076, w_eco38077, w_eco38078, w_eco38079, w_eco38080, w_eco38081, w_eco38082, w_eco38083, w_eco38084, w_eco38085, w_eco38086, w_eco38087, w_eco38088, w_eco38089, w_eco38090, w_eco38091, w_eco38092, w_eco38093, w_eco38094, w_eco38095, w_eco38096, w_eco38097, w_eco38098, w_eco38099, w_eco38100, w_eco38101, w_eco38102, w_eco38103, w_eco38104, w_eco38105, w_eco38106, w_eco38107, w_eco38108, w_eco38109, w_eco38110, w_eco38111, w_eco38112, w_eco38113, w_eco38114, w_eco38115, w_eco38116, w_eco38117, w_eco38118, w_eco38119, w_eco38120, w_eco38121, w_eco38122, w_eco38123, w_eco38124, w_eco38125, w_eco38126, w_eco38127, w_eco38128, w_eco38129, w_eco38130, w_eco38131, w_eco38132, w_eco38133, w_eco38134, w_eco38135, w_eco38136, w_eco38137, w_eco38138, w_eco38139, w_eco38140, w_eco38141, w_eco38142, w_eco38143, w_eco38144, w_eco38145, w_eco38146, w_eco38147, w_eco38148, w_eco38149, w_eco38150, w_eco38151, w_eco38152, w_eco38153, w_eco38154, w_eco38155, w_eco38156, w_eco38157, w_eco38158, w_eco38159, w_eco38160, w_eco38161, w_eco38162, w_eco38163, w_eco38164, w_eco38165, w_eco38166, w_eco38167, w_eco38168, w_eco38169, w_eco38170, w_eco38171, w_eco38172, w_eco38173, w_eco38174, w_eco38175, w_eco38176, w_eco38177, w_eco38178, w_eco38179, w_eco38180, w_eco38181, w_eco38182, w_eco38183, w_eco38184, w_eco38185, w_eco38186, w_eco38187, w_eco38188, w_eco38189, w_eco38190, w_eco38191, w_eco38192, w_eco38193, w_eco38194, w_eco38195, w_eco38196, w_eco38197, w_eco38198, w_eco38199, w_eco38200, w_eco38201, w_eco38202, w_eco38203, w_eco38204, w_eco38205, w_eco38206, w_eco38207, w_eco38208, w_eco38209, w_eco38210, w_eco38211, w_eco38212, w_eco38213, w_eco38214, w_eco38215, w_eco38216, w_eco38217, w_eco38218, w_eco38219, w_eco38220, w_eco38221, w_eco38222, w_eco38223, w_eco38224, w_eco38225, w_eco38226, w_eco38227, w_eco38228, w_eco38229, w_eco38230, w_eco38231, w_eco38232, w_eco38233, w_eco38234, w_eco38235, w_eco38236, w_eco38237, w_eco38238, w_eco38239, w_eco38240, w_eco38241, w_eco38242, w_eco38243, w_eco38244, w_eco38245, w_eco38246, w_eco38247, w_eco38248, w_eco38249, w_eco38250, w_eco38251, w_eco38252, w_eco38253, w_eco38254, w_eco38255, w_eco38256, w_eco38257, w_eco38258, w_eco38259, w_eco38260, w_eco38261, w_eco38262, w_eco38263, w_eco38264, w_eco38265, w_eco38266, w_eco38267, w_eco38268, w_eco38269, w_eco38270, w_eco38271, w_eco38272, w_eco38273, w_eco38274, w_eco38275, w_eco38276, w_eco38277, w_eco38278, w_eco38279, w_eco38280, w_eco38281, w_eco38282, w_eco38283, w_eco38284, w_eco38285, w_eco38286, w_eco38287, w_eco38288, w_eco38289, w_eco38290, w_eco38291, w_eco38292, w_eco38293, w_eco38294, w_eco38295, w_eco38296, w_eco38297, w_eco38298, w_eco38299, w_eco38300, w_eco38301, w_eco38302, w_eco38303, w_eco38304, w_eco38305, w_eco38306, w_eco38307, w_eco38308, w_eco38309, w_eco38310, w_eco38311, w_eco38312, w_eco38313, w_eco38314, w_eco38315, w_eco38316, w_eco38317, w_eco38318, w_eco38319, w_eco38320, w_eco38321, w_eco38322, w_eco38323, w_eco38324, w_eco38325, w_eco38326, w_eco38327, w_eco38328, w_eco38329, w_eco38330, w_eco38331, w_eco38332, w_eco38333, w_eco38334, w_eco38335, w_eco38336, w_eco38337, w_eco38338, w_eco38339, w_eco38340, w_eco38341, w_eco38342, w_eco38343, w_eco38344, w_eco38345, w_eco38346, w_eco38347, w_eco38348, w_eco38349, w_eco38350, w_eco38351, w_eco38352, w_eco38353, w_eco38354, w_eco38355, w_eco38356, w_eco38357, w_eco38358, w_eco38359, w_eco38360, w_eco38361, w_eco38362, w_eco38363, w_eco38364, w_eco38365, w_eco38366, w_eco38367, w_eco38368, w_eco38369, w_eco38370, w_eco38371, w_eco38372, w_eco38373, w_eco38374, w_eco38375, w_eco38376, w_eco38377, w_eco38378, w_eco38379, w_eco38380, w_eco38381, w_eco38382, w_eco38383, w_eco38384, w_eco38385, w_eco38386, w_eco38387, w_eco38388, w_eco38389, w_eco38390, w_eco38391, w_eco38392, w_eco38393, w_eco38394, w_eco38395, w_eco38396, w_eco38397, w_eco38398, w_eco38399, w_eco38400, w_eco38401, w_eco38402, w_eco38403, w_eco38404, w_eco38405, w_eco38406, w_eco38407, w_eco38408, w_eco38409, w_eco38410, w_eco38411, w_eco38412, w_eco38413, w_eco38414, w_eco38415, w_eco38416, w_eco38417, w_eco38418, w_eco38419, w_eco38420, w_eco38421, w_eco38422, w_eco38423, w_eco38424, w_eco38425, w_eco38426, w_eco38427, w_eco38428, w_eco38429, w_eco38430, w_eco38431, w_eco38432, w_eco38433, w_eco38434, w_eco38435, w_eco38436, w_eco38437, w_eco38438, w_eco38439, w_eco38440, w_eco38441, w_eco38442, w_eco38443, w_eco38444, w_eco38445, w_eco38446, w_eco38447, w_eco38448, w_eco38449, w_eco38450, w_eco38451, w_eco38452, w_eco38453, w_eco38454, w_eco38455, w_eco38456, w_eco38457, w_eco38458, w_eco38459, w_eco38460, w_eco38461, w_eco38462, w_eco38463, w_eco38464, w_eco38465, w_eco38466, w_eco38467, w_eco38468, w_eco38469, w_eco38470, w_eco38471, w_eco38472, w_eco38473, w_eco38474, w_eco38475, w_eco38476, w_eco38477, w_eco38478, w_eco38479, w_eco38480, w_eco38481, w_eco38482, w_eco38483, w_eco38484, w_eco38485, w_eco38486, w_eco38487, w_eco38488, w_eco38489, w_eco38490, w_eco38491, w_eco38492, w_eco38493, w_eco38494, w_eco38495, w_eco38496, w_eco38497, w_eco38498, w_eco38499, w_eco38500, w_eco38501, w_eco38502, w_eco38503, w_eco38504, w_eco38505, w_eco38506, w_eco38507, w_eco38508, w_eco38509, w_eco38510, w_eco38511, w_eco38512, w_eco38513, w_eco38514, w_eco38515, w_eco38516, w_eco38517, w_eco38518, w_eco38519, w_eco38520, w_eco38521, w_eco38522, w_eco38523, w_eco38524, w_eco38525, w_eco38526, w_eco38527, w_eco38528, w_eco38529, w_eco38530, w_eco38531, w_eco38532, w_eco38533, w_eco38534, w_eco38535, w_eco38536, w_eco38537, w_eco38538, w_eco38539, w_eco38540, w_eco38541, w_eco38542, w_eco38543, w_eco38544, w_eco38545, w_eco38546, w_eco38547, w_eco38548, w_eco38549, w_eco38550, w_eco38551, w_eco38552, w_eco38553, w_eco38554, w_eco38555, w_eco38556, w_eco38557, w_eco38558, w_eco38559, w_eco38560, w_eco38561, w_eco38562, w_eco38563, w_eco38564, w_eco38565, w_eco38566, w_eco38567, w_eco38568, w_eco38569, w_eco38570, w_eco38571, w_eco38572, w_eco38573, w_eco38574, w_eco38575, w_eco38576, w_eco38577, w_eco38578, w_eco38579, w_eco38580, w_eco38581, w_eco38582, w_eco38583, w_eco38584, w_eco38585, w_eco38586, w_eco38587, w_eco38588, w_eco38589, w_eco38590, w_eco38591, w_eco38592, w_eco38593, w_eco38594, w_eco38595, w_eco38596, w_eco38597, w_eco38598, w_eco38599, w_eco38600, w_eco38601, w_eco38602, w_eco38603, w_eco38604, w_eco38605, w_eco38606, w_eco38607, w_eco38608, w_eco38609, w_eco38610, w_eco38611, w_eco38612, w_eco38613, w_eco38614, w_eco38615, w_eco38616, w_eco38617, w_eco38618, w_eco38619, w_eco38620, w_eco38621, w_eco38622, w_eco38623, w_eco38624, w_eco38625, w_eco38626, w_eco38627, w_eco38628, w_eco38629, w_eco38630, w_eco38631, w_eco38632, w_eco38633, w_eco38634, w_eco38635, w_eco38636, w_eco38637, w_eco38638, w_eco38639, w_eco38640, w_eco38641, w_eco38642, w_eco38643, w_eco38644, w_eco38645, w_eco38646, w_eco38647, w_eco38648, w_eco38649, w_eco38650, w_eco38651, w_eco38652, w_eco38653, w_eco38654, w_eco38655, w_eco38656, w_eco38657, w_eco38658, w_eco38659, w_eco38660, w_eco38661, w_eco38662, w_eco38663, w_eco38664, w_eco38665, w_eco38666, w_eco38667, w_eco38668, w_eco38669, w_eco38670, w_eco38671, w_eco38672, w_eco38673, w_eco38674, w_eco38675, w_eco38676, w_eco38677, w_eco38678, w_eco38679, w_eco38680, w_eco38681, w_eco38682, w_eco38683, w_eco38684, w_eco38685, w_eco38686, w_eco38687, w_eco38688, w_eco38689, w_eco38690, w_eco38691, w_eco38692, w_eco38693, w_eco38694, w_eco38695, w_eco38696, w_eco38697, w_eco38698, w_eco38699, w_eco38700, w_eco38701, w_eco38702, w_eco38703, w_eco38704, w_eco38705, w_eco38706, w_eco38707, w_eco38708, w_eco38709, w_eco38710, w_eco38711, w_eco38712, w_eco38713, w_eco38714, w_eco38715, w_eco38716, w_eco38717, w_eco38718, w_eco38719, w_eco38720, w_eco38721, w_eco38722, w_eco38723, w_eco38724, w_eco38725, w_eco38726, w_eco38727, w_eco38728, w_eco38729, w_eco38730, w_eco38731, w_eco38732, w_eco38733, w_eco38734, w_eco38735, w_eco38736, w_eco38737, w_eco38738, w_eco38739, w_eco38740, w_eco38741, w_eco38742, w_eco38743, w_eco38744, w_eco38745, w_eco38746, w_eco38747, w_eco38748, w_eco38749, w_eco38750, w_eco38751, w_eco38752, w_eco38753, w_eco38754, w_eco38755, w_eco38756, w_eco38757, w_eco38758, w_eco38759, w_eco38760, w_eco38761, w_eco38762, w_eco38763, w_eco38764, w_eco38765, w_eco38766, w_eco38767, w_eco38768, w_eco38769, w_eco38770, w_eco38771, w_eco38772, w_eco38773, w_eco38774, w_eco38775, w_eco38776, w_eco38777, w_eco38778, w_eco38779, w_eco38780, w_eco38781, w_eco38782, w_eco38783, w_eco38784, w_eco38785, w_eco38786, w_eco38787, w_eco38788, w_eco38789, w_eco38790, w_eco38791, w_eco38792, w_eco38793, w_eco38794, w_eco38795, w_eco38796, w_eco38797, w_eco38798, w_eco38799, w_eco38800, w_eco38801, w_eco38802, w_eco38803, w_eco38804, w_eco38805, w_eco38806, w_eco38807, w_eco38808, w_eco38809, w_eco38810, w_eco38811, w_eco38812, w_eco38813, w_eco38814, w_eco38815, w_eco38816, w_eco38817, w_eco38818, w_eco38819, w_eco38820, w_eco38821, w_eco38822, w_eco38823, w_eco38824, w_eco38825, w_eco38826, w_eco38827, w_eco38828, w_eco38829, w_eco38830, w_eco38831, w_eco38832, w_eco38833, w_eco38834, w_eco38835, w_eco38836, w_eco38837, w_eco38838, w_eco38839, w_eco38840, w_eco38841, w_eco38842, w_eco38843, w_eco38844, w_eco38845, w_eco38846, w_eco38847, w_eco38848, w_eco38849, w_eco38850, w_eco38851, w_eco38852, w_eco38853, w_eco38854, w_eco38855, w_eco38856, w_eco38857, w_eco38858, w_eco38859, w_eco38860, w_eco38861, w_eco38862, w_eco38863, w_eco38864, w_eco38865, w_eco38866, w_eco38867, w_eco38868, w_eco38869, w_eco38870, w_eco38871, w_eco38872, w_eco38873, w_eco38874, w_eco38875, w_eco38876, w_eco38877, w_eco38878, w_eco38879, w_eco38880, w_eco38881, w_eco38882, w_eco38883, w_eco38884, w_eco38885, w_eco38886, w_eco38887, w_eco38888, w_eco38889, w_eco38890, w_eco38891, w_eco38892, w_eco38893, w_eco38894, w_eco38895, w_eco38896, w_eco38897, w_eco38898, w_eco38899, w_eco38900, w_eco38901, w_eco38902, w_eco38903, w_eco38904, w_eco38905, w_eco38906, w_eco38907, w_eco38908, w_eco38909, w_eco38910, w_eco38911, w_eco38912, w_eco38913, w_eco38914, w_eco38915, w_eco38916, w_eco38917, w_eco38918, w_eco38919, w_eco38920, w_eco38921, w_eco38922, w_eco38923, w_eco38924, w_eco38925, w_eco38926, w_eco38927, w_eco38928, w_eco38929, w_eco38930, w_eco38931, w_eco38932, w_eco38933, w_eco38934, w_eco38935, w_eco38936, w_eco38937, w_eco38938, w_eco38939, w_eco38940, w_eco38941, w_eco38942, w_eco38943, w_eco38944, w_eco38945, w_eco38946, w_eco38947, w_eco38948, w_eco38949, w_eco38950, w_eco38951, w_eco38952, w_eco38953, w_eco38954, w_eco38955, w_eco38956, w_eco38957, w_eco38958, w_eco38959, w_eco38960, w_eco38961, w_eco38962, w_eco38963, w_eco38964, w_eco38965, w_eco38966, w_eco38967, w_eco38968, w_eco38969, w_eco38970, w_eco38971, w_eco38972, w_eco38973, w_eco38974, w_eco38975, w_eco38976, w_eco38977, w_eco38978, w_eco38979, w_eco38980, w_eco38981, w_eco38982, w_eco38983, w_eco38984, w_eco38985, w_eco38986, w_eco38987, w_eco38988, w_eco38989, w_eco38990, w_eco38991, w_eco38992, w_eco38993, w_eco38994, w_eco38995, w_eco38996, w_eco38997, w_eco38998, w_eco38999, w_eco39000, w_eco39001, w_eco39002, w_eco39003, w_eco39004, w_eco39005, w_eco39006, w_eco39007, w_eco39008, w_eco39009, w_eco39010, w_eco39011, w_eco39012, w_eco39013, w_eco39014, w_eco39015, w_eco39016, w_eco39017, w_eco39018, w_eco39019, w_eco39020, w_eco39021, w_eco39022, w_eco39023, w_eco39024, w_eco39025, w_eco39026, w_eco39027, w_eco39028, w_eco39029, w_eco39030, w_eco39031, w_eco39032, w_eco39033, w_eco39034, w_eco39035, w_eco39036, w_eco39037, w_eco39038, w_eco39039, w_eco39040, w_eco39041, w_eco39042, w_eco39043, w_eco39044, w_eco39045, w_eco39046, w_eco39047, w_eco39048, w_eco39049, w_eco39050, w_eco39051, w_eco39052, w_eco39053, w_eco39054, w_eco39055, w_eco39056, w_eco39057, w_eco39058, w_eco39059, w_eco39060, w_eco39061, w_eco39062, w_eco39063, w_eco39064, w_eco39065, w_eco39066, w_eco39067, w_eco39068, w_eco39069, w_eco39070, w_eco39071, w_eco39072, w_eco39073, w_eco39074, w_eco39075, w_eco39076, w_eco39077, w_eco39078, w_eco39079, w_eco39080, w_eco39081, w_eco39082, w_eco39083, w_eco39084, w_eco39085, w_eco39086, w_eco39087, w_eco39088, w_eco39089, w_eco39090, w_eco39091, w_eco39092, w_eco39093, w_eco39094, w_eco39095, w_eco39096, w_eco39097, w_eco39098, w_eco39099, w_eco39100, w_eco39101, w_eco39102, w_eco39103, w_eco39104, w_eco39105, w_eco39106, w_eco39107, w_eco39108, w_eco39109, w_eco39110, w_eco39111, w_eco39112, w_eco39113, w_eco39114, w_eco39115, w_eco39116, w_eco39117, w_eco39118, w_eco39119, w_eco39120, w_eco39121, w_eco39122, w_eco39123, w_eco39124, w_eco39125, w_eco39126, w_eco39127, w_eco39128, w_eco39129, w_eco39130, w_eco39131, w_eco39132, w_eco39133, w_eco39134, w_eco39135, w_eco39136, w_eco39137, w_eco39138, w_eco39139, w_eco39140, w_eco39141, w_eco39142, w_eco39143, w_eco39144, w_eco39145, w_eco39146, w_eco39147, w_eco39148, w_eco39149, w_eco39150, w_eco39151, w_eco39152, w_eco39153, w_eco39154, w_eco39155, w_eco39156, w_eco39157, w_eco39158, w_eco39159, w_eco39160, w_eco39161, w_eco39162, w_eco39163, w_eco39164, w_eco39165, w_eco39166, w_eco39167, w_eco39168, w_eco39169, w_eco39170, w_eco39171, w_eco39172, w_eco39173, w_eco39174, w_eco39175, w_eco39176, w_eco39177, w_eco39178, w_eco39179, w_eco39180, w_eco39181, w_eco39182, w_eco39183, w_eco39184, w_eco39185, w_eco39186, w_eco39187, w_eco39188, w_eco39189, w_eco39190, w_eco39191, w_eco39192, w_eco39193, w_eco39194, w_eco39195, w_eco39196, w_eco39197, w_eco39198, w_eco39199, w_eco39200, w_eco39201, w_eco39202, w_eco39203, w_eco39204, w_eco39205, w_eco39206, w_eco39207, w_eco39208, w_eco39209, w_eco39210, w_eco39211, w_eco39212, w_eco39213, w_eco39214, w_eco39215, w_eco39216, w_eco39217, w_eco39218, w_eco39219, w_eco39220, w_eco39221, w_eco39222, w_eco39223, w_eco39224, w_eco39225, w_eco39226, w_eco39227, w_eco39228, w_eco39229, w_eco39230, w_eco39231, w_eco39232, w_eco39233, w_eco39234, w_eco39235, w_eco39236, w_eco39237, w_eco39238, w_eco39239, w_eco39240, w_eco39241, w_eco39242, w_eco39243, w_eco39244, w_eco39245, w_eco39246, w_eco39247, w_eco39248, w_eco39249, w_eco39250, w_eco39251, w_eco39252, w_eco39253, w_eco39254, w_eco39255, w_eco39256, w_eco39257, w_eco39258, w_eco39259, w_eco39260, w_eco39261, w_eco39262, w_eco39263, w_eco39264, w_eco39265, w_eco39266, w_eco39267, w_eco39268, w_eco39269, w_eco39270, w_eco39271, w_eco39272, w_eco39273, w_eco39274, w_eco39275, w_eco39276, w_eco39277, w_eco39278, w_eco39279, w_eco39280, w_eco39281, w_eco39282, w_eco39283, w_eco39284, w_eco39285, w_eco39286, w_eco39287, w_eco39288, w_eco39289, w_eco39290, w_eco39291, w_eco39292, w_eco39293, w_eco39294, w_eco39295, w_eco39296, w_eco39297, w_eco39298, w_eco39299, w_eco39300, w_eco39301, w_eco39302, w_eco39303, w_eco39304, w_eco39305, w_eco39306, w_eco39307, w_eco39308, w_eco39309, w_eco39310, w_eco39311, w_eco39312, w_eco39313, w_eco39314, w_eco39315, w_eco39316, w_eco39317, w_eco39318, w_eco39319, w_eco39320, w_eco39321, w_eco39322, w_eco39323, w_eco39324, w_eco39325, w_eco39326, w_eco39327, w_eco39328, w_eco39329, w_eco39330, w_eco39331, w_eco39332, w_eco39333, w_eco39334, w_eco39335, w_eco39336, w_eco39337, w_eco39338, w_eco39339, w_eco39340, w_eco39341, w_eco39342, w_eco39343, w_eco39344, w_eco39345, w_eco39346, w_eco39347, w_eco39348, w_eco39349, w_eco39350, w_eco39351, w_eco39352, w_eco39353, w_eco39354, w_eco39355, w_eco39356, w_eco39357, w_eco39358, w_eco39359, w_eco39360, w_eco39361, w_eco39362, w_eco39363, w_eco39364, w_eco39365, w_eco39366, w_eco39367, w_eco39368, w_eco39369, w_eco39370, w_eco39371, w_eco39372, w_eco39373, w_eco39374, w_eco39375, w_eco39376, w_eco39377, w_eco39378, w_eco39379, w_eco39380, w_eco39381, w_eco39382, w_eco39383, w_eco39384, w_eco39385, w_eco39386, w_eco39387, w_eco39388, w_eco39389, w_eco39390, w_eco39391, w_eco39392, w_eco39393, w_eco39394, w_eco39395, w_eco39396, w_eco39397, w_eco39398, w_eco39399, w_eco39400, w_eco39401, w_eco39402, w_eco39403, w_eco39404, w_eco39405, w_eco39406, w_eco39407, w_eco39408, w_eco39409, w_eco39410, w_eco39411, w_eco39412, w_eco39413, w_eco39414, w_eco39415, w_eco39416, w_eco39417, w_eco39418, w_eco39419, w_eco39420, w_eco39421, w_eco39422, w_eco39423, w_eco39424, w_eco39425, w_eco39426, w_eco39427, w_eco39428, w_eco39429, w_eco39430, w_eco39431, w_eco39432, w_eco39433, w_eco39434, w_eco39435, w_eco39436, w_eco39437, w_eco39438, w_eco39439, w_eco39440, w_eco39441, w_eco39442, w_eco39443, w_eco39444, w_eco39445, w_eco39446, w_eco39447, w_eco39448, w_eco39449, w_eco39450, w_eco39451, w_eco39452, w_eco39453, w_eco39454, w_eco39455, w_eco39456, w_eco39457, w_eco39458, w_eco39459, w_eco39460, w_eco39461, w_eco39462, w_eco39463, w_eco39464, w_eco39465, w_eco39466, w_eco39467, w_eco39468, w_eco39469, w_eco39470, w_eco39471, w_eco39472, w_eco39473, w_eco39474, w_eco39475, w_eco39476, w_eco39477, w_eco39478, w_eco39479, w_eco39480, w_eco39481, w_eco39482, w_eco39483, w_eco39484, w_eco39485, w_eco39486, w_eco39487, w_eco39488, w_eco39489, w_eco39490, w_eco39491, w_eco39492, w_eco39493, w_eco39494, w_eco39495, w_eco39496, w_eco39497, w_eco39498, w_eco39499, w_eco39500, w_eco39501, w_eco39502, w_eco39503, w_eco39504, w_eco39505, w_eco39506, w_eco39507, w_eco39508, w_eco39509, w_eco39510, w_eco39511, w_eco39512, w_eco39513, w_eco39514, w_eco39515, w_eco39516, w_eco39517, w_eco39518, w_eco39519, w_eco39520, w_eco39521, w_eco39522, w_eco39523, w_eco39524, w_eco39525, w_eco39526, w_eco39527, w_eco39528, w_eco39529, w_eco39530, w_eco39531, w_eco39532, w_eco39533, w_eco39534, w_eco39535, w_eco39536, w_eco39537, w_eco39538, w_eco39539, w_eco39540, w_eco39541, w_eco39542, w_eco39543, w_eco39544, w_eco39545, w_eco39546, w_eco39547, w_eco39548, w_eco39549, w_eco39550, w_eco39551, w_eco39552, w_eco39553, w_eco39554, w_eco39555, w_eco39556, w_eco39557, w_eco39558, w_eco39559, w_eco39560, w_eco39561, w_eco39562, w_eco39563, w_eco39564, w_eco39565, w_eco39566, w_eco39567, w_eco39568, w_eco39569, w_eco39570, w_eco39571, w_eco39572, w_eco39573, w_eco39574, w_eco39575, w_eco39576, w_eco39577, w_eco39578, w_eco39579, w_eco39580, w_eco39581, w_eco39582, w_eco39583, w_eco39584, w_eco39585, w_eco39586, w_eco39587, w_eco39588, w_eco39589, w_eco39590, w_eco39591, w_eco39592, w_eco39593, w_eco39594, w_eco39595, w_eco39596, w_eco39597, w_eco39598, w_eco39599, w_eco39600, w_eco39601, w_eco39602, w_eco39603, w_eco39604, w_eco39605, w_eco39606, w_eco39607, w_eco39608, w_eco39609, w_eco39610, w_eco39611, w_eco39612, w_eco39613, w_eco39614, w_eco39615, w_eco39616, w_eco39617, w_eco39618, w_eco39619, w_eco39620, w_eco39621, w_eco39622, w_eco39623, w_eco39624, w_eco39625, w_eco39626, w_eco39627, w_eco39628, w_eco39629, w_eco39630, w_eco39631, w_eco39632, w_eco39633, w_eco39634, w_eco39635, w_eco39636, w_eco39637, w_eco39638, w_eco39639, w_eco39640, w_eco39641, w_eco39642, w_eco39643, w_eco39644, w_eco39645, w_eco39646, w_eco39647, w_eco39648, w_eco39649, w_eco39650, w_eco39651, w_eco39652, w_eco39653, w_eco39654, w_eco39655, w_eco39656, w_eco39657, w_eco39658, w_eco39659, w_eco39660, w_eco39661, w_eco39662, w_eco39663, w_eco39664, w_eco39665, w_eco39666, w_eco39667, w_eco39668, w_eco39669, w_eco39670, w_eco39671, w_eco39672, w_eco39673, w_eco39674, w_eco39675, w_eco39676, w_eco39677, w_eco39678, w_eco39679, w_eco39680, w_eco39681, w_eco39682, w_eco39683, w_eco39684, w_eco39685, w_eco39686, w_eco39687, w_eco39688, w_eco39689, w_eco39690, w_eco39691, w_eco39692, w_eco39693, w_eco39694, w_eco39695, w_eco39696, w_eco39697, w_eco39698, w_eco39699, w_eco39700, w_eco39701, w_eco39702, w_eco39703, w_eco39704, w_eco39705, w_eco39706, w_eco39707, w_eco39708, w_eco39709, w_eco39710, w_eco39711, w_eco39712, w_eco39713, w_eco39714, w_eco39715, w_eco39716, w_eco39717, w_eco39718, w_eco39719, w_eco39720, w_eco39721, w_eco39722, w_eco39723, w_eco39724, w_eco39725, w_eco39726, w_eco39727, w_eco39728, w_eco39729, w_eco39730, w_eco39731, w_eco39732, w_eco39733, w_eco39734, w_eco39735, w_eco39736, w_eco39737, w_eco39738, w_eco39739, w_eco39740, w_eco39741, w_eco39742, w_eco39743, w_eco39744, w_eco39745, w_eco39746, w_eco39747, w_eco39748, w_eco39749, w_eco39750, w_eco39751, w_eco39752, w_eco39753, w_eco39754, w_eco39755, w_eco39756, w_eco39757, w_eco39758, w_eco39759, w_eco39760, w_eco39761, w_eco39762, w_eco39763, w_eco39764, w_eco39765, w_eco39766, w_eco39767, w_eco39768, w_eco39769, w_eco39770, w_eco39771, w_eco39772, w_eco39773, w_eco39774, w_eco39775, w_eco39776, w_eco39777, w_eco39778, w_eco39779, w_eco39780, w_eco39781, w_eco39782, w_eco39783, w_eco39784, w_eco39785, w_eco39786, w_eco39787, w_eco39788, w_eco39789, w_eco39790, w_eco39791, w_eco39792, w_eco39793, w_eco39794, w_eco39795, w_eco39796, w_eco39797, w_eco39798, w_eco39799, w_eco39800, w_eco39801, w_eco39802, w_eco39803, w_eco39804, w_eco39805, w_eco39806, w_eco39807, w_eco39808, w_eco39809, w_eco39810, w_eco39811, w_eco39812, w_eco39813, w_eco39814, w_eco39815, w_eco39816, w_eco39817, w_eco39818, w_eco39819, w_eco39820, w_eco39821, w_eco39822, w_eco39823, w_eco39824, w_eco39825, w_eco39826, w_eco39827, w_eco39828, w_eco39829, w_eco39830, w_eco39831, w_eco39832, w_eco39833, w_eco39834, w_eco39835, w_eco39836, w_eco39837, w_eco39838, w_eco39839, w_eco39840, w_eco39841, w_eco39842, w_eco39843, w_eco39844, w_eco39845, w_eco39846, w_eco39847, w_eco39848, w_eco39849, w_eco39850, w_eco39851, w_eco39852, w_eco39853, w_eco39854, w_eco39855, w_eco39856, w_eco39857, w_eco39858, w_eco39859, w_eco39860, w_eco39861, w_eco39862, w_eco39863, w_eco39864, w_eco39865, w_eco39866, w_eco39867, w_eco39868, w_eco39869, w_eco39870, w_eco39871, w_eco39872, w_eco39873, w_eco39874, w_eco39875, w_eco39876, w_eco39877, w_eco39878, w_eco39879, w_eco39880, w_eco39881, w_eco39882, w_eco39883, w_eco39884, w_eco39885, w_eco39886, w_eco39887, w_eco39888, w_eco39889, w_eco39890, w_eco39891, w_eco39892, w_eco39893, w_eco39894, w_eco39895, w_eco39896, w_eco39897, w_eco39898, w_eco39899, w_eco39900, w_eco39901, w_eco39902, w_eco39903, w_eco39904, w_eco39905, w_eco39906, w_eco39907, w_eco39908, w_eco39909, w_eco39910, w_eco39911, w_eco39912, w_eco39913, w_eco39914, w_eco39915, w_eco39916, w_eco39917, w_eco39918, w_eco39919, w_eco39920, w_eco39921, w_eco39922, w_eco39923, w_eco39924, w_eco39925, w_eco39926, w_eco39927, w_eco39928, w_eco39929, w_eco39930, w_eco39931, w_eco39932, w_eco39933, w_eco39934, w_eco39935, w_eco39936, w_eco39937, w_eco39938, w_eco39939, w_eco39940, w_eco39941, w_eco39942, w_eco39943, w_eco39944, w_eco39945, w_eco39946, w_eco39947, w_eco39948, w_eco39949, w_eco39950, w_eco39951, w_eco39952, w_eco39953, w_eco39954, w_eco39955, w_eco39956, w_eco39957, w_eco39958, w_eco39959, w_eco39960, w_eco39961, w_eco39962, w_eco39963, w_eco39964, w_eco39965, w_eco39966, w_eco39967, w_eco39968, w_eco39969, w_eco39970, w_eco39971, w_eco39972, w_eco39973, w_eco39974, w_eco39975, w_eco39976, w_eco39977, w_eco39978, w_eco39979, w_eco39980, w_eco39981, w_eco39982, w_eco39983, w_eco39984, w_eco39985, w_eco39986, w_eco39987, w_eco39988, w_eco39989, w_eco39990, w_eco39991, w_eco39992, w_eco39993, w_eco39994, w_eco39995, w_eco39996, w_eco39997, w_eco39998, w_eco39999, w_eco40000, w_eco40001, w_eco40002, w_eco40003, w_eco40004, w_eco40005, w_eco40006, w_eco40007, w_eco40008, w_eco40009, w_eco40010, w_eco40011, w_eco40012, w_eco40013, w_eco40014, w_eco40015, w_eco40016, w_eco40017, w_eco40018, w_eco40019, w_eco40020, w_eco40021, w_eco40022, w_eco40023, w_eco40024, w_eco40025, w_eco40026, w_eco40027, w_eco40028, w_eco40029, w_eco40030, w_eco40031, w_eco40032, w_eco40033, w_eco40034, w_eco40035, w_eco40036, w_eco40037, w_eco40038, w_eco40039, w_eco40040, w_eco40041, w_eco40042, w_eco40043, w_eco40044, w_eco40045, w_eco40046, w_eco40047, w_eco40048, w_eco40049, w_eco40050, w_eco40051, w_eco40052, w_eco40053, w_eco40054, w_eco40055, w_eco40056, w_eco40057, w_eco40058, w_eco40059, w_eco40060, w_eco40061, w_eco40062, w_eco40063, w_eco40064, w_eco40065, w_eco40066, w_eco40067, w_eco40068, w_eco40069, w_eco40070, w_eco40071, w_eco40072, w_eco40073, w_eco40074, w_eco40075, w_eco40076, w_eco40077, w_eco40078, w_eco40079, w_eco40080, w_eco40081, w_eco40082, w_eco40083, w_eco40084, w_eco40085, w_eco40086, w_eco40087, w_eco40088, w_eco40089, w_eco40090, w_eco40091, w_eco40092, w_eco40093, w_eco40094, w_eco40095, w_eco40096, w_eco40097, w_eco40098, w_eco40099, w_eco40100, w_eco40101, w_eco40102, w_eco40103, w_eco40104, w_eco40105, w_eco40106, w_eco40107, w_eco40108, w_eco40109, w_eco40110, w_eco40111, w_eco40112, w_eco40113, w_eco40114, w_eco40115, w_eco40116, w_eco40117, w_eco40118, w_eco40119, w_eco40120, w_eco40121, w_eco40122, w_eco40123, w_eco40124, w_eco40125, w_eco40126, w_eco40127, w_eco40128, w_eco40129, w_eco40130, w_eco40131, w_eco40132, w_eco40133, w_eco40134, w_eco40135, w_eco40136, w_eco40137, w_eco40138, w_eco40139, w_eco40140, w_eco40141, w_eco40142, w_eco40143, w_eco40144, w_eco40145, w_eco40146, w_eco40147, w_eco40148, w_eco40149, w_eco40150, w_eco40151, w_eco40152, w_eco40153, w_eco40154, w_eco40155, w_eco40156, w_eco40157, w_eco40158, w_eco40159, w_eco40160, w_eco40161, w_eco40162, w_eco40163, w_eco40164, w_eco40165, w_eco40166, w_eco40167, w_eco40168, w_eco40169, w_eco40170, w_eco40171, w_eco40172, w_eco40173, w_eco40174, w_eco40175, w_eco40176, w_eco40177, w_eco40178, w_eco40179, w_eco40180, w_eco40181, w_eco40182, w_eco40183, w_eco40184, w_eco40185, w_eco40186, w_eco40187, w_eco40188, w_eco40189, w_eco40190, w_eco40191, w_eco40192, w_eco40193, w_eco40194, w_eco40195, w_eco40196, w_eco40197, w_eco40198, w_eco40199, w_eco40200, w_eco40201, w_eco40202, w_eco40203, w_eco40204, w_eco40205, w_eco40206, w_eco40207, w_eco40208, w_eco40209, w_eco40210, w_eco40211, w_eco40212, w_eco40213, w_eco40214, w_eco40215, w_eco40216, w_eco40217, w_eco40218, w_eco40219, w_eco40220, w_eco40221, w_eco40222, w_eco40223, w_eco40224, w_eco40225, w_eco40226, w_eco40227, w_eco40228, w_eco40229, w_eco40230, w_eco40231, w_eco40232, w_eco40233, w_eco40234, w_eco40235, w_eco40236, w_eco40237, w_eco40238, w_eco40239, w_eco40240, w_eco40241, w_eco40242, w_eco40243, w_eco40244, w_eco40245, w_eco40246, w_eco40247, w_eco40248, w_eco40249, w_eco40250, w_eco40251, w_eco40252, w_eco40253, w_eco40254, w_eco40255, w_eco40256, w_eco40257, w_eco40258, w_eco40259, w_eco40260, w_eco40261, w_eco40262, w_eco40263, w_eco40264, w_eco40265, w_eco40266, w_eco40267, w_eco40268, w_eco40269, w_eco40270, w_eco40271, w_eco40272, w_eco40273, w_eco40274, w_eco40275, w_eco40276, w_eco40277, w_eco40278, w_eco40279, w_eco40280, w_eco40281, w_eco40282, w_eco40283, w_eco40284, w_eco40285, w_eco40286, w_eco40287, w_eco40288, w_eco40289, w_eco40290, w_eco40291, w_eco40292, w_eco40293, w_eco40294, w_eco40295, w_eco40296, w_eco40297, w_eco40298, w_eco40299, w_eco40300, w_eco40301, w_eco40302, w_eco40303, w_eco40304, w_eco40305, w_eco40306, w_eco40307, w_eco40308, w_eco40309, w_eco40310, w_eco40311, w_eco40312, w_eco40313, w_eco40314, w_eco40315, w_eco40316, w_eco40317, w_eco40318, w_eco40319, w_eco40320, w_eco40321, w_eco40322, w_eco40323, w_eco40324, w_eco40325, w_eco40326, w_eco40327, w_eco40328, w_eco40329, w_eco40330, w_eco40331, w_eco40332, w_eco40333, w_eco40334, w_eco40335, w_eco40336, w_eco40337, w_eco40338, w_eco40339, w_eco40340, w_eco40341, w_eco40342, w_eco40343, w_eco40344, w_eco40345, w_eco40346, w_eco40347, w_eco40348, w_eco40349, w_eco40350, w_eco40351, w_eco40352, w_eco40353, w_eco40354, w_eco40355, w_eco40356, w_eco40357, w_eco40358, w_eco40359, w_eco40360, w_eco40361, w_eco40362, w_eco40363, w_eco40364, w_eco40365, w_eco40366, w_eco40367, w_eco40368, w_eco40369, w_eco40370, w_eco40371, w_eco40372, w_eco40373, w_eco40374, w_eco40375, w_eco40376, w_eco40377, w_eco40378, w_eco40379, w_eco40380, w_eco40381, w_eco40382, w_eco40383, w_eco40384, w_eco40385, w_eco40386, w_eco40387, w_eco40388, w_eco40389, w_eco40390, w_eco40391, w_eco40392, w_eco40393, w_eco40394, w_eco40395, w_eco40396, w_eco40397, w_eco40398, w_eco40399, w_eco40400, w_eco40401, w_eco40402, w_eco40403, w_eco40404, w_eco40405, w_eco40406, w_eco40407, w_eco40408, w_eco40409, w_eco40410, w_eco40411, w_eco40412, w_eco40413, w_eco40414, w_eco40415, w_eco40416, w_eco40417, w_eco40418, w_eco40419, w_eco40420, w_eco40421, w_eco40422, w_eco40423, w_eco40424, w_eco40425, w_eco40426, w_eco40427, w_eco40428, w_eco40429, w_eco40430, w_eco40431, w_eco40432, w_eco40433, w_eco40434, w_eco40435, w_eco40436, w_eco40437, w_eco40438, w_eco40439, w_eco40440, w_eco40441, w_eco40442, w_eco40443, w_eco40444, w_eco40445, w_eco40446, w_eco40447, w_eco40448, w_eco40449, w_eco40450, w_eco40451, w_eco40452, w_eco40453, w_eco40454, w_eco40455, w_eco40456, w_eco40457, w_eco40458, w_eco40459, w_eco40460, w_eco40461, w_eco40462, w_eco40463, w_eco40464, w_eco40465, w_eco40466, w_eco40467, w_eco40468, w_eco40469, w_eco40470, w_eco40471, w_eco40472, w_eco40473, w_eco40474, w_eco40475, w_eco40476, w_eco40477, w_eco40478, w_eco40479, w_eco40480, w_eco40481, w_eco40482, w_eco40483, w_eco40484, w_eco40485, w_eco40486, w_eco40487, w_eco40488, w_eco40489, w_eco40490, w_eco40491, w_eco40492, w_eco40493, w_eco40494, w_eco40495, w_eco40496, w_eco40497, w_eco40498, w_eco40499, w_eco40500, w_eco40501, w_eco40502, w_eco40503, w_eco40504, w_eco40505, w_eco40506, w_eco40507, w_eco40508, w_eco40509, w_eco40510, w_eco40511, w_eco40512, w_eco40513, w_eco40514, w_eco40515, w_eco40516, w_eco40517, w_eco40518, w_eco40519, w_eco40520, w_eco40521, w_eco40522, w_eco40523, w_eco40524, w_eco40525, w_eco40526, w_eco40527, w_eco40528, w_eco40529, w_eco40530, w_eco40531, w_eco40532, w_eco40533, w_eco40534, w_eco40535, w_eco40536, w_eco40537, w_eco40538, w_eco40539, w_eco40540, w_eco40541, w_eco40542, w_eco40543, w_eco40544, w_eco40545, w_eco40546, w_eco40547, w_eco40548, w_eco40549, w_eco40550, w_eco40551, w_eco40552, w_eco40553, w_eco40554, w_eco40555, w_eco40556, w_eco40557, w_eco40558, w_eco40559, w_eco40560, w_eco40561, w_eco40562, w_eco40563, w_eco40564, w_eco40565, w_eco40566, w_eco40567, w_eco40568, w_eco40569, w_eco40570, w_eco40571, w_eco40572, w_eco40573, w_eco40574, w_eco40575, w_eco40576, w_eco40577, w_eco40578, w_eco40579, w_eco40580, w_eco40581, w_eco40582, w_eco40583, w_eco40584, w_eco40585, w_eco40586, w_eco40587, w_eco40588, w_eco40589, w_eco40590, w_eco40591, w_eco40592, w_eco40593, w_eco40594, w_eco40595, w_eco40596, w_eco40597, w_eco40598, w_eco40599, w_eco40600, w_eco40601, w_eco40602, w_eco40603, w_eco40604, w_eco40605, w_eco40606, w_eco40607, w_eco40608, w_eco40609, w_eco40610, w_eco40611, w_eco40612, w_eco40613, w_eco40614, w_eco40615, w_eco40616, w_eco40617, w_eco40618, w_eco40619, w_eco40620, w_eco40621, w_eco40622, w_eco40623, w_eco40624, w_eco40625, w_eco40626, w_eco40627, w_eco40628, w_eco40629, w_eco40630, w_eco40631, w_eco40632, w_eco40633, w_eco40634, w_eco40635, w_eco40636, w_eco40637, w_eco40638, w_eco40639, w_eco40640, w_eco40641, w_eco40642, w_eco40643, w_eco40644, w_eco40645, w_eco40646, w_eco40647, w_eco40648, w_eco40649, w_eco40650, w_eco40651, w_eco40652, w_eco40653, w_eco40654, w_eco40655, w_eco40656, w_eco40657, w_eco40658, w_eco40659, w_eco40660, w_eco40661, w_eco40662, w_eco40663, w_eco40664, w_eco40665, w_eco40666, w_eco40667, w_eco40668, w_eco40669, w_eco40670, w_eco40671, w_eco40672, w_eco40673, w_eco40674, w_eco40675, w_eco40676, w_eco40677, w_eco40678, w_eco40679, w_eco40680, w_eco40681, w_eco40682, w_eco40683, w_eco40684, w_eco40685, w_eco40686, w_eco40687, w_eco40688, w_eco40689, w_eco40690, w_eco40691, w_eco40692, w_eco40693, w_eco40694, w_eco40695, w_eco40696, w_eco40697, w_eco40698, w_eco40699, w_eco40700, w_eco40701, w_eco40702, w_eco40703, w_eco40704, w_eco40705, w_eco40706, w_eco40707, w_eco40708, w_eco40709, w_eco40710, w_eco40711, w_eco40712, w_eco40713, w_eco40714, w_eco40715, w_eco40716, w_eco40717, w_eco40718, w_eco40719, w_eco40720, w_eco40721, w_eco40722, w_eco40723, w_eco40724, w_eco40725, w_eco40726, w_eco40727, w_eco40728, w_eco40729, w_eco40730, w_eco40731, w_eco40732, w_eco40733, w_eco40734, w_eco40735, w_eco40736, w_eco40737, w_eco40738, w_eco40739, w_eco40740, w_eco40741, w_eco40742, w_eco40743, w_eco40744, w_eco40745, w_eco40746, w_eco40747, w_eco40748, w_eco40749, w_eco40750, w_eco40751, w_eco40752, w_eco40753, w_eco40754, w_eco40755, w_eco40756, w_eco40757, w_eco40758, w_eco40759, w_eco40760, w_eco40761, w_eco40762, w_eco40763, w_eco40764, w_eco40765, w_eco40766, w_eco40767, w_eco40768, w_eco40769, w_eco40770, w_eco40771, w_eco40772, w_eco40773, w_eco40774, w_eco40775, w_eco40776, w_eco40777, w_eco40778, w_eco40779, w_eco40780, w_eco40781, w_eco40782, w_eco40783, w_eco40784, w_eco40785, w_eco40786, w_eco40787, w_eco40788, w_eco40789, w_eco40790, w_eco40791, w_eco40792, w_eco40793, w_eco40794, w_eco40795, w_eco40796, w_eco40797, w_eco40798, w_eco40799, w_eco40800, w_eco40801, w_eco40802, w_eco40803, w_eco40804, w_eco40805, w_eco40806, w_eco40807, w_eco40808, w_eco40809, w_eco40810, w_eco40811, w_eco40812, w_eco40813, w_eco40814, w_eco40815, w_eco40816, w_eco40817, w_eco40818, w_eco40819, w_eco40820, w_eco40821, w_eco40822, w_eco40823, w_eco40824, w_eco40825, w_eco40826, w_eco40827, w_eco40828, w_eco40829, w_eco40830, w_eco40831, w_eco40832, w_eco40833, w_eco40834, w_eco40835, w_eco40836, w_eco40837, w_eco40838, w_eco40839, w_eco40840, w_eco40841, w_eco40842, w_eco40843, w_eco40844, w_eco40845, w_eco40846, w_eco40847, w_eco40848, w_eco40849, w_eco40850, w_eco40851, w_eco40852, w_eco40853, w_eco40854, w_eco40855, w_eco40856, w_eco40857, w_eco40858, w_eco40859, w_eco40860, w_eco40861, w_eco40862, w_eco40863, w_eco40864, w_eco40865, w_eco40866, w_eco40867, w_eco40868, w_eco40869, w_eco40870, w_eco40871, w_eco40872, w_eco40873, w_eco40874, w_eco40875, w_eco40876, w_eco40877, w_eco40878, w_eco40879, w_eco40880, w_eco40881, w_eco40882, w_eco40883, w_eco40884, w_eco40885, w_eco40886, w_eco40887, w_eco40888, w_eco40889, w_eco40890, w_eco40891, w_eco40892, w_eco40893, w_eco40894, w_eco40895, w_eco40896, w_eco40897, w_eco40898, w_eco40899, w_eco40900, w_eco40901, w_eco40902, w_eco40903, w_eco40904, w_eco40905, w_eco40906, w_eco40907, w_eco40908, w_eco40909, w_eco40910, w_eco40911, w_eco40912, w_eco40913, w_eco40914, w_eco40915, w_eco40916, w_eco40917, w_eco40918, w_eco40919, w_eco40920, w_eco40921, w_eco40922, w_eco40923, w_eco40924, w_eco40925, w_eco40926, w_eco40927, w_eco40928, w_eco40929, w_eco40930, w_eco40931, w_eco40932, w_eco40933, w_eco40934, w_eco40935, w_eco40936, w_eco40937, w_eco40938, w_eco40939, w_eco40940, w_eco40941, w_eco40942, w_eco40943, w_eco40944, w_eco40945, w_eco40946, w_eco40947, w_eco40948, w_eco40949, w_eco40950, w_eco40951, w_eco40952, w_eco40953, w_eco40954, w_eco40955, w_eco40956, w_eco40957, w_eco40958, w_eco40959, w_eco40960, w_eco40961, w_eco40962, w_eco40963, w_eco40964, w_eco40965, w_eco40966, w_eco40967, w_eco40968, w_eco40969, w_eco40970, w_eco40971, w_eco40972, w_eco40973, w_eco40974, w_eco40975, w_eco40976, w_eco40977, w_eco40978, w_eco40979, w_eco40980, w_eco40981, w_eco40982, w_eco40983, w_eco40984, w_eco40985, w_eco40986, w_eco40987, w_eco40988, w_eco40989, w_eco40990, w_eco40991, w_eco40992, w_eco40993, w_eco40994, w_eco40995, w_eco40996, w_eco40997, w_eco40998, w_eco40999, w_eco41000, w_eco41001, w_eco41002, w_eco41003, w_eco41004, w_eco41005, w_eco41006, w_eco41007, w_eco41008, w_eco41009, w_eco41010, w_eco41011, w_eco41012, w_eco41013, w_eco41014, w_eco41015, w_eco41016, w_eco41017, w_eco41018, w_eco41019, w_eco41020, w_eco41021, w_eco41022, w_eco41023, w_eco41024, w_eco41025, w_eco41026, w_eco41027, w_eco41028, w_eco41029, w_eco41030, w_eco41031, w_eco41032, w_eco41033, w_eco41034, w_eco41035, w_eco41036, w_eco41037, w_eco41038, w_eco41039, w_eco41040, w_eco41041, w_eco41042, w_eco41043, w_eco41044, w_eco41045, w_eco41046, w_eco41047, w_eco41048, w_eco41049, w_eco41050, w_eco41051, w_eco41052, w_eco41053, w_eco41054, w_eco41055, w_eco41056, w_eco41057, w_eco41058, w_eco41059, w_eco41060, w_eco41061, w_eco41062, w_eco41063, w_eco41064, w_eco41065, w_eco41066, w_eco41067, w_eco41068, w_eco41069, w_eco41070, w_eco41071, w_eco41072, w_eco41073, w_eco41074, w_eco41075, w_eco41076, w_eco41077, w_eco41078, w_eco41079, w_eco41080, w_eco41081, w_eco41082, w_eco41083, w_eco41084, w_eco41085, w_eco41086, w_eco41087, w_eco41088, w_eco41089, w_eco41090, w_eco41091, w_eco41092, w_eco41093, w_eco41094, w_eco41095, w_eco41096, w_eco41097, w_eco41098, w_eco41099, w_eco41100, w_eco41101, w_eco41102, w_eco41103, w_eco41104, w_eco41105, w_eco41106, w_eco41107, w_eco41108, w_eco41109, w_eco41110, w_eco41111, w_eco41112, w_eco41113, w_eco41114, w_eco41115, w_eco41116, w_eco41117, w_eco41118, w_eco41119, w_eco41120, w_eco41121, w_eco41122, w_eco41123, w_eco41124, w_eco41125, w_eco41126, w_eco41127, w_eco41128, w_eco41129, w_eco41130, w_eco41131, w_eco41132, w_eco41133, w_eco41134, w_eco41135, w_eco41136, w_eco41137, w_eco41138, w_eco41139, w_eco41140, w_eco41141, w_eco41142, w_eco41143, w_eco41144, w_eco41145, w_eco41146, w_eco41147, w_eco41148, w_eco41149, w_eco41150, w_eco41151, w_eco41152, w_eco41153, w_eco41154, w_eco41155, w_eco41156, w_eco41157, w_eco41158, w_eco41159, w_eco41160, w_eco41161, w_eco41162, w_eco41163, w_eco41164, w_eco41165, w_eco41166, w_eco41167, w_eco41168, w_eco41169, w_eco41170, w_eco41171, w_eco41172, w_eco41173, w_eco41174, w_eco41175, w_eco41176, w_eco41177, w_eco41178, w_eco41179, w_eco41180, w_eco41181, w_eco41182, w_eco41183, w_eco41184, w_eco41185, w_eco41186, w_eco41187, w_eco41188, w_eco41189, w_eco41190, w_eco41191, w_eco41192, w_eco41193, w_eco41194, w_eco41195, w_eco41196, w_eco41197, w_eco41198, w_eco41199, w_eco41200, w_eco41201, w_eco41202, w_eco41203, w_eco41204, w_eco41205, w_eco41206, w_eco41207, w_eco41208, w_eco41209, w_eco41210, w_eco41211, w_eco41212, w_eco41213, w_eco41214, w_eco41215, w_eco41216, w_eco41217, w_eco41218, w_eco41219, w_eco41220, w_eco41221, w_eco41222, w_eco41223, w_eco41224, w_eco41225, w_eco41226, w_eco41227, w_eco41228, w_eco41229, w_eco41230, w_eco41231, w_eco41232, w_eco41233, w_eco41234, w_eco41235, w_eco41236, w_eco41237, w_eco41238, w_eco41239, w_eco41240, w_eco41241, w_eco41242, w_eco41243, w_eco41244, w_eco41245, w_eco41246, w_eco41247, w_eco41248, w_eco41249, w_eco41250, w_eco41251, w_eco41252, w_eco41253, w_eco41254, w_eco41255, w_eco41256, w_eco41257, w_eco41258, w_eco41259, w_eco41260, w_eco41261, w_eco41262, w_eco41263, w_eco41264, w_eco41265, w_eco41266, w_eco41267, w_eco41268, w_eco41269, w_eco41270, w_eco41271, w_eco41272, w_eco41273, w_eco41274, w_eco41275, w_eco41276, w_eco41277, w_eco41278, w_eco41279, w_eco41280, w_eco41281, w_eco41282, w_eco41283, w_eco41284, w_eco41285, w_eco41286, w_eco41287, w_eco41288, w_eco41289, w_eco41290, w_eco41291, w_eco41292, w_eco41293, w_eco41294, w_eco41295, w_eco41296, w_eco41297, w_eco41298, w_eco41299, w_eco41300, w_eco41301, w_eco41302, w_eco41303, w_eco41304, w_eco41305, w_eco41306, w_eco41307, w_eco41308, w_eco41309, w_eco41310, w_eco41311, w_eco41312, w_eco41313, w_eco41314, w_eco41315, w_eco41316, w_eco41317, w_eco41318, w_eco41319, w_eco41320, w_eco41321, w_eco41322, w_eco41323, w_eco41324, w_eco41325, w_eco41326, w_eco41327, w_eco41328, w_eco41329, w_eco41330, w_eco41331, w_eco41332, w_eco41333, w_eco41334, w_eco41335, w_eco41336, w_eco41337, w_eco41338, w_eco41339, w_eco41340, w_eco41341, w_eco41342, w_eco41343, w_eco41344, w_eco41345, w_eco41346, w_eco41347, w_eco41348, w_eco41349, w_eco41350, w_eco41351, w_eco41352, w_eco41353, w_eco41354, w_eco41355, w_eco41356, w_eco41357, w_eco41358, w_eco41359, w_eco41360, w_eco41361, w_eco41362, w_eco41363, w_eco41364, w_eco41365, w_eco41366, w_eco41367, w_eco41368, w_eco41369, w_eco41370, w_eco41371, w_eco41372, w_eco41373, w_eco41374, w_eco41375, w_eco41376, w_eco41377, w_eco41378, w_eco41379, w_eco41380, w_eco41381, w_eco41382, w_eco41383, w_eco41384, w_eco41385, w_eco41386, w_eco41387, w_eco41388, w_eco41389, w_eco41390, w_eco41391, w_eco41392, w_eco41393, w_eco41394, w_eco41395, w_eco41396, w_eco41397, w_eco41398, w_eco41399, w_eco41400, w_eco41401, w_eco41402, w_eco41403, w_eco41404, w_eco41405, w_eco41406, w_eco41407, w_eco41408, w_eco41409, w_eco41410, w_eco41411, w_eco41412, w_eco41413, w_eco41414, w_eco41415, w_eco41416, w_eco41417, w_eco41418, w_eco41419, w_eco41420, w_eco41421, w_eco41422, w_eco41423, w_eco41424, w_eco41425, w_eco41426, w_eco41427, w_eco41428, w_eco41429, w_eco41430, w_eco41431, w_eco41432, w_eco41433, w_eco41434, w_eco41435, w_eco41436, w_eco41437, w_eco41438, w_eco41439, w_eco41440, w_eco41441, w_eco41442, w_eco41443, w_eco41444, w_eco41445, w_eco41446, w_eco41447, w_eco41448, w_eco41449, w_eco41450, w_eco41451, w_eco41452, w_eco41453, w_eco41454, w_eco41455, w_eco41456, w_eco41457, w_eco41458, w_eco41459, w_eco41460, w_eco41461, w_eco41462, w_eco41463, w_eco41464, w_eco41465, w_eco41466, w_eco41467, w_eco41468, w_eco41469, w_eco41470, w_eco41471, w_eco41472, w_eco41473, w_eco41474, w_eco41475, w_eco41476, w_eco41477, w_eco41478, w_eco41479, w_eco41480, w_eco41481, w_eco41482, w_eco41483, w_eco41484, w_eco41485, w_eco41486, w_eco41487, w_eco41488, w_eco41489, w_eco41490, w_eco41491, w_eco41492, w_eco41493, w_eco41494, w_eco41495, w_eco41496, w_eco41497, w_eco41498, w_eco41499, w_eco41500, w_eco41501, w_eco41502, w_eco41503, w_eco41504, w_eco41505, w_eco41506, w_eco41507, w_eco41508, w_eco41509, w_eco41510, w_eco41511, w_eco41512, w_eco41513, w_eco41514, w_eco41515, w_eco41516, w_eco41517, w_eco41518, w_eco41519, w_eco41520, w_eco41521, w_eco41522, w_eco41523, w_eco41524, w_eco41525, w_eco41526, w_eco41527, w_eco41528, w_eco41529, w_eco41530, w_eco41531, w_eco41532, w_eco41533, w_eco41534, w_eco41535, w_eco41536, w_eco41537, w_eco41538, w_eco41539, w_eco41540, w_eco41541, w_eco41542, w_eco41543, w_eco41544, w_eco41545, w_eco41546, w_eco41547, w_eco41548, w_eco41549, w_eco41550, w_eco41551, w_eco41552, w_eco41553, w_eco41554, w_eco41555, w_eco41556, w_eco41557, w_eco41558, w_eco41559, w_eco41560, w_eco41561, w_eco41562, w_eco41563, w_eco41564, w_eco41565, w_eco41566, w_eco41567, w_eco41568, w_eco41569, w_eco41570, w_eco41571, w_eco41572, w_eco41573, w_eco41574, w_eco41575, w_eco41576, w_eco41577, w_eco41578, w_eco41579, w_eco41580, w_eco41581, w_eco41582, w_eco41583, w_eco41584, w_eco41585, w_eco41586, w_eco41587, w_eco41588, w_eco41589, w_eco41590, w_eco41591, w_eco41592, w_eco41593, w_eco41594, w_eco41595, w_eco41596, w_eco41597, w_eco41598, w_eco41599, w_eco41600, w_eco41601, w_eco41602, w_eco41603, w_eco41604, w_eco41605, w_eco41606, w_eco41607, w_eco41608, w_eco41609, w_eco41610, w_eco41611, w_eco41612, w_eco41613, w_eco41614, w_eco41615, w_eco41616, w_eco41617, w_eco41618, w_eco41619, w_eco41620, w_eco41621, w_eco41622, w_eco41623, w_eco41624, w_eco41625, w_eco41626, w_eco41627, w_eco41628, w_eco41629, w_eco41630, w_eco41631, w_eco41632, w_eco41633, w_eco41634, w_eco41635, w_eco41636, w_eco41637, w_eco41638, w_eco41639, w_eco41640, w_eco41641, w_eco41642, w_eco41643, w_eco41644, w_eco41645, w_eco41646, w_eco41647, w_eco41648, w_eco41649, w_eco41650, w_eco41651, w_eco41652, w_eco41653, w_eco41654, w_eco41655, w_eco41656, w_eco41657, w_eco41658, w_eco41659, w_eco41660, w_eco41661, w_eco41662, w_eco41663, w_eco41664, w_eco41665, w_eco41666, w_eco41667, w_eco41668, w_eco41669, w_eco41670, w_eco41671, w_eco41672, w_eco41673, w_eco41674, w_eco41675, w_eco41676, w_eco41677, w_eco41678, w_eco41679, w_eco41680, w_eco41681, w_eco41682, w_eco41683, w_eco41684, w_eco41685, w_eco41686, w_eco41687, w_eco41688, w_eco41689, w_eco41690, w_eco41691, w_eco41692, w_eco41693, w_eco41694, w_eco41695, w_eco41696, w_eco41697, w_eco41698, w_eco41699, w_eco41700, w_eco41701, w_eco41702, w_eco41703, w_eco41704, w_eco41705, w_eco41706, w_eco41707, w_eco41708, w_eco41709, w_eco41710, w_eco41711, w_eco41712, w_eco41713, w_eco41714, w_eco41715, w_eco41716, w_eco41717, w_eco41718, w_eco41719, w_eco41720, w_eco41721, w_eco41722, w_eco41723, w_eco41724, w_eco41725, w_eco41726, w_eco41727, w_eco41728, w_eco41729, w_eco41730, w_eco41731, w_eco41732, w_eco41733, w_eco41734, w_eco41735, w_eco41736, w_eco41737, w_eco41738, w_eco41739, w_eco41740, w_eco41741, w_eco41742, w_eco41743, w_eco41744, w_eco41745, w_eco41746, w_eco41747, w_eco41748, w_eco41749, w_eco41750, w_eco41751, w_eco41752, w_eco41753, w_eco41754, w_eco41755, w_eco41756, w_eco41757, w_eco41758, w_eco41759, w_eco41760, w_eco41761, w_eco41762, w_eco41763, w_eco41764, w_eco41765, w_eco41766, w_eco41767, w_eco41768, w_eco41769, w_eco41770, w_eco41771, w_eco41772, w_eco41773, w_eco41774, w_eco41775, w_eco41776, w_eco41777, w_eco41778, w_eco41779, w_eco41780, w_eco41781, w_eco41782, w_eco41783, w_eco41784, w_eco41785, w_eco41786, w_eco41787, w_eco41788, w_eco41789, w_eco41790, w_eco41791, w_eco41792, w_eco41793, w_eco41794, w_eco41795, w_eco41796, w_eco41797, w_eco41798, w_eco41799, w_eco41800, w_eco41801, w_eco41802, w_eco41803, w_eco41804, w_eco41805, w_eco41806, w_eco41807, w_eco41808, w_eco41809, w_eco41810, w_eco41811, w_eco41812, w_eco41813, w_eco41814, w_eco41815, w_eco41816, w_eco41817, w_eco41818, w_eco41819, w_eco41820, w_eco41821, w_eco41822, w_eco41823, w_eco41824, w_eco41825, w_eco41826, w_eco41827, w_eco41828, w_eco41829, w_eco41830, w_eco41831, w_eco41832, w_eco41833, w_eco41834, w_eco41835, w_eco41836, w_eco41837, w_eco41838, w_eco41839, w_eco41840, w_eco41841, w_eco41842, w_eco41843, w_eco41844, w_eco41845, w_eco41846, w_eco41847, w_eco41848, w_eco41849, w_eco41850, w_eco41851, w_eco41852, w_eco41853, w_eco41854, w_eco41855, w_eco41856, w_eco41857, w_eco41858, w_eco41859, w_eco41860, w_eco41861, w_eco41862, w_eco41863, w_eco41864, w_eco41865, w_eco41866, w_eco41867, w_eco41868, w_eco41869, w_eco41870, w_eco41871, w_eco41872, w_eco41873, w_eco41874, w_eco41875, w_eco41876, w_eco41877, w_eco41878, w_eco41879, w_eco41880, w_eco41881, w_eco41882, w_eco41883, w_eco41884, w_eco41885, w_eco41886, w_eco41887, w_eco41888, w_eco41889, w_eco41890, w_eco41891, w_eco41892, w_eco41893, w_eco41894, w_eco41895, w_eco41896, w_eco41897, w_eco41898, w_eco41899, w_eco41900, w_eco41901, w_eco41902, w_eco41903, w_eco41904, w_eco41905, w_eco41906, w_eco41907, w_eco41908, w_eco41909, w_eco41910, w_eco41911, w_eco41912, w_eco41913, w_eco41914, w_eco41915, w_eco41916, w_eco41917, w_eco41918, w_eco41919, w_eco41920, w_eco41921, w_eco41922, w_eco41923, w_eco41924, w_eco41925, w_eco41926, w_eco41927, w_eco41928, w_eco41929, w_eco41930, w_eco41931, w_eco41932, w_eco41933, w_eco41934, w_eco41935, w_eco41936, w_eco41937, w_eco41938, w_eco41939, w_eco41940, w_eco41941, w_eco41942, w_eco41943, w_eco41944, w_eco41945, w_eco41946, w_eco41947, w_eco41948, w_eco41949, w_eco41950, w_eco41951, w_eco41952, w_eco41953, w_eco41954, w_eco41955, w_eco41956, w_eco41957, w_eco41958, w_eco41959, w_eco41960, w_eco41961, w_eco41962, w_eco41963, w_eco41964, w_eco41965, w_eco41966, w_eco41967, w_eco41968, w_eco41969, w_eco41970, w_eco41971, w_eco41972, w_eco41973, w_eco41974, w_eco41975, w_eco41976, w_eco41977, w_eco41978, w_eco41979, w_eco41980, w_eco41981, w_eco41982, w_eco41983, w_eco41984, w_eco41985, w_eco41986, w_eco41987, w_eco41988, w_eco41989, w_eco41990, w_eco41991, w_eco41992, w_eco41993, w_eco41994, w_eco41995, w_eco41996, w_eco41997, w_eco41998, w_eco41999, w_eco42000, w_eco42001, w_eco42002, w_eco42003, w_eco42004, w_eco42005, w_eco42006, w_eco42007, w_eco42008, w_eco42009, w_eco42010, w_eco42011, w_eco42012, w_eco42013, w_eco42014, w_eco42015, w_eco42016, w_eco42017, w_eco42018, w_eco42019, w_eco42020, w_eco42021, w_eco42022, w_eco42023, w_eco42024, w_eco42025, w_eco42026, w_eco42027, w_eco42028, w_eco42029, w_eco42030, w_eco42031, w_eco42032, w_eco42033, w_eco42034, w_eco42035, w_eco42036, w_eco42037, w_eco42038, w_eco42039, w_eco42040, w_eco42041, w_eco42042, w_eco42043, w_eco42044, w_eco42045, w_eco42046, w_eco42047, w_eco42048, w_eco42049, w_eco42050, w_eco42051, w_eco42052, w_eco42053, w_eco42054, w_eco42055, w_eco42056, w_eco42057, w_eco42058, w_eco42059, w_eco42060, w_eco42061, w_eco42062, w_eco42063, w_eco42064, w_eco42065, w_eco42066, w_eco42067, w_eco42068, w_eco42069, w_eco42070, w_eco42071, w_eco42072, w_eco42073, w_eco42074, w_eco42075, w_eco42076, w_eco42077, w_eco42078, w_eco42079, w_eco42080, w_eco42081, w_eco42082, w_eco42083, w_eco42084, w_eco42085, w_eco42086, w_eco42087, w_eco42088, w_eco42089, w_eco42090, w_eco42091, w_eco42092, w_eco42093, w_eco42094, w_eco42095, w_eco42096, w_eco42097, w_eco42098, w_eco42099, w_eco42100, w_eco42101, w_eco42102, w_eco42103, w_eco42104, w_eco42105, w_eco42106, w_eco42107, w_eco42108, w_eco42109, w_eco42110, w_eco42111, w_eco42112, w_eco42113, w_eco42114, w_eco42115, w_eco42116, w_eco42117, w_eco42118, w_eco42119, w_eco42120, w_eco42121, w_eco42122, w_eco42123, w_eco42124, w_eco42125, w_eco42126, w_eco42127, w_eco42128, w_eco42129, w_eco42130, w_eco42131, w_eco42132, w_eco42133, w_eco42134, w_eco42135, w_eco42136, w_eco42137, w_eco42138, w_eco42139, w_eco42140, w_eco42141, w_eco42142, w_eco42143, w_eco42144, w_eco42145, w_eco42146, w_eco42147, w_eco42148, w_eco42149, w_eco42150, w_eco42151, w_eco42152, w_eco42153, w_eco42154, w_eco42155, w_eco42156, w_eco42157, w_eco42158, w_eco42159, w_eco42160, w_eco42161, w_eco42162, w_eco42163, w_eco42164, w_eco42165, w_eco42166, w_eco42167, w_eco42168, w_eco42169, w_eco42170, w_eco42171, w_eco42172, w_eco42173, w_eco42174, w_eco42175, w_eco42176, w_eco42177, w_eco42178, w_eco42179, w_eco42180, w_eco42181, w_eco42182, w_eco42183, w_eco42184, w_eco42185, w_eco42186, w_eco42187, w_eco42188, w_eco42189, w_eco42190, w_eco42191, w_eco42192, w_eco42193, w_eco42194, w_eco42195, w_eco42196, w_eco42197, w_eco42198, w_eco42199, w_eco42200, w_eco42201, w_eco42202, w_eco42203, w_eco42204, w_eco42205, w_eco42206, w_eco42207, w_eco42208, w_eco42209, w_eco42210, w_eco42211, w_eco42212, w_eco42213, w_eco42214, w_eco42215, w_eco42216, w_eco42217, w_eco42218, w_eco42219, w_eco42220, w_eco42221, w_eco42222, w_eco42223, w_eco42224, w_eco42225, w_eco42226, w_eco42227, w_eco42228, w_eco42229, w_eco42230, w_eco42231, w_eco42232, w_eco42233, w_eco42234, w_eco42235, w_eco42236, w_eco42237, w_eco42238, w_eco42239, w_eco42240, w_eco42241, w_eco42242, w_eco42243, w_eco42244, w_eco42245, w_eco42246, w_eco42247, w_eco42248, w_eco42249, w_eco42250, w_eco42251, w_eco42252, w_eco42253, w_eco42254, w_eco42255, w_eco42256, w_eco42257, w_eco42258, w_eco42259, w_eco42260, w_eco42261, w_eco42262, w_eco42263, w_eco42264, w_eco42265, w_eco42266, w_eco42267, w_eco42268, w_eco42269, w_eco42270, w_eco42271, w_eco42272, w_eco42273, w_eco42274, w_eco42275, w_eco42276, w_eco42277, w_eco42278, w_eco42279, w_eco42280, w_eco42281, w_eco42282, w_eco42283, w_eco42284, w_eco42285, w_eco42286, w_eco42287, w_eco42288, w_eco42289, w_eco42290, w_eco42291, w_eco42292, w_eco42293, w_eco42294, w_eco42295, w_eco42296, w_eco42297, w_eco42298, w_eco42299, w_eco42300, w_eco42301, w_eco42302, w_eco42303, w_eco42304, w_eco42305, w_eco42306, w_eco42307, w_eco42308, w_eco42309, w_eco42310, w_eco42311, w_eco42312, w_eco42313, w_eco42314, w_eco42315, w_eco42316, w_eco42317, w_eco42318, w_eco42319, w_eco42320, w_eco42321, w_eco42322, w_eco42323, w_eco42324, w_eco42325, w_eco42326, w_eco42327, w_eco42328, w_eco42329, w_eco42330, w_eco42331, w_eco42332, w_eco42333, w_eco42334, w_eco42335, w_eco42336, w_eco42337, w_eco42338, w_eco42339, w_eco42340, w_eco42341, w_eco42342, w_eco42343, w_eco42344, w_eco42345, w_eco42346, w_eco42347, w_eco42348, w_eco42349, w_eco42350, w_eco42351, w_eco42352, w_eco42353, w_eco42354, w_eco42355, w_eco42356, w_eco42357, w_eco42358, w_eco42359, w_eco42360, w_eco42361, w_eco42362, w_eco42363, w_eco42364, w_eco42365, w_eco42366, w_eco42367, w_eco42368, w_eco42369, w_eco42370, w_eco42371, w_eco42372, w_eco42373, w_eco42374, w_eco42375, w_eco42376, w_eco42377, w_eco42378, w_eco42379, w_eco42380, w_eco42381, w_eco42382, w_eco42383, w_eco42384, w_eco42385, w_eco42386, w_eco42387, w_eco42388, w_eco42389, w_eco42390, w_eco42391, w_eco42392, w_eco42393, w_eco42394, w_eco42395, w_eco42396, w_eco42397, w_eco42398, w_eco42399, w_eco42400, w_eco42401, w_eco42402, w_eco42403, w_eco42404, w_eco42405, w_eco42406, w_eco42407, w_eco42408, w_eco42409, w_eco42410, w_eco42411, w_eco42412, w_eco42413, w_eco42414, w_eco42415, w_eco42416, w_eco42417, w_eco42418, w_eco42419, w_eco42420, w_eco42421, w_eco42422, w_eco42423, w_eco42424, w_eco42425, w_eco42426, w_eco42427, w_eco42428, w_eco42429, w_eco42430, w_eco42431, w_eco42432, w_eco42433, w_eco42434, w_eco42435, w_eco42436, w_eco42437, w_eco42438, w_eco42439, w_eco42440, w_eco42441, w_eco42442, w_eco42443, w_eco42444, w_eco42445, w_eco42446, w_eco42447, w_eco42448, w_eco42449, w_eco42450, w_eco42451, w_eco42452, w_eco42453, w_eco42454, w_eco42455, w_eco42456, w_eco42457, w_eco42458, w_eco42459, w_eco42460, w_eco42461, w_eco42462, w_eco42463, w_eco42464, w_eco42465, w_eco42466, w_eco42467, w_eco42468, w_eco42469, w_eco42470, w_eco42471, w_eco42472, w_eco42473, w_eco42474, w_eco42475, w_eco42476, w_eco42477, w_eco42478, w_eco42479, w_eco42480, w_eco42481, w_eco42482, w_eco42483, w_eco42484, w_eco42485, w_eco42486, w_eco42487, w_eco42488, w_eco42489, w_eco42490, w_eco42491, w_eco42492, w_eco42493, w_eco42494, w_eco42495, w_eco42496, w_eco42497, w_eco42498, w_eco42499, w_eco42500, w_eco42501, w_eco42502, w_eco42503, w_eco42504, w_eco42505, w_eco42506, w_eco42507, w_eco42508, w_eco42509, w_eco42510, w_eco42511, w_eco42512, w_eco42513, w_eco42514, w_eco42515, w_eco42516, w_eco42517, w_eco42518, w_eco42519, w_eco42520, w_eco42521, w_eco42522, w_eco42523, w_eco42524, w_eco42525, w_eco42526, w_eco42527, w_eco42528, w_eco42529, w_eco42530, w_eco42531, w_eco42532, w_eco42533, w_eco42534, w_eco42535, w_eco42536, w_eco42537, w_eco42538, w_eco42539, w_eco42540, w_eco42541, w_eco42542, w_eco42543, w_eco42544, w_eco42545, w_eco42546, w_eco42547, w_eco42548, w_eco42549, w_eco42550, w_eco42551, w_eco42552, w_eco42553, w_eco42554, w_eco42555, w_eco42556, w_eco42557, w_eco42558, w_eco42559, w_eco42560, w_eco42561, w_eco42562, w_eco42563, w_eco42564, w_eco42565, w_eco42566, w_eco42567, w_eco42568, w_eco42569, w_eco42570, w_eco42571, w_eco42572, w_eco42573, w_eco42574, w_eco42575, w_eco42576, w_eco42577, w_eco42578, w_eco42579, w_eco42580, w_eco42581, w_eco42582, w_eco42583, w_eco42584, w_eco42585, w_eco42586, w_eco42587, w_eco42588, w_eco42589, w_eco42590, w_eco42591, w_eco42592, w_eco42593, w_eco42594, w_eco42595, w_eco42596, w_eco42597, w_eco42598, w_eco42599, w_eco42600, w_eco42601, w_eco42602, w_eco42603, w_eco42604, w_eco42605, w_eco42606, w_eco42607, w_eco42608, w_eco42609, w_eco42610, w_eco42611, w_eco42612, w_eco42613, w_eco42614, w_eco42615, w_eco42616, w_eco42617, w_eco42618, w_eco42619, w_eco42620, w_eco42621, w_eco42622, w_eco42623, w_eco42624, w_eco42625, w_eco42626, w_eco42627, w_eco42628, w_eco42629, w_eco42630, w_eco42631, w_eco42632, w_eco42633, w_eco42634, w_eco42635, w_eco42636, w_eco42637, w_eco42638, w_eco42639, w_eco42640, w_eco42641, w_eco42642, w_eco42643, w_eco42644, w_eco42645, w_eco42646, w_eco42647, w_eco42648, w_eco42649, w_eco42650, w_eco42651, w_eco42652, w_eco42653, w_eco42654, w_eco42655, w_eco42656, w_eco42657, w_eco42658, w_eco42659, w_eco42660, w_eco42661, w_eco42662, w_eco42663, w_eco42664, w_eco42665, w_eco42666, w_eco42667, w_eco42668, w_eco42669, w_eco42670, w_eco42671, w_eco42672, w_eco42673, w_eco42674, w_eco42675, w_eco42676, w_eco42677, w_eco42678, w_eco42679, w_eco42680, w_eco42681, w_eco42682, w_eco42683, w_eco42684, w_eco42685, w_eco42686, w_eco42687, w_eco42688, w_eco42689, w_eco42690, w_eco42691, w_eco42692, w_eco42693, w_eco42694, w_eco42695, w_eco42696, w_eco42697, w_eco42698, w_eco42699, w_eco42700, w_eco42701, w_eco42702, w_eco42703, w_eco42704, w_eco42705, w_eco42706, w_eco42707, w_eco42708, w_eco42709, w_eco42710, w_eco42711, w_eco42712, w_eco42713, w_eco42714, w_eco42715, w_eco42716, w_eco42717, w_eco42718, w_eco42719, w_eco42720, w_eco42721, w_eco42722, w_eco42723, w_eco42724, w_eco42725, w_eco42726, w_eco42727, w_eco42728, w_eco42729, w_eco42730, w_eco42731, w_eco42732, w_eco42733, w_eco42734, w_eco42735, w_eco42736, w_eco42737, w_eco42738, w_eco42739, w_eco42740, w_eco42741, w_eco42742, w_eco42743, w_eco42744, w_eco42745, w_eco42746, w_eco42747, w_eco42748, w_eco42749, w_eco42750, w_eco42751, w_eco42752, w_eco42753, w_eco42754, w_eco42755, w_eco42756, w_eco42757, w_eco42758, w_eco42759, w_eco42760, w_eco42761, w_eco42762, w_eco42763, w_eco42764, w_eco42765, w_eco42766, w_eco42767, w_eco42768, w_eco42769, w_eco42770, w_eco42771, w_eco42772, w_eco42773, w_eco42774, w_eco42775, w_eco42776, w_eco42777, w_eco42778, w_eco42779, w_eco42780, w_eco42781, w_eco42782, w_eco42783, w_eco42784, w_eco42785, w_eco42786, w_eco42787, w_eco42788, w_eco42789, w_eco42790, w_eco42791, w_eco42792, w_eco42793, w_eco42794, w_eco42795, w_eco42796, w_eco42797, w_eco42798, w_eco42799, w_eco42800, w_eco42801, w_eco42802, w_eco42803, w_eco42804, w_eco42805, w_eco42806, w_eco42807, w_eco42808, w_eco42809, w_eco42810, w_eco42811, w_eco42812, w_eco42813, w_eco42814, w_eco42815, w_eco42816, w_eco42817, w_eco42818, w_eco42819, w_eco42820, w_eco42821, w_eco42822, w_eco42823, w_eco42824, w_eco42825, w_eco42826, w_eco42827, w_eco42828, w_eco42829, w_eco42830, w_eco42831, w_eco42832, w_eco42833, w_eco42834, w_eco42835, w_eco42836, w_eco42837, w_eco42838, w_eco42839, w_eco42840, w_eco42841, w_eco42842, w_eco42843, w_eco42844, w_eco42845, w_eco42846, w_eco42847, w_eco42848, w_eco42849, w_eco42850, w_eco42851, w_eco42852, w_eco42853, w_eco42854, w_eco42855, w_eco42856, w_eco42857, w_eco42858, w_eco42859, w_eco42860, w_eco42861, w_eco42862, w_eco42863, w_eco42864, w_eco42865, w_eco42866, w_eco42867, w_eco42868, w_eco42869, w_eco42870, w_eco42871, w_eco42872, w_eco42873, w_eco42874, w_eco42875, w_eco42876, w_eco42877, w_eco42878, w_eco42879, w_eco42880, w_eco42881, w_eco42882, w_eco42883, w_eco42884, w_eco42885, w_eco42886, w_eco42887, w_eco42888, w_eco42889, w_eco42890, w_eco42891, w_eco42892, w_eco42893, w_eco42894, w_eco42895, w_eco42896, w_eco42897, w_eco42898, w_eco42899, w_eco42900, w_eco42901, w_eco42902, w_eco42903, w_eco42904, w_eco42905, w_eco42906, w_eco42907, w_eco42908, w_eco42909, w_eco42910, w_eco42911, w_eco42912, w_eco42913, w_eco42914, w_eco42915, w_eco42916, w_eco42917, w_eco42918, w_eco42919, w_eco42920, w_eco42921, w_eco42922, w_eco42923, w_eco42924, w_eco42925, w_eco42926, w_eco42927, w_eco42928, w_eco42929, w_eco42930, w_eco42931, w_eco42932, w_eco42933, w_eco42934, w_eco42935, w_eco42936, w_eco42937, w_eco42938, w_eco42939, w_eco42940, w_eco42941, w_eco42942, w_eco42943, w_eco42944, w_eco42945, w_eco42946, w_eco42947, w_eco42948, w_eco42949, w_eco42950, w_eco42951, w_eco42952, w_eco42953, w_eco42954, w_eco42955, w_eco42956, w_eco42957, w_eco42958, w_eco42959, w_eco42960, w_eco42961, w_eco42962, w_eco42963, w_eco42964, w_eco42965, w_eco42966, w_eco42967, w_eco42968, w_eco42969, w_eco42970, w_eco42971, w_eco42972, w_eco42973, w_eco42974, w_eco42975, w_eco42976, w_eco42977, w_eco42978, w_eco42979, w_eco42980, w_eco42981, w_eco42982, w_eco42983, w_eco42984, w_eco42985, w_eco42986, w_eco42987, w_eco42988, w_eco42989, w_eco42990, w_eco42991, w_eco42992, w_eco42993, w_eco42994, w_eco42995, w_eco42996, w_eco42997, w_eco42998, w_eco42999, w_eco43000, w_eco43001, w_eco43002, w_eco43003, w_eco43004, w_eco43005, w_eco43006, w_eco43007, w_eco43008, w_eco43009, w_eco43010, w_eco43011, w_eco43012, w_eco43013, w_eco43014, w_eco43015, w_eco43016, w_eco43017, w_eco43018, w_eco43019, w_eco43020, w_eco43021, w_eco43022, w_eco43023, w_eco43024, w_eco43025, w_eco43026, w_eco43027, w_eco43028, w_eco43029, w_eco43030, w_eco43031, w_eco43032, w_eco43033, w_eco43034, w_eco43035, w_eco43036, w_eco43037, w_eco43038, w_eco43039, w_eco43040, w_eco43041, w_eco43042, w_eco43043, w_eco43044, w_eco43045, w_eco43046, w_eco43047, w_eco43048, w_eco43049, w_eco43050, w_eco43051, w_eco43052, w_eco43053, w_eco43054, w_eco43055, w_eco43056, w_eco43057, w_eco43058, w_eco43059, w_eco43060, w_eco43061, w_eco43062, w_eco43063, w_eco43064, w_eco43065, w_eco43066, w_eco43067, w_eco43068, w_eco43069, w_eco43070, w_eco43071, w_eco43072, w_eco43073, w_eco43074, w_eco43075, w_eco43076, w_eco43077, w_eco43078, w_eco43079, w_eco43080, w_eco43081, w_eco43082, w_eco43083, w_eco43084, w_eco43085, w_eco43086, w_eco43087, w_eco43088, w_eco43089, w_eco43090, w_eco43091, w_eco43092, w_eco43093, w_eco43094, w_eco43095, w_eco43096, w_eco43097, w_eco43098, w_eco43099, w_eco43100, w_eco43101, w_eco43102, w_eco43103, w_eco43104, w_eco43105, w_eco43106, w_eco43107, w_eco43108, w_eco43109, w_eco43110, w_eco43111, w_eco43112, w_eco43113, w_eco43114, w_eco43115, w_eco43116, w_eco43117, w_eco43118, w_eco43119, w_eco43120, w_eco43121, w_eco43122, w_eco43123, w_eco43124, w_eco43125, w_eco43126, w_eco43127, w_eco43128, w_eco43129, w_eco43130, w_eco43131, w_eco43132, w_eco43133, w_eco43134, w_eco43135, w_eco43136, w_eco43137, w_eco43138, w_eco43139, w_eco43140, w_eco43141, w_eco43142, w_eco43143, w_eco43144, w_eco43145, w_eco43146, w_eco43147, w_eco43148, w_eco43149, w_eco43150, w_eco43151, w_eco43152, w_eco43153, w_eco43154, w_eco43155, w_eco43156, w_eco43157, w_eco43158, w_eco43159, w_eco43160, w_eco43161, w_eco43162, w_eco43163, w_eco43164, w_eco43165, w_eco43166, w_eco43167, w_eco43168, w_eco43169, w_eco43170, w_eco43171, w_eco43172, w_eco43173, w_eco43174, w_eco43175, w_eco43176, w_eco43177, w_eco43178, w_eco43179, w_eco43180, w_eco43181, w_eco43182, w_eco43183, w_eco43184, w_eco43185, w_eco43186, w_eco43187, w_eco43188, w_eco43189, w_eco43190, w_eco43191, w_eco43192, w_eco43193, w_eco43194, w_eco43195, w_eco43196, w_eco43197, w_eco43198, w_eco43199, w_eco43200, w_eco43201, w_eco43202, w_eco43203, w_eco43204, w_eco43205, w_eco43206, w_eco43207, w_eco43208, w_eco43209, w_eco43210, w_eco43211, w_eco43212, w_eco43213, w_eco43214, w_eco43215, w_eco43216, w_eco43217, w_eco43218, w_eco43219, w_eco43220, w_eco43221, w_eco43222, w_eco43223, w_eco43224, w_eco43225, w_eco43226, w_eco43227, w_eco43228, w_eco43229, w_eco43230, w_eco43231, w_eco43232, w_eco43233, w_eco43234, w_eco43235, w_eco43236, w_eco43237, w_eco43238, w_eco43239, w_eco43240, w_eco43241, w_eco43242, w_eco43243, w_eco43244, w_eco43245, w_eco43246, w_eco43247, w_eco43248, w_eco43249, w_eco43250, w_eco43251, w_eco43252, w_eco43253, w_eco43254, w_eco43255, w_eco43256, w_eco43257, w_eco43258, w_eco43259, w_eco43260, w_eco43261, w_eco43262, w_eco43263, w_eco43264, w_eco43265, w_eco43266, w_eco43267, w_eco43268, w_eco43269, w_eco43270, w_eco43271, w_eco43272, w_eco43273, w_eco43274, w_eco43275, w_eco43276, w_eco43277, w_eco43278, w_eco43279, w_eco43280, w_eco43281, w_eco43282, w_eco43283, w_eco43284, w_eco43285, w_eco43286, w_eco43287, w_eco43288, w_eco43289, w_eco43290, w_eco43291, w_eco43292, w_eco43293, w_eco43294, w_eco43295, w_eco43296, w_eco43297, w_eco43298, w_eco43299, w_eco43300, w_eco43301, w_eco43302, w_eco43303, w_eco43304, w_eco43305, w_eco43306, w_eco43307, w_eco43308, w_eco43309, w_eco43310, w_eco43311, w_eco43312, w_eco43313, w_eco43314, w_eco43315, w_eco43316, w_eco43317, w_eco43318, w_eco43319, w_eco43320, w_eco43321, w_eco43322, w_eco43323, w_eco43324, w_eco43325, w_eco43326, w_eco43327, w_eco43328, w_eco43329, w_eco43330, w_eco43331, w_eco43332, w_eco43333, w_eco43334, w_eco43335, w_eco43336, w_eco43337, w_eco43338, w_eco43339, w_eco43340, w_eco43341, w_eco43342, w_eco43343, w_eco43344, w_eco43345, w_eco43346, w_eco43347, w_eco43348, w_eco43349, w_eco43350, w_eco43351, w_eco43352, w_eco43353, w_eco43354, w_eco43355, w_eco43356, w_eco43357, w_eco43358, w_eco43359, w_eco43360, w_eco43361, w_eco43362, w_eco43363, w_eco43364, w_eco43365, w_eco43366, w_eco43367, w_eco43368, w_eco43369, w_eco43370, w_eco43371, w_eco43372, w_eco43373, w_eco43374, w_eco43375, w_eco43376, w_eco43377, w_eco43378, w_eco43379, w_eco43380, w_eco43381, w_eco43382, w_eco43383, w_eco43384, w_eco43385, w_eco43386, w_eco43387, w_eco43388, w_eco43389, w_eco43390, w_eco43391, w_eco43392, w_eco43393, w_eco43394, w_eco43395, w_eco43396, w_eco43397, w_eco43398, w_eco43399, w_eco43400, w_eco43401, w_eco43402, w_eco43403, w_eco43404, w_eco43405, w_eco43406, w_eco43407, w_eco43408, w_eco43409, w_eco43410, w_eco43411, w_eco43412, w_eco43413, w_eco43414, w_eco43415, w_eco43416, w_eco43417, w_eco43418, w_eco43419, w_eco43420, w_eco43421, w_eco43422, w_eco43423, w_eco43424, w_eco43425, w_eco43426, w_eco43427, w_eco43428, w_eco43429, w_eco43430, w_eco43431, w_eco43432, w_eco43433, w_eco43434, w_eco43435, w_eco43436, w_eco43437, w_eco43438, w_eco43439, w_eco43440, w_eco43441, w_eco43442, w_eco43443, w_eco43444, w_eco43445, w_eco43446, w_eco43447, w_eco43448, w_eco43449, w_eco43450, w_eco43451, w_eco43452, w_eco43453, w_eco43454, w_eco43455, w_eco43456, w_eco43457, w_eco43458, w_eco43459, w_eco43460, w_eco43461, w_eco43462, w_eco43463, w_eco43464, w_eco43465, w_eco43466, w_eco43467, w_eco43468, w_eco43469, w_eco43470, w_eco43471, w_eco43472, w_eco43473, w_eco43474, w_eco43475, w_eco43476, w_eco43477, w_eco43478, w_eco43479, w_eco43480, w_eco43481, w_eco43482, w_eco43483, w_eco43484, w_eco43485, w_eco43486, w_eco43487, w_eco43488, w_eco43489, w_eco43490, w_eco43491, w_eco43492, w_eco43493, w_eco43494, w_eco43495, w_eco43496, w_eco43497, w_eco43498, w_eco43499, w_eco43500, w_eco43501, w_eco43502, w_eco43503, w_eco43504, w_eco43505, w_eco43506, w_eco43507, w_eco43508, w_eco43509, w_eco43510, w_eco43511, w_eco43512, w_eco43513, w_eco43514, w_eco43515, w_eco43516, w_eco43517, w_eco43518, w_eco43519, w_eco43520, w_eco43521, w_eco43522, w_eco43523, w_eco43524, w_eco43525, w_eco43526, w_eco43527, w_eco43528, w_eco43529, w_eco43530, w_eco43531, w_eco43532, w_eco43533, w_eco43534, w_eco43535, w_eco43536, w_eco43537, w_eco43538, w_eco43539, w_eco43540, w_eco43541, w_eco43542, w_eco43543, w_eco43544, w_eco43545, w_eco43546, w_eco43547, w_eco43548, w_eco43549, w_eco43550, w_eco43551, w_eco43552, w_eco43553, w_eco43554, w_eco43555, w_eco43556, w_eco43557, w_eco43558, w_eco43559, w_eco43560, w_eco43561, w_eco43562, w_eco43563, w_eco43564, w_eco43565, w_eco43566, w_eco43567, w_eco43568, w_eco43569, w_eco43570, w_eco43571, w_eco43572, w_eco43573, w_eco43574, w_eco43575, w_eco43576, w_eco43577, w_eco43578, w_eco43579, w_eco43580, w_eco43581, w_eco43582, w_eco43583, w_eco43584, w_eco43585, w_eco43586, w_eco43587, w_eco43588, w_eco43589, w_eco43590, w_eco43591, w_eco43592, w_eco43593, w_eco43594, w_eco43595, w_eco43596, w_eco43597, w_eco43598, w_eco43599, w_eco43600, w_eco43601, w_eco43602, w_eco43603, w_eco43604, w_eco43605, w_eco43606, w_eco43607, w_eco43608, w_eco43609, w_eco43610, w_eco43611, w_eco43612, w_eco43613, w_eco43614, w_eco43615, w_eco43616, w_eco43617, w_eco43618, w_eco43619, w_eco43620, w_eco43621, w_eco43622, w_eco43623, w_eco43624, w_eco43625, w_eco43626, w_eco43627, w_eco43628, w_eco43629, w_eco43630, w_eco43631, w_eco43632, w_eco43633, w_eco43634, w_eco43635, w_eco43636, w_eco43637, w_eco43638, w_eco43639, w_eco43640, w_eco43641, w_eco43642, w_eco43643, w_eco43644, w_eco43645, w_eco43646, w_eco43647, w_eco43648, w_eco43649, w_eco43650, w_eco43651, w_eco43652, w_eco43653, w_eco43654, w_eco43655, w_eco43656, w_eco43657, w_eco43658, w_eco43659, w_eco43660, w_eco43661, w_eco43662, w_eco43663, w_eco43664, w_eco43665, w_eco43666, w_eco43667, w_eco43668, w_eco43669, w_eco43670, w_eco43671, w_eco43672, w_eco43673, w_eco43674, w_eco43675, w_eco43676, w_eco43677, w_eco43678, w_eco43679, w_eco43680, w_eco43681, w_eco43682, w_eco43683, w_eco43684, w_eco43685, w_eco43686, w_eco43687, w_eco43688, w_eco43689, w_eco43690, w_eco43691, w_eco43692, w_eco43693, w_eco43694, w_eco43695, w_eco43696, w_eco43697, w_eco43698, w_eco43699, w_eco43700, w_eco43701, w_eco43702, w_eco43703, w_eco43704, w_eco43705, w_eco43706, w_eco43707, w_eco43708, w_eco43709, w_eco43710, w_eco43711, w_eco43712, w_eco43713, w_eco43714, w_eco43715, w_eco43716, w_eco43717, w_eco43718, w_eco43719, w_eco43720, w_eco43721, w_eco43722, w_eco43723, w_eco43724, w_eco43725, w_eco43726, w_eco43727, w_eco43728, w_eco43729, w_eco43730, w_eco43731, w_eco43732, w_eco43733, w_eco43734, w_eco43735, w_eco43736, w_eco43737, w_eco43738, w_eco43739, w_eco43740, w_eco43741, w_eco43742, w_eco43743, w_eco43744, w_eco43745, w_eco43746, w_eco43747, w_eco43748, w_eco43749, w_eco43750, w_eco43751, w_eco43752, w_eco43753, w_eco43754, w_eco43755, w_eco43756, w_eco43757, w_eco43758, w_eco43759, w_eco43760, w_eco43761, w_eco43762, w_eco43763, w_eco43764, w_eco43765, w_eco43766, w_eco43767, w_eco43768, w_eco43769, w_eco43770, w_eco43771, w_eco43772, w_eco43773, w_eco43774, w_eco43775, w_eco43776, w_eco43777, w_eco43778, w_eco43779, w_eco43780, w_eco43781, w_eco43782, w_eco43783, w_eco43784, w_eco43785, w_eco43786, w_eco43787, w_eco43788, w_eco43789, w_eco43790, w_eco43791, w_eco43792, w_eco43793, w_eco43794, w_eco43795, w_eco43796, w_eco43797, w_eco43798, w_eco43799, w_eco43800, w_eco43801, w_eco43802, w_eco43803, w_eco43804, w_eco43805, w_eco43806, w_eco43807, w_eco43808, w_eco43809, w_eco43810, w_eco43811, w_eco43812, w_eco43813, w_eco43814, w_eco43815, w_eco43816, w_eco43817, w_eco43818, w_eco43819, w_eco43820, w_eco43821, w_eco43822, w_eco43823, w_eco43824, w_eco43825, w_eco43826, w_eco43827, w_eco43828, w_eco43829, w_eco43830, w_eco43831, w_eco43832, w_eco43833, w_eco43834, w_eco43835, w_eco43836, w_eco43837, w_eco43838, w_eco43839, w_eco43840, w_eco43841, w_eco43842, w_eco43843, w_eco43844, w_eco43845, w_eco43846, w_eco43847, w_eco43848, w_eco43849, w_eco43850, w_eco43851, w_eco43852, w_eco43853, w_eco43854, w_eco43855, w_eco43856, w_eco43857, w_eco43858, w_eco43859, w_eco43860, w_eco43861, w_eco43862, w_eco43863, w_eco43864, w_eco43865, w_eco43866, w_eco43867, w_eco43868, w_eco43869, w_eco43870, w_eco43871, w_eco43872, w_eco43873, w_eco43874, w_eco43875, w_eco43876, w_eco43877, w_eco43878, w_eco43879, w_eco43880, w_eco43881, w_eco43882, w_eco43883, w_eco43884, w_eco43885, w_eco43886, w_eco43887, w_eco43888, w_eco43889, w_eco43890, w_eco43891, w_eco43892, w_eco43893, w_eco43894, w_eco43895, w_eco43896, w_eco43897, w_eco43898, w_eco43899, w_eco43900, w_eco43901, w_eco43902, w_eco43903, w_eco43904, w_eco43905, w_eco43906, w_eco43907, w_eco43908, w_eco43909, w_eco43910, w_eco43911, w_eco43912, w_eco43913, w_eco43914, w_eco43915, w_eco43916, w_eco43917, w_eco43918, w_eco43919, w_eco43920, w_eco43921, w_eco43922, w_eco43923, w_eco43924, w_eco43925, w_eco43926, w_eco43927, w_eco43928, w_eco43929, w_eco43930, w_eco43931, w_eco43932, w_eco43933, w_eco43934, w_eco43935, w_eco43936, w_eco43937, w_eco43938, w_eco43939, w_eco43940, w_eco43941, w_eco43942, w_eco43943, w_eco43944, w_eco43945, w_eco43946, w_eco43947, w_eco43948, w_eco43949, w_eco43950, w_eco43951, w_eco43952, w_eco43953, w_eco43954, w_eco43955, w_eco43956, w_eco43957, w_eco43958, w_eco43959, w_eco43960, w_eco43961, w_eco43962, w_eco43963, w_eco43964, w_eco43965, w_eco43966, w_eco43967, w_eco43968, w_eco43969, w_eco43970, w_eco43971, w_eco43972, w_eco43973, w_eco43974, w_eco43975, w_eco43976, w_eco43977, w_eco43978, w_eco43979, w_eco43980, w_eco43981, w_eco43982, w_eco43983, w_eco43984, w_eco43985, w_eco43986, w_eco43987, w_eco43988, w_eco43989, w_eco43990, w_eco43991, w_eco43992, w_eco43993, w_eco43994, w_eco43995, w_eco43996, w_eco43997, w_eco43998, w_eco43999, w_eco44000, w_eco44001, w_eco44002, w_eco44003, w_eco44004, w_eco44005, w_eco44006, w_eco44007, w_eco44008, w_eco44009, w_eco44010, w_eco44011, w_eco44012, w_eco44013, w_eco44014, w_eco44015, w_eco44016, w_eco44017, w_eco44018, w_eco44019, w_eco44020, w_eco44021, w_eco44022, w_eco44023, w_eco44024, w_eco44025, w_eco44026, w_eco44027, w_eco44028, w_eco44029, w_eco44030, w_eco44031, w_eco44032, w_eco44033, w_eco44034, w_eco44035, w_eco44036, w_eco44037, w_eco44038, w_eco44039, w_eco44040, w_eco44041, w_eco44042, w_eco44043, w_eco44044, w_eco44045, w_eco44046, w_eco44047, w_eco44048, w_eco44049, w_eco44050, w_eco44051, w_eco44052, w_eco44053, w_eco44054, w_eco44055, w_eco44056, w_eco44057, w_eco44058, w_eco44059, w_eco44060, w_eco44061, w_eco44062, w_eco44063, w_eco44064, w_eco44065, w_eco44066, w_eco44067, w_eco44068, w_eco44069, w_eco44070, w_eco44071, w_eco44072, w_eco44073, w_eco44074, w_eco44075, w_eco44076, w_eco44077, w_eco44078, w_eco44079, w_eco44080, w_eco44081, w_eco44082, w_eco44083, w_eco44084, w_eco44085, w_eco44086, w_eco44087, w_eco44088, w_eco44089, w_eco44090, w_eco44091, w_eco44092, w_eco44093, w_eco44094, w_eco44095, w_eco44096, w_eco44097, w_eco44098, w_eco44099, w_eco44100, w_eco44101, w_eco44102, w_eco44103, w_eco44104, w_eco44105, w_eco44106, w_eco44107, w_eco44108, w_eco44109, w_eco44110, w_eco44111, w_eco44112, w_eco44113, w_eco44114, w_eco44115, w_eco44116, w_eco44117, w_eco44118, w_eco44119, w_eco44120, w_eco44121, w_eco44122, w_eco44123, w_eco44124, w_eco44125, w_eco44126, w_eco44127, w_eco44128, w_eco44129, w_eco44130, w_eco44131, w_eco44132, w_eco44133, w_eco44134, w_eco44135, w_eco44136, w_eco44137, w_eco44138, w_eco44139, w_eco44140, w_eco44141, w_eco44142, w_eco44143, w_eco44144, w_eco44145, w_eco44146, w_eco44147, w_eco44148, w_eco44149, w_eco44150, w_eco44151, w_eco44152, w_eco44153, w_eco44154, w_eco44155, w_eco44156, w_eco44157, w_eco44158, w_eco44159, w_eco44160, w_eco44161, w_eco44162, w_eco44163, w_eco44164, w_eco44165, w_eco44166, w_eco44167, w_eco44168, w_eco44169, w_eco44170, w_eco44171, w_eco44172, w_eco44173, w_eco44174, w_eco44175, w_eco44176, w_eco44177, w_eco44178, w_eco44179, w_eco44180, w_eco44181, w_eco44182, w_eco44183, w_eco44184, w_eco44185, w_eco44186, w_eco44187, w_eco44188, w_eco44189, w_eco44190, w_eco44191, w_eco44192, w_eco44193, w_eco44194, w_eco44195, w_eco44196, w_eco44197, w_eco44198, w_eco44199, w_eco44200, w_eco44201, w_eco44202, w_eco44203, w_eco44204, w_eco44205, w_eco44206, w_eco44207, w_eco44208, w_eco44209, w_eco44210, w_eco44211, w_eco44212, w_eco44213, w_eco44214, w_eco44215, w_eco44216, w_eco44217, w_eco44218, w_eco44219, w_eco44220, w_eco44221, w_eco44222, w_eco44223, w_eco44224, w_eco44225, w_eco44226, w_eco44227, w_eco44228, w_eco44229, w_eco44230, w_eco44231, w_eco44232, w_eco44233, w_eco44234, w_eco44235, w_eco44236, w_eco44237, w_eco44238, w_eco44239, w_eco44240, w_eco44241, w_eco44242, w_eco44243, w_eco44244, w_eco44245, w_eco44246, w_eco44247, w_eco44248, w_eco44249, w_eco44250, w_eco44251, w_eco44252, w_eco44253, w_eco44254, w_eco44255, w_eco44256, w_eco44257, w_eco44258, w_eco44259, w_eco44260, w_eco44261, w_eco44262, w_eco44263, w_eco44264, w_eco44265, w_eco44266, w_eco44267, w_eco44268, w_eco44269, w_eco44270, w_eco44271, w_eco44272, w_eco44273, w_eco44274, w_eco44275, w_eco44276, w_eco44277, w_eco44278, w_eco44279, w_eco44280, w_eco44281, w_eco44282, w_eco44283, w_eco44284, w_eco44285, w_eco44286, w_eco44287, w_eco44288, w_eco44289, w_eco44290, w_eco44291, w_eco44292, w_eco44293, w_eco44294, w_eco44295, w_eco44296, w_eco44297, w_eco44298, w_eco44299, w_eco44300, w_eco44301, w_eco44302, w_eco44303, w_eco44304, w_eco44305, w_eco44306, w_eco44307, w_eco44308, w_eco44309, w_eco44310, w_eco44311, w_eco44312, w_eco44313, w_eco44314, w_eco44315, w_eco44316, w_eco44317, w_eco44318, w_eco44319, w_eco44320, w_eco44321, w_eco44322, w_eco44323, w_eco44324, w_eco44325, w_eco44326, w_eco44327, w_eco44328, w_eco44329, w_eco44330, w_eco44331, w_eco44332, w_eco44333, w_eco44334, w_eco44335, w_eco44336, w_eco44337, w_eco44338, w_eco44339, w_eco44340, w_eco44341, w_eco44342, w_eco44343, w_eco44344, w_eco44345, w_eco44346, w_eco44347, w_eco44348, w_eco44349, w_eco44350, w_eco44351, w_eco44352, w_eco44353, w_eco44354, w_eco44355, w_eco44356, w_eco44357, w_eco44358, w_eco44359, w_eco44360, w_eco44361, w_eco44362, w_eco44363, w_eco44364, w_eco44365, w_eco44366, w_eco44367, w_eco44368, w_eco44369, w_eco44370, w_eco44371, w_eco44372, w_eco44373, w_eco44374, w_eco44375, w_eco44376, w_eco44377, w_eco44378, w_eco44379, w_eco44380, w_eco44381, w_eco44382, w_eco44383, w_eco44384, w_eco44385, w_eco44386, w_eco44387, w_eco44388, w_eco44389, w_eco44390, w_eco44391, w_eco44392, w_eco44393, w_eco44394, w_eco44395, w_eco44396, w_eco44397, w_eco44398, w_eco44399, w_eco44400, w_eco44401, w_eco44402, w_eco44403, w_eco44404, w_eco44405, w_eco44406, w_eco44407, w_eco44408, w_eco44409, w_eco44410, w_eco44411, w_eco44412, w_eco44413, w_eco44414, w_eco44415, w_eco44416, w_eco44417, w_eco44418, w_eco44419, w_eco44420, w_eco44421, w_eco44422, w_eco44423, w_eco44424, w_eco44425, w_eco44426, w_eco44427, w_eco44428, w_eco44429, w_eco44430, w_eco44431, w_eco44432, w_eco44433, w_eco44434, w_eco44435, w_eco44436, w_eco44437, w_eco44438, w_eco44439, w_eco44440, w_eco44441, w_eco44442, w_eco44443, w_eco44444, w_eco44445, w_eco44446, w_eco44447, w_eco44448, w_eco44449, w_eco44450, w_eco44451, w_eco44452, w_eco44453, w_eco44454, w_eco44455, w_eco44456, w_eco44457, w_eco44458, w_eco44459, w_eco44460, w_eco44461, w_eco44462, w_eco44463, w_eco44464, w_eco44465, w_eco44466, w_eco44467, w_eco44468, w_eco44469, w_eco44470, w_eco44471, w_eco44472, w_eco44473, w_eco44474, w_eco44475, w_eco44476, w_eco44477, w_eco44478, w_eco44479, w_eco44480, w_eco44481, w_eco44482, w_eco44483, w_eco44484, w_eco44485, w_eco44486, w_eco44487, w_eco44488, w_eco44489, w_eco44490, w_eco44491, w_eco44492, w_eco44493, w_eco44494, w_eco44495, w_eco44496, w_eco44497, w_eco44498, w_eco44499, w_eco44500, w_eco44501, w_eco44502, w_eco44503, w_eco44504, w_eco44505, w_eco44506, w_eco44507, w_eco44508, w_eco44509, w_eco44510, w_eco44511, w_eco44512, w_eco44513, w_eco44514, w_eco44515, w_eco44516, w_eco44517, w_eco44518, w_eco44519, w_eco44520, w_eco44521, w_eco44522, w_eco44523, w_eco44524, w_eco44525, w_eco44526, w_eco44527, w_eco44528, w_eco44529, w_eco44530, w_eco44531, w_eco44532, w_eco44533, w_eco44534, w_eco44535, w_eco44536, w_eco44537, w_eco44538, w_eco44539, w_eco44540, w_eco44541, w_eco44542, w_eco44543, w_eco44544, w_eco44545, w_eco44546, w_eco44547, w_eco44548, w_eco44549, w_eco44550, w_eco44551, w_eco44552, w_eco44553, w_eco44554, w_eco44555, w_eco44556, w_eco44557, w_eco44558, w_eco44559, w_eco44560, w_eco44561, w_eco44562, w_eco44563, w_eco44564, w_eco44565, w_eco44566, w_eco44567, w_eco44568, w_eco44569, w_eco44570, w_eco44571, w_eco44572, w_eco44573, w_eco44574, w_eco44575, w_eco44576, w_eco44577, w_eco44578, w_eco44579, w_eco44580, w_eco44581, w_eco44582, w_eco44583, w_eco44584, w_eco44585, w_eco44586, w_eco44587, w_eco44588, w_eco44589, w_eco44590, w_eco44591, w_eco44592, w_eco44593, w_eco44594, w_eco44595, w_eco44596, w_eco44597, w_eco44598, w_eco44599, w_eco44600, w_eco44601, w_eco44602, w_eco44603, w_eco44604, w_eco44605, w_eco44606, w_eco44607, w_eco44608, w_eco44609, w_eco44610, w_eco44611, w_eco44612, w_eco44613, w_eco44614, w_eco44615, w_eco44616, w_eco44617, w_eco44618, w_eco44619, w_eco44620, w_eco44621, w_eco44622, w_eco44623, w_eco44624, w_eco44625, w_eco44626, w_eco44627, w_eco44628, w_eco44629, w_eco44630, w_eco44631, w_eco44632, w_eco44633, w_eco44634, w_eco44635, w_eco44636, w_eco44637, w_eco44638, w_eco44639, w_eco44640, w_eco44641, w_eco44642, w_eco44643, w_eco44644, w_eco44645, w_eco44646, w_eco44647, w_eco44648, w_eco44649, w_eco44650, w_eco44651, w_eco44652, w_eco44653, w_eco44654, w_eco44655, w_eco44656, w_eco44657, w_eco44658, w_eco44659, w_eco44660, w_eco44661, w_eco44662, w_eco44663, w_eco44664, w_eco44665, w_eco44666, w_eco44667, w_eco44668, w_eco44669, w_eco44670, w_eco44671, w_eco44672, w_eco44673, w_eco44674, w_eco44675, w_eco44676, w_eco44677, w_eco44678, w_eco44679, w_eco44680, w_eco44681, w_eco44682, w_eco44683, w_eco44684, w_eco44685, w_eco44686, w_eco44687, w_eco44688, w_eco44689, w_eco44690, w_eco44691, w_eco44692, w_eco44693, w_eco44694, w_eco44695, w_eco44696, w_eco44697, w_eco44698, w_eco44699, w_eco44700, w_eco44701, w_eco44702, w_eco44703, w_eco44704, w_eco44705, w_eco44706, w_eco44707, w_eco44708, w_eco44709, w_eco44710, w_eco44711, w_eco44712, w_eco44713, w_eco44714, w_eco44715, w_eco44716, w_eco44717, w_eco44718, w_eco44719, w_eco44720, w_eco44721, w_eco44722, w_eco44723, w_eco44724, w_eco44725, w_eco44726, w_eco44727, w_eco44728, w_eco44729, w_eco44730, w_eco44731, w_eco44732, w_eco44733, w_eco44734, w_eco44735, w_eco44736, w_eco44737, w_eco44738, w_eco44739, w_eco44740, w_eco44741, w_eco44742, w_eco44743, w_eco44744, w_eco44745, w_eco44746, w_eco44747, w_eco44748, w_eco44749, w_eco44750, w_eco44751, w_eco44752, w_eco44753, w_eco44754, w_eco44755, w_eco44756, w_eco44757, w_eco44758, w_eco44759, w_eco44760, w_eco44761, w_eco44762, w_eco44763, w_eco44764, w_eco44765, w_eco44766, w_eco44767, w_eco44768, w_eco44769, w_eco44770, w_eco44771, w_eco44772, w_eco44773, w_eco44774, w_eco44775, w_eco44776, w_eco44777, w_eco44778, w_eco44779, w_eco44780, w_eco44781, w_eco44782, w_eco44783, w_eco44784, w_eco44785, w_eco44786, w_eco44787, w_eco44788, w_eco44789, w_eco44790, w_eco44791, w_eco44792, w_eco44793, w_eco44794, w_eco44795, w_eco44796, w_eco44797, w_eco44798, w_eco44799, w_eco44800, w_eco44801, w_eco44802, w_eco44803, w_eco44804, w_eco44805, w_eco44806, w_eco44807, w_eco44808, w_eco44809, w_eco44810, w_eco44811, w_eco44812, w_eco44813, w_eco44814, w_eco44815, w_eco44816, w_eco44817, w_eco44818, w_eco44819, w_eco44820, w_eco44821, w_eco44822, w_eco44823, w_eco44824, w_eco44825, w_eco44826, w_eco44827, w_eco44828, w_eco44829, w_eco44830, w_eco44831, w_eco44832, w_eco44833, w_eco44834, w_eco44835, w_eco44836, w_eco44837, w_eco44838, w_eco44839, w_eco44840, w_eco44841, w_eco44842, w_eco44843, w_eco44844, w_eco44845, w_eco44846, w_eco44847, w_eco44848, w_eco44849, w_eco44850, w_eco44851, w_eco44852, w_eco44853, w_eco44854, w_eco44855, w_eco44856, w_eco44857, w_eco44858, w_eco44859, w_eco44860, w_eco44861, w_eco44862, w_eco44863, w_eco44864, w_eco44865, w_eco44866, w_eco44867, w_eco44868, w_eco44869, w_eco44870, w_eco44871, w_eco44872, w_eco44873, w_eco44874, w_eco44875, w_eco44876, w_eco44877, w_eco44878, w_eco44879, w_eco44880, w_eco44881, w_eco44882, w_eco44883, w_eco44884, w_eco44885, w_eco44886, w_eco44887, w_eco44888, w_eco44889, w_eco44890, w_eco44891, w_eco44892, w_eco44893, w_eco44894, w_eco44895, w_eco44896, w_eco44897, w_eco44898, w_eco44899, w_eco44900, w_eco44901, w_eco44902, w_eco44903, w_eco44904, w_eco44905, w_eco44906, w_eco44907, w_eco44908, w_eco44909, w_eco44910, w_eco44911, w_eco44912, w_eco44913, w_eco44914, w_eco44915, w_eco44916, w_eco44917, w_eco44918, w_eco44919, w_eco44920, w_eco44921, w_eco44922, w_eco44923, w_eco44924, w_eco44925, w_eco44926, w_eco44927, w_eco44928, w_eco44929, w_eco44930, w_eco44931, w_eco44932, w_eco44933, w_eco44934, w_eco44935, w_eco44936, w_eco44937, w_eco44938, w_eco44939, w_eco44940, w_eco44941, w_eco44942, w_eco44943, w_eco44944, w_eco44945, w_eco44946, w_eco44947, w_eco44948, w_eco44949, w_eco44950, w_eco44951, w_eco44952, w_eco44953, w_eco44954, w_eco44955, w_eco44956, w_eco44957, w_eco44958, w_eco44959, w_eco44960, w_eco44961, w_eco44962, w_eco44963, w_eco44964, w_eco44965, w_eco44966, w_eco44967, w_eco44968, w_eco44969, w_eco44970, w_eco44971, w_eco44972, w_eco44973, w_eco44974, w_eco44975, w_eco44976, w_eco44977, w_eco44978, w_eco44979, w_eco44980, w_eco44981, w_eco44982, w_eco44983, w_eco44984, w_eco44985, w_eco44986, w_eco44987, w_eco44988, w_eco44989, w_eco44990, w_eco44991, w_eco44992, w_eco44993, w_eco44994, w_eco44995, w_eco44996, w_eco44997, w_eco44998, w_eco44999, w_eco45000, w_eco45001, w_eco45002, w_eco45003, w_eco45004, w_eco45005, w_eco45006, w_eco45007, w_eco45008, w_eco45009, w_eco45010, w_eco45011, w_eco45012, w_eco45013, w_eco45014, w_eco45015, w_eco45016, w_eco45017, w_eco45018, w_eco45019, w_eco45020, w_eco45021, w_eco45022, w_eco45023, w_eco45024, w_eco45025, w_eco45026, w_eco45027, w_eco45028, w_eco45029, w_eco45030, w_eco45031, w_eco45032, w_eco45033, w_eco45034, w_eco45035, w_eco45036, w_eco45037, w_eco45038, w_eco45039, w_eco45040, w_eco45041, w_eco45042, w_eco45043, w_eco45044, w_eco45045, w_eco45046, w_eco45047, w_eco45048, w_eco45049, w_eco45050, w_eco45051, w_eco45052, w_eco45053, w_eco45054, w_eco45055, w_eco45056, w_eco45057, w_eco45058, w_eco45059, w_eco45060, w_eco45061, w_eco45062, w_eco45063, w_eco45064, w_eco45065, w_eco45066, w_eco45067, w_eco45068, w_eco45069, w_eco45070, w_eco45071, w_eco45072, w_eco45073, w_eco45074, w_eco45075, w_eco45076, w_eco45077, w_eco45078, w_eco45079, w_eco45080, w_eco45081, w_eco45082, w_eco45083, w_eco45084, w_eco45085, w_eco45086, w_eco45087, w_eco45088, w_eco45089, w_eco45090, w_eco45091, w_eco45092, w_eco45093, w_eco45094, w_eco45095, w_eco45096, w_eco45097, w_eco45098, w_eco45099, w_eco45100, w_eco45101, w_eco45102, w_eco45103, w_eco45104, w_eco45105, w_eco45106, w_eco45107, w_eco45108, w_eco45109, w_eco45110, w_eco45111, w_eco45112, w_eco45113, w_eco45114, w_eco45115, w_eco45116, w_eco45117, w_eco45118, w_eco45119, w_eco45120, w_eco45121, w_eco45122, w_eco45123, w_eco45124, w_eco45125, w_eco45126, w_eco45127, w_eco45128, w_eco45129, w_eco45130, w_eco45131, w_eco45132, w_eco45133, w_eco45134, w_eco45135, w_eco45136, w_eco45137, w_eco45138, w_eco45139, w_eco45140, w_eco45141, w_eco45142, w_eco45143, w_eco45144, w_eco45145, w_eco45146, w_eco45147, w_eco45148, w_eco45149, w_eco45150, w_eco45151, w_eco45152, w_eco45153, w_eco45154, w_eco45155, w_eco45156, w_eco45157, w_eco45158, w_eco45159, w_eco45160, w_eco45161, w_eco45162, w_eco45163, w_eco45164, w_eco45165, w_eco45166, w_eco45167, w_eco45168, w_eco45169, w_eco45170, w_eco45171, w_eco45172, w_eco45173, w_eco45174, w_eco45175, w_eco45176, w_eco45177, w_eco45178, w_eco45179, w_eco45180, w_eco45181, w_eco45182, w_eco45183, w_eco45184, w_eco45185, w_eco45186, w_eco45187, w_eco45188, w_eco45189, w_eco45190, w_eco45191, w_eco45192, w_eco45193, w_eco45194, w_eco45195, w_eco45196, w_eco45197, w_eco45198, w_eco45199, w_eco45200, w_eco45201, w_eco45202, w_eco45203, w_eco45204, w_eco45205, w_eco45206, w_eco45207, w_eco45208, w_eco45209, w_eco45210, w_eco45211, w_eco45212, w_eco45213, w_eco45214, w_eco45215, w_eco45216, w_eco45217, w_eco45218, w_eco45219, w_eco45220, w_eco45221, w_eco45222, w_eco45223, w_eco45224, w_eco45225, w_eco45226, w_eco45227, w_eco45228, w_eco45229, w_eco45230, w_eco45231, w_eco45232, w_eco45233, w_eco45234, w_eco45235, w_eco45236, w_eco45237, w_eco45238, w_eco45239, w_eco45240, w_eco45241, w_eco45242, w_eco45243, w_eco45244, w_eco45245, w_eco45246, w_eco45247, w_eco45248, w_eco45249, w_eco45250, w_eco45251, w_eco45252, w_eco45253, w_eco45254, w_eco45255, w_eco45256, w_eco45257, w_eco45258, w_eco45259, w_eco45260, w_eco45261, w_eco45262, w_eco45263, w_eco45264, w_eco45265, w_eco45266, w_eco45267, w_eco45268, w_eco45269, w_eco45270, w_eco45271, w_eco45272, w_eco45273, w_eco45274, w_eco45275, w_eco45276, w_eco45277, w_eco45278, w_eco45279, w_eco45280, w_eco45281, w_eco45282, w_eco45283, w_eco45284, w_eco45285, w_eco45286, w_eco45287, w_eco45288, w_eco45289, w_eco45290, w_eco45291, w_eco45292, w_eco45293, w_eco45294, w_eco45295, w_eco45296, w_eco45297, w_eco45298, w_eco45299, w_eco45300, w_eco45301, w_eco45302, w_eco45303, w_eco45304, w_eco45305, w_eco45306, w_eco45307, w_eco45308, w_eco45309, w_eco45310, w_eco45311, w_eco45312, w_eco45313, w_eco45314, w_eco45315, w_eco45316, w_eco45317, w_eco45318, w_eco45319, w_eco45320, w_eco45321, w_eco45322, w_eco45323, w_eco45324, w_eco45325, w_eco45326, w_eco45327, w_eco45328, w_eco45329, w_eco45330, w_eco45331, w_eco45332, w_eco45333, w_eco45334, w_eco45335, w_eco45336, w_eco45337, w_eco45338, w_eco45339, w_eco45340, w_eco45341, w_eco45342, w_eco45343, w_eco45344, w_eco45345, w_eco45346, w_eco45347, w_eco45348, w_eco45349, w_eco45350, w_eco45351, w_eco45352, w_eco45353, w_eco45354, w_eco45355, w_eco45356, w_eco45357, w_eco45358, w_eco45359, w_eco45360, w_eco45361, w_eco45362, w_eco45363, w_eco45364, w_eco45365, w_eco45366, w_eco45367, w_eco45368, w_eco45369, w_eco45370, w_eco45371, w_eco45372, w_eco45373, w_eco45374, w_eco45375, w_eco45376, w_eco45377, w_eco45378, w_eco45379, w_eco45380, w_eco45381, w_eco45382, w_eco45383, w_eco45384, w_eco45385, w_eco45386, w_eco45387, w_eco45388, w_eco45389, w_eco45390, w_eco45391, w_eco45392, w_eco45393, w_eco45394, w_eco45395, w_eco45396, w_eco45397, w_eco45398, w_eco45399, w_eco45400, w_eco45401, w_eco45402, w_eco45403, w_eco45404, w_eco45405, w_eco45406, w_eco45407, w_eco45408, w_eco45409, w_eco45410, w_eco45411, w_eco45412, w_eco45413, w_eco45414, w_eco45415, w_eco45416, w_eco45417, w_eco45418, w_eco45419, w_eco45420, w_eco45421, w_eco45422, w_eco45423, w_eco45424, w_eco45425, w_eco45426, w_eco45427, w_eco45428, w_eco45429, w_eco45430, w_eco45431, w_eco45432, w_eco45433, w_eco45434, w_eco45435, w_eco45436, w_eco45437, w_eco45438, w_eco45439, w_eco45440, w_eco45441, w_eco45442, w_eco45443, w_eco45444, w_eco45445, w_eco45446, w_eco45447, w_eco45448, w_eco45449, w_eco45450, w_eco45451, w_eco45452, w_eco45453, w_eco45454, w_eco45455, w_eco45456, w_eco45457, w_eco45458, w_eco45459, w_eco45460, w_eco45461, w_eco45462, w_eco45463, w_eco45464, w_eco45465, w_eco45466, w_eco45467, w_eco45468, w_eco45469, w_eco45470, w_eco45471, w_eco45472, w_eco45473, w_eco45474, w_eco45475, w_eco45476, w_eco45477, w_eco45478, w_eco45479, w_eco45480, w_eco45481, w_eco45482, w_eco45483, w_eco45484, w_eco45485, w_eco45486, w_eco45487, w_eco45488, w_eco45489, w_eco45490, w_eco45491, w_eco45492, w_eco45493, w_eco45494, w_eco45495, w_eco45496, w_eco45497, w_eco45498, w_eco45499, w_eco45500, w_eco45501, w_eco45502, w_eco45503, w_eco45504, w_eco45505, w_eco45506, w_eco45507, w_eco45508, w_eco45509, w_eco45510, w_eco45511, w_eco45512, w_eco45513, w_eco45514, w_eco45515, w_eco45516, w_eco45517, w_eco45518, w_eco45519, w_eco45520, w_eco45521, w_eco45522, w_eco45523, w_eco45524, w_eco45525, w_eco45526, w_eco45527, w_eco45528, w_eco45529, w_eco45530, w_eco45531, w_eco45532, w_eco45533, w_eco45534, w_eco45535, w_eco45536, w_eco45537, w_eco45538, w_eco45539, w_eco45540, w_eco45541, w_eco45542, w_eco45543, w_eco45544, w_eco45545, w_eco45546, w_eco45547, w_eco45548, w_eco45549, w_eco45550, w_eco45551, w_eco45552, w_eco45553, w_eco45554, w_eco45555, w_eco45556, w_eco45557, w_eco45558, w_eco45559, w_eco45560, w_eco45561, w_eco45562, w_eco45563, w_eco45564, w_eco45565, w_eco45566, w_eco45567, w_eco45568, w_eco45569, w_eco45570, w_eco45571, w_eco45572, w_eco45573, w_eco45574, w_eco45575, w_eco45576, w_eco45577, w_eco45578, w_eco45579, w_eco45580, w_eco45581, w_eco45582, w_eco45583, w_eco45584, w_eco45585, w_eco45586, w_eco45587, w_eco45588, w_eco45589, w_eco45590, w_eco45591, w_eco45592, w_eco45593, w_eco45594, w_eco45595, w_eco45596, w_eco45597, w_eco45598, w_eco45599, w_eco45600, w_eco45601, w_eco45602, w_eco45603, w_eco45604, w_eco45605, w_eco45606, w_eco45607, w_eco45608, w_eco45609, w_eco45610, w_eco45611, w_eco45612, w_eco45613, w_eco45614, w_eco45615, w_eco45616, w_eco45617, w_eco45618, w_eco45619, w_eco45620, w_eco45621, w_eco45622, w_eco45623, w_eco45624, w_eco45625, w_eco45626, w_eco45627, w_eco45628, w_eco45629, w_eco45630, w_eco45631, w_eco45632, w_eco45633, w_eco45634, w_eco45635, w_eco45636, w_eco45637, w_eco45638, w_eco45639, w_eco45640, w_eco45641, w_eco45642, w_eco45643, w_eco45644, w_eco45645, w_eco45646, w_eco45647, w_eco45648, w_eco45649, w_eco45650, w_eco45651, w_eco45652, w_eco45653, w_eco45654, w_eco45655, w_eco45656, w_eco45657, w_eco45658, w_eco45659, w_eco45660, w_eco45661, w_eco45662, w_eco45663, w_eco45664, w_eco45665, w_eco45666, w_eco45667, w_eco45668, w_eco45669, w_eco45670, w_eco45671, w_eco45672, w_eco45673, w_eco45674, w_eco45675, w_eco45676, w_eco45677, w_eco45678, w_eco45679, w_eco45680, w_eco45681, w_eco45682, w_eco45683, w_eco45684, w_eco45685, w_eco45686, w_eco45687, w_eco45688, w_eco45689, w_eco45690, w_eco45691, w_eco45692, w_eco45693, w_eco45694, w_eco45695, w_eco45696, w_eco45697, w_eco45698, w_eco45699, w_eco45700, w_eco45701, w_eco45702, w_eco45703, w_eco45704, w_eco45705, w_eco45706, w_eco45707, w_eco45708, w_eco45709, w_eco45710, w_eco45711, w_eco45712, w_eco45713, w_eco45714, w_eco45715, w_eco45716, w_eco45717, w_eco45718, w_eco45719, w_eco45720, w_eco45721, w_eco45722, w_eco45723, w_eco45724, w_eco45725, w_eco45726, w_eco45727, w_eco45728, w_eco45729, w_eco45730, w_eco45731, w_eco45732, w_eco45733, w_eco45734, w_eco45735, w_eco45736, w_eco45737, w_eco45738, w_eco45739, w_eco45740, w_eco45741, w_eco45742, w_eco45743, w_eco45744, w_eco45745, w_eco45746, w_eco45747, w_eco45748, w_eco45749, w_eco45750, w_eco45751, w_eco45752, w_eco45753, w_eco45754, w_eco45755, w_eco45756, w_eco45757, w_eco45758, w_eco45759, w_eco45760, w_eco45761, w_eco45762, w_eco45763, w_eco45764, w_eco45765, w_eco45766, w_eco45767, w_eco45768, w_eco45769, w_eco45770, w_eco45771, w_eco45772, w_eco45773, w_eco45774, w_eco45775, w_eco45776, w_eco45777, w_eco45778, w_eco45779, w_eco45780, w_eco45781, w_eco45782, w_eco45783, w_eco45784, w_eco45785, w_eco45786, w_eco45787, w_eco45788, w_eco45789, w_eco45790, w_eco45791, w_eco45792, w_eco45793, w_eco45794, w_eco45795, w_eco45796, w_eco45797, w_eco45798, w_eco45799, w_eco45800, w_eco45801, w_eco45802, w_eco45803, w_eco45804, w_eco45805, w_eco45806, w_eco45807, w_eco45808, w_eco45809, w_eco45810, w_eco45811, w_eco45812, w_eco45813, w_eco45814, w_eco45815, w_eco45816, w_eco45817, w_eco45818, w_eco45819, w_eco45820, w_eco45821, w_eco45822, w_eco45823, w_eco45824, w_eco45825, w_eco45826, w_eco45827, w_eco45828, w_eco45829, w_eco45830, w_eco45831, w_eco45832, w_eco45833, w_eco45834, w_eco45835, w_eco45836, w_eco45837, w_eco45838, w_eco45839, w_eco45840, w_eco45841, w_eco45842, w_eco45843, w_eco45844, w_eco45845, w_eco45846, w_eco45847, w_eco45848, w_eco45849, w_eco45850, w_eco45851, w_eco45852, w_eco45853, w_eco45854, w_eco45855, w_eco45856, w_eco45857, w_eco45858, w_eco45859, w_eco45860, w_eco45861, w_eco45862, w_eco45863, w_eco45864, w_eco45865, w_eco45866, w_eco45867, w_eco45868, w_eco45869, w_eco45870, w_eco45871, w_eco45872, w_eco45873, w_eco45874, w_eco45875, w_eco45876, w_eco45877, w_eco45878, w_eco45879, w_eco45880, w_eco45881, w_eco45882, w_eco45883, w_eco45884, w_eco45885, w_eco45886, w_eco45887, w_eco45888, w_eco45889, w_eco45890, w_eco45891, w_eco45892, w_eco45893, w_eco45894, w_eco45895, w_eco45896, w_eco45897, w_eco45898, w_eco45899, w_eco45900, w_eco45901, w_eco45902, w_eco45903, w_eco45904, w_eco45905, w_eco45906, w_eco45907, w_eco45908, w_eco45909, w_eco45910, w_eco45911, w_eco45912, w_eco45913, w_eco45914, w_eco45915, w_eco45916, w_eco45917, w_eco45918, w_eco45919, w_eco45920, w_eco45921, w_eco45922, w_eco45923, w_eco45924, w_eco45925, w_eco45926, w_eco45927, w_eco45928, w_eco45929, w_eco45930, w_eco45931, w_eco45932, w_eco45933, w_eco45934, w_eco45935, w_eco45936, w_eco45937, w_eco45938, w_eco45939, w_eco45940, w_eco45941, w_eco45942, w_eco45943, w_eco45944, w_eco45945, w_eco45946, w_eco45947, w_eco45948, w_eco45949, w_eco45950, w_eco45951, w_eco45952, w_eco45953, w_eco45954, w_eco45955, w_eco45956, w_eco45957, w_eco45958, w_eco45959, w_eco45960, w_eco45961, w_eco45962, w_eco45963, w_eco45964, w_eco45965, w_eco45966, w_eco45967, w_eco45968, w_eco45969, w_eco45970, w_eco45971, w_eco45972, w_eco45973, w_eco45974, w_eco45975, w_eco45976, w_eco45977, w_eco45978, w_eco45979, w_eco45980, w_eco45981, w_eco45982, w_eco45983, w_eco45984, w_eco45985, w_eco45986, w_eco45987, w_eco45988, w_eco45989, w_eco45990, w_eco45991, w_eco45992, w_eco45993, w_eco45994, w_eco45995, w_eco45996, w_eco45997, w_eco45998, w_eco45999, w_eco46000, w_eco46001, w_eco46002, w_eco46003, w_eco46004, w_eco46005, w_eco46006, w_eco46007, w_eco46008, w_eco46009, w_eco46010, w_eco46011, w_eco46012, w_eco46013, w_eco46014, w_eco46015, w_eco46016, w_eco46017, w_eco46018, w_eco46019, w_eco46020, w_eco46021, w_eco46022, w_eco46023, w_eco46024, w_eco46025, w_eco46026, w_eco46027, w_eco46028, w_eco46029, w_eco46030, w_eco46031, w_eco46032, w_eco46033, w_eco46034, w_eco46035, w_eco46036, w_eco46037, w_eco46038, w_eco46039, w_eco46040, w_eco46041, w_eco46042, w_eco46043, w_eco46044, w_eco46045, w_eco46046, w_eco46047, w_eco46048, w_eco46049, w_eco46050, w_eco46051, w_eco46052, w_eco46053, w_eco46054, w_eco46055, w_eco46056, w_eco46057, w_eco46058, w_eco46059, w_eco46060, w_eco46061, w_eco46062, w_eco46063, w_eco46064, w_eco46065, w_eco46066, w_eco46067, w_eco46068, w_eco46069, w_eco46070, w_eco46071, w_eco46072, w_eco46073, w_eco46074, w_eco46075, w_eco46076, w_eco46077, w_eco46078, w_eco46079, w_eco46080, w_eco46081, w_eco46082, w_eco46083, w_eco46084, w_eco46085, w_eco46086, w_eco46087, w_eco46088, w_eco46089, w_eco46090, w_eco46091, w_eco46092, w_eco46093, w_eco46094, w_eco46095, w_eco46096, w_eco46097, w_eco46098, w_eco46099, w_eco46100, w_eco46101, w_eco46102, w_eco46103, w_eco46104, w_eco46105, w_eco46106, w_eco46107, w_eco46108, w_eco46109, w_eco46110, w_eco46111, w_eco46112, w_eco46113, w_eco46114, w_eco46115, w_eco46116, w_eco46117, w_eco46118, w_eco46119, w_eco46120, w_eco46121, w_eco46122, w_eco46123, w_eco46124, w_eco46125, w_eco46126, w_eco46127, w_eco46128, w_eco46129, w_eco46130, w_eco46131, w_eco46132, w_eco46133, w_eco46134, w_eco46135, w_eco46136, w_eco46137, w_eco46138, w_eco46139, w_eco46140, w_eco46141, w_eco46142, w_eco46143, w_eco46144, w_eco46145, w_eco46146, w_eco46147, w_eco46148, w_eco46149, w_eco46150, w_eco46151, w_eco46152, w_eco46153, w_eco46154, w_eco46155, w_eco46156, w_eco46157, w_eco46158, w_eco46159, w_eco46160, w_eco46161, w_eco46162, w_eco46163, w_eco46164, w_eco46165, w_eco46166, w_eco46167, w_eco46168, w_eco46169, w_eco46170, w_eco46171, w_eco46172, w_eco46173, w_eco46174, w_eco46175, w_eco46176, w_eco46177, w_eco46178, w_eco46179, w_eco46180, w_eco46181, w_eco46182, w_eco46183, w_eco46184, w_eco46185, w_eco46186, w_eco46187, w_eco46188, w_eco46189, w_eco46190, w_eco46191, w_eco46192, w_eco46193, w_eco46194, w_eco46195, w_eco46196, w_eco46197, w_eco46198, w_eco46199, w_eco46200, w_eco46201, w_eco46202, w_eco46203, w_eco46204, w_eco46205, w_eco46206, w_eco46207, w_eco46208, w_eco46209, w_eco46210, w_eco46211, w_eco46212, w_eco46213, w_eco46214, w_eco46215, w_eco46216, w_eco46217, w_eco46218, w_eco46219, w_eco46220, w_eco46221, w_eco46222, w_eco46223, w_eco46224, w_eco46225, w_eco46226, w_eco46227, w_eco46228, w_eco46229, w_eco46230, w_eco46231, w_eco46232, w_eco46233, w_eco46234, w_eco46235, w_eco46236, w_eco46237, w_eco46238, w_eco46239, w_eco46240, w_eco46241, w_eco46242, w_eco46243, w_eco46244, w_eco46245, w_eco46246, w_eco46247, w_eco46248, w_eco46249, w_eco46250, w_eco46251, w_eco46252, w_eco46253, w_eco46254, w_eco46255, w_eco46256, w_eco46257, w_eco46258, w_eco46259, w_eco46260, w_eco46261, w_eco46262, w_eco46263, w_eco46264, w_eco46265, w_eco46266, w_eco46267, w_eco46268, w_eco46269, w_eco46270, w_eco46271, w_eco46272, w_eco46273, w_eco46274, w_eco46275, w_eco46276, w_eco46277, w_eco46278, w_eco46279, w_eco46280, w_eco46281, w_eco46282, w_eco46283, w_eco46284, w_eco46285, w_eco46286, w_eco46287, w_eco46288, w_eco46289, w_eco46290, w_eco46291, w_eco46292, w_eco46293, w_eco46294, w_eco46295, w_eco46296, w_eco46297, w_eco46298, w_eco46299, w_eco46300, w_eco46301, w_eco46302, w_eco46303, w_eco46304, w_eco46305, w_eco46306, w_eco46307, w_eco46308, w_eco46309, w_eco46310, w_eco46311, w_eco46312, w_eco46313, w_eco46314, w_eco46315, w_eco46316, w_eco46317, w_eco46318, w_eco46319, w_eco46320, w_eco46321, w_eco46322, w_eco46323, w_eco46324, w_eco46325, w_eco46326, w_eco46327, w_eco46328, w_eco46329, w_eco46330, w_eco46331, w_eco46332, w_eco46333, w_eco46334, w_eco46335, w_eco46336, w_eco46337, w_eco46338, w_eco46339, w_eco46340, w_eco46341, w_eco46342, w_eco46343, w_eco46344, w_eco46345, w_eco46346, w_eco46347, w_eco46348, w_eco46349, w_eco46350, w_eco46351, w_eco46352, w_eco46353, w_eco46354, w_eco46355, w_eco46356, w_eco46357, w_eco46358, w_eco46359, w_eco46360, w_eco46361, w_eco46362, w_eco46363, w_eco46364, w_eco46365, w_eco46366, w_eco46367, w_eco46368, w_eco46369, w_eco46370, w_eco46371, w_eco46372, w_eco46373, w_eco46374, w_eco46375, w_eco46376, w_eco46377, w_eco46378, w_eco46379, w_eco46380, w_eco46381, w_eco46382, w_eco46383, w_eco46384, w_eco46385, w_eco46386, w_eco46387, w_eco46388, w_eco46389, w_eco46390, w_eco46391, w_eco46392, w_eco46393, w_eco46394, w_eco46395, w_eco46396, w_eco46397, w_eco46398, w_eco46399, w_eco46400, w_eco46401, w_eco46402, w_eco46403, w_eco46404, w_eco46405, w_eco46406, w_eco46407, w_eco46408, w_eco46409, w_eco46410, w_eco46411, w_eco46412, w_eco46413, w_eco46414, w_eco46415, w_eco46416, w_eco46417, w_eco46418, w_eco46419, w_eco46420, w_eco46421, w_eco46422, w_eco46423, w_eco46424, w_eco46425, w_eco46426, w_eco46427, w_eco46428, w_eco46429, w_eco46430, w_eco46431, w_eco46432, w_eco46433, w_eco46434, w_eco46435, w_eco46436, w_eco46437, w_eco46438, w_eco46439, w_eco46440, w_eco46441, w_eco46442, w_eco46443, w_eco46444, w_eco46445, w_eco46446, w_eco46447, w_eco46448, w_eco46449, w_eco46450, w_eco46451, w_eco46452, w_eco46453, w_eco46454, w_eco46455, w_eco46456, w_eco46457, w_eco46458, w_eco46459, w_eco46460, w_eco46461, w_eco46462, w_eco46463, w_eco46464, w_eco46465, w_eco46466, w_eco46467, w_eco46468, w_eco46469, w_eco46470, w_eco46471, w_eco46472, w_eco46473, w_eco46474, w_eco46475, w_eco46476, w_eco46477, w_eco46478, w_eco46479, w_eco46480, w_eco46481, w_eco46482, w_eco46483, w_eco46484, w_eco46485, w_eco46486, w_eco46487, w_eco46488, w_eco46489, w_eco46490, w_eco46491, w_eco46492, w_eco46493, w_eco46494, w_eco46495, w_eco46496, w_eco46497, w_eco46498, w_eco46499, w_eco46500, w_eco46501, w_eco46502, w_eco46503, w_eco46504, w_eco46505, w_eco46506, w_eco46507, w_eco46508, w_eco46509, w_eco46510, w_eco46511, w_eco46512, w_eco46513, w_eco46514, w_eco46515, w_eco46516, w_eco46517, w_eco46518, w_eco46519, w_eco46520, w_eco46521, w_eco46522, w_eco46523, w_eco46524, w_eco46525, w_eco46526, w_eco46527, w_eco46528, w_eco46529, w_eco46530, w_eco46531, w_eco46532, w_eco46533, w_eco46534, w_eco46535, w_eco46536, w_eco46537, w_eco46538, w_eco46539, w_eco46540, w_eco46541, w_eco46542, w_eco46543, w_eco46544, w_eco46545, w_eco46546, w_eco46547, w_eco46548, w_eco46549, w_eco46550, w_eco46551, w_eco46552, w_eco46553, w_eco46554, w_eco46555, w_eco46556, w_eco46557, w_eco46558, w_eco46559, w_eco46560, w_eco46561, w_eco46562, w_eco46563, w_eco46564, w_eco46565, w_eco46566, w_eco46567, w_eco46568, w_eco46569, w_eco46570, w_eco46571, w_eco46572, w_eco46573, w_eco46574, w_eco46575, w_eco46576, w_eco46577, w_eco46578, w_eco46579, w_eco46580, w_eco46581, w_eco46582, w_eco46583, w_eco46584, w_eco46585, w_eco46586, w_eco46587, w_eco46588, w_eco46589, w_eco46590, w_eco46591, w_eco46592, w_eco46593, w_eco46594, w_eco46595, w_eco46596, w_eco46597, w_eco46598, w_eco46599, w_eco46600, w_eco46601, w_eco46602, w_eco46603, w_eco46604, w_eco46605, w_eco46606, w_eco46607, w_eco46608, w_eco46609, w_eco46610, w_eco46611, w_eco46612, w_eco46613, w_eco46614, w_eco46615, w_eco46616, w_eco46617, w_eco46618, w_eco46619, w_eco46620, w_eco46621, w_eco46622, w_eco46623, w_eco46624, w_eco46625, w_eco46626, w_eco46627, w_eco46628, w_eco46629, w_eco46630, w_eco46631, w_eco46632, w_eco46633, w_eco46634, w_eco46635, w_eco46636, w_eco46637, w_eco46638, w_eco46639, w_eco46640, w_eco46641, w_eco46642, w_eco46643, w_eco46644, w_eco46645, w_eco46646, w_eco46647, w_eco46648, w_eco46649, w_eco46650, w_eco46651, w_eco46652, w_eco46653, w_eco46654, w_eco46655, w_eco46656, w_eco46657, w_eco46658, w_eco46659, w_eco46660, w_eco46661, w_eco46662, w_eco46663, w_eco46664, w_eco46665, w_eco46666, w_eco46667, w_eco46668, w_eco46669, w_eco46670, w_eco46671, w_eco46672, w_eco46673, w_eco46674, w_eco46675, w_eco46676, w_eco46677, w_eco46678, w_eco46679, w_eco46680, w_eco46681, w_eco46682, w_eco46683, w_eco46684, w_eco46685, w_eco46686, w_eco46687, w_eco46688, w_eco46689, w_eco46690, w_eco46691, w_eco46692, w_eco46693, w_eco46694, w_eco46695, w_eco46696, w_eco46697, w_eco46698, w_eco46699, w_eco46700, w_eco46701, w_eco46702, w_eco46703, w_eco46704, w_eco46705, w_eco46706, w_eco46707, w_eco46708, w_eco46709, w_eco46710, w_eco46711, w_eco46712, w_eco46713, w_eco46714, w_eco46715, w_eco46716, w_eco46717, w_eco46718, w_eco46719, w_eco46720, w_eco46721, w_eco46722, w_eco46723, w_eco46724, w_eco46725, w_eco46726, w_eco46727, w_eco46728, w_eco46729, w_eco46730, w_eco46731, w_eco46732, w_eco46733, w_eco46734, w_eco46735, w_eco46736, w_eco46737, w_eco46738, w_eco46739, w_eco46740, w_eco46741, w_eco46742, w_eco46743, w_eco46744, w_eco46745, w_eco46746, w_eco46747, w_eco46748, w_eco46749, w_eco46750, w_eco46751, w_eco46752, w_eco46753, w_eco46754, w_eco46755, w_eco46756, w_eco46757, w_eco46758, w_eco46759, w_eco46760, w_eco46761, w_eco46762, w_eco46763, w_eco46764, w_eco46765, w_eco46766, w_eco46767, w_eco46768, w_eco46769, w_eco46770, w_eco46771, w_eco46772, w_eco46773, w_eco46774, w_eco46775, w_eco46776, w_eco46777, w_eco46778, w_eco46779, w_eco46780, w_eco46781, w_eco46782, w_eco46783, w_eco46784, w_eco46785, w_eco46786, w_eco46787, w_eco46788, w_eco46789, w_eco46790, w_eco46791, w_eco46792, w_eco46793, w_eco46794, w_eco46795, w_eco46796, w_eco46797, w_eco46798, w_eco46799, w_eco46800, w_eco46801, w_eco46802, w_eco46803, w_eco46804, w_eco46805, w_eco46806, w_eco46807, w_eco46808, w_eco46809, w_eco46810, w_eco46811, w_eco46812, w_eco46813, w_eco46814, w_eco46815, w_eco46816, w_eco46817, w_eco46818, w_eco46819, w_eco46820, w_eco46821, w_eco46822, w_eco46823, w_eco46824, w_eco46825, w_eco46826, w_eco46827, w_eco46828, w_eco46829, w_eco46830, w_eco46831, w_eco46832, w_eco46833, w_eco46834, w_eco46835, w_eco46836, w_eco46837, w_eco46838, w_eco46839, w_eco46840, w_eco46841, w_eco46842, w_eco46843, w_eco46844, w_eco46845, w_eco46846, w_eco46847, w_eco46848, w_eco46849, w_eco46850, w_eco46851, w_eco46852, w_eco46853, w_eco46854, w_eco46855, w_eco46856, w_eco46857, w_eco46858, w_eco46859, w_eco46860, w_eco46861, w_eco46862, w_eco46863, w_eco46864, w_eco46865, w_eco46866, w_eco46867, w_eco46868, w_eco46869, w_eco46870, w_eco46871, w_eco46872, w_eco46873, w_eco46874, w_eco46875, w_eco46876, w_eco46877, w_eco46878, w_eco46879, w_eco46880, w_eco46881, w_eco46882, w_eco46883, w_eco46884, w_eco46885, w_eco46886, w_eco46887, w_eco46888, w_eco46889, w_eco46890, w_eco46891, w_eco46892, w_eco46893, w_eco46894, w_eco46895, w_eco46896, w_eco46897, w_eco46898, w_eco46899, w_eco46900, w_eco46901, w_eco46902, w_eco46903, w_eco46904, w_eco46905, w_eco46906, w_eco46907, w_eco46908, w_eco46909, w_eco46910, w_eco46911, w_eco46912, w_eco46913, w_eco46914, w_eco46915, w_eco46916, w_eco46917, w_eco46918, w_eco46919, w_eco46920, w_eco46921, w_eco46922, w_eco46923, w_eco46924, w_eco46925, w_eco46926, w_eco46927, w_eco46928, w_eco46929, w_eco46930, w_eco46931, w_eco46932, w_eco46933, w_eco46934, w_eco46935, w_eco46936, w_eco46937, w_eco46938, w_eco46939, w_eco46940, w_eco46941, w_eco46942, w_eco46943, w_eco46944, w_eco46945, w_eco46946, w_eco46947, w_eco46948, w_eco46949, w_eco46950, w_eco46951, w_eco46952, w_eco46953, w_eco46954, w_eco46955, w_eco46956, w_eco46957, w_eco46958, w_eco46959, w_eco46960, w_eco46961, w_eco46962, w_eco46963, w_eco46964, w_eco46965, w_eco46966, w_eco46967, w_eco46968, w_eco46969, w_eco46970, w_eco46971, w_eco46972, w_eco46973, w_eco46974, w_eco46975, w_eco46976, w_eco46977, w_eco46978, w_eco46979, w_eco46980, w_eco46981, w_eco46982, w_eco46983, w_eco46984, w_eco46985, w_eco46986, w_eco46987, w_eco46988, w_eco46989, w_eco46990, w_eco46991, w_eco46992, w_eco46993, w_eco46994, w_eco46995, w_eco46996, w_eco46997, w_eco46998, w_eco46999, w_eco47000, w_eco47001, w_eco47002, w_eco47003, w_eco47004, w_eco47005, w_eco47006, w_eco47007, w_eco47008, w_eco47009, w_eco47010, w_eco47011, w_eco47012, w_eco47013, w_eco47014, w_eco47015, w_eco47016, w_eco47017, w_eco47018, w_eco47019, w_eco47020, w_eco47021, w_eco47022, w_eco47023, w_eco47024, w_eco47025, w_eco47026, w_eco47027, w_eco47028, w_eco47029, w_eco47030, w_eco47031, w_eco47032, w_eco47033, w_eco47034, w_eco47035, w_eco47036, w_eco47037, w_eco47038, w_eco47039, w_eco47040, w_eco47041, w_eco47042, w_eco47043, w_eco47044, w_eco47045, w_eco47046, w_eco47047, w_eco47048, w_eco47049, w_eco47050, w_eco47051, w_eco47052, w_eco47053, w_eco47054, w_eco47055, w_eco47056, w_eco47057, w_eco47058, w_eco47059, w_eco47060, w_eco47061, w_eco47062, w_eco47063, w_eco47064, w_eco47065, w_eco47066, w_eco47067, w_eco47068, w_eco47069, w_eco47070, w_eco47071, w_eco47072, w_eco47073, w_eco47074, w_eco47075, w_eco47076, w_eco47077, w_eco47078, w_eco47079, w_eco47080, w_eco47081, w_eco47082, w_eco47083, w_eco47084, w_eco47085, w_eco47086, w_eco47087, w_eco47088, w_eco47089, w_eco47090, w_eco47091, w_eco47092, w_eco47093, w_eco47094, w_eco47095, w_eco47096, w_eco47097, w_eco47098, w_eco47099, w_eco47100, w_eco47101, w_eco47102, w_eco47103, w_eco47104, w_eco47105, w_eco47106, w_eco47107, w_eco47108, w_eco47109, w_eco47110, w_eco47111, w_eco47112, w_eco47113, w_eco47114, w_eco47115, w_eco47116, w_eco47117, w_eco47118, w_eco47119, w_eco47120, w_eco47121, w_eco47122, w_eco47123, w_eco47124, w_eco47125, w_eco47126, w_eco47127, w_eco47128, w_eco47129, w_eco47130, w_eco47131, w_eco47132, w_eco47133, w_eco47134, w_eco47135, w_eco47136, w_eco47137, w_eco47138, w_eco47139, w_eco47140, w_eco47141, w_eco47142, w_eco47143, w_eco47144, w_eco47145, w_eco47146, w_eco47147, w_eco47148, w_eco47149, w_eco47150, w_eco47151, w_eco47152, w_eco47153, w_eco47154, w_eco47155, w_eco47156, w_eco47157, w_eco47158, w_eco47159, w_eco47160, w_eco47161, w_eco47162, w_eco47163, w_eco47164, w_eco47165, w_eco47166, w_eco47167, w_eco47168, w_eco47169, w_eco47170, w_eco47171, w_eco47172, w_eco47173, w_eco47174, w_eco47175, w_eco47176, w_eco47177, w_eco47178, w_eco47179, w_eco47180, w_eco47181, w_eco47182, w_eco47183, w_eco47184, w_eco47185, w_eco47186, w_eco47187, w_eco47188, w_eco47189, w_eco47190, w_eco47191, w_eco47192, w_eco47193, w_eco47194, w_eco47195, w_eco47196, w_eco47197, w_eco47198, w_eco47199, w_eco47200, w_eco47201, w_eco47202, w_eco47203, w_eco47204, w_eco47205, w_eco47206, w_eco47207, w_eco47208, w_eco47209, w_eco47210, w_eco47211, w_eco47212, w_eco47213, w_eco47214, w_eco47215, w_eco47216, w_eco47217, w_eco47218, w_eco47219, w_eco47220, w_eco47221, w_eco47222, w_eco47223, w_eco47224, w_eco47225, w_eco47226, w_eco47227, w_eco47228, w_eco47229, w_eco47230, w_eco47231, w_eco47232, w_eco47233, w_eco47234, w_eco47235, w_eco47236, w_eco47237, w_eco47238, w_eco47239, w_eco47240, w_eco47241, w_eco47242, w_eco47243, w_eco47244, w_eco47245, w_eco47246, w_eco47247, w_eco47248, w_eco47249, w_eco47250, w_eco47251, w_eco47252, w_eco47253, w_eco47254, w_eco47255, w_eco47256, w_eco47257, w_eco47258, w_eco47259, w_eco47260, w_eco47261, w_eco47262, w_eco47263, w_eco47264, w_eco47265, w_eco47266, w_eco47267, w_eco47268, w_eco47269, w_eco47270, w_eco47271, w_eco47272, w_eco47273, w_eco47274, w_eco47275, w_eco47276, w_eco47277, w_eco47278, w_eco47279, w_eco47280, w_eco47281, w_eco47282, w_eco47283, w_eco47284, w_eco47285, w_eco47286, w_eco47287, w_eco47288, w_eco47289, w_eco47290, w_eco47291, w_eco47292, w_eco47293, w_eco47294, w_eco47295, w_eco47296, w_eco47297, w_eco47298, w_eco47299, w_eco47300, w_eco47301, w_eco47302, w_eco47303, w_eco47304, w_eco47305, w_eco47306, w_eco47307, w_eco47308, w_eco47309, w_eco47310, w_eco47311, w_eco47312, w_eco47313, w_eco47314, w_eco47315, w_eco47316, w_eco47317, w_eco47318, w_eco47319, w_eco47320, w_eco47321, w_eco47322, w_eco47323, w_eco47324, w_eco47325, w_eco47326, w_eco47327, w_eco47328, w_eco47329, w_eco47330, w_eco47331, w_eco47332, w_eco47333, w_eco47334, w_eco47335, w_eco47336, w_eco47337, w_eco47338, w_eco47339, w_eco47340, w_eco47341, w_eco47342, w_eco47343, w_eco47344, w_eco47345, w_eco47346, w_eco47347, w_eco47348, w_eco47349, w_eco47350, w_eco47351, w_eco47352, w_eco47353, w_eco47354, w_eco47355, w_eco47356, w_eco47357, w_eco47358, w_eco47359, w_eco47360, w_eco47361, w_eco47362, w_eco47363, w_eco47364, w_eco47365, w_eco47366, w_eco47367, w_eco47368, w_eco47369, w_eco47370, w_eco47371, w_eco47372, w_eco47373, w_eco47374, w_eco47375, w_eco47376, w_eco47377, w_eco47378, w_eco47379, w_eco47380, w_eco47381, w_eco47382, w_eco47383, w_eco47384, w_eco47385, w_eco47386, w_eco47387, w_eco47388, w_eco47389, w_eco47390, w_eco47391, w_eco47392, w_eco47393, w_eco47394, w_eco47395, w_eco47396, w_eco47397, w_eco47398, w_eco47399, w_eco47400, w_eco47401, w_eco47402, w_eco47403, w_eco47404, w_eco47405, w_eco47406, w_eco47407, w_eco47408, w_eco47409, w_eco47410, w_eco47411, w_eco47412, w_eco47413, w_eco47414, w_eco47415, w_eco47416, w_eco47417, w_eco47418, w_eco47419, w_eco47420, w_eco47421, w_eco47422, w_eco47423, w_eco47424, w_eco47425, w_eco47426, w_eco47427, w_eco47428, w_eco47429, w_eco47430, w_eco47431, w_eco47432, w_eco47433, w_eco47434, w_eco47435, w_eco47436, w_eco47437, w_eco47438, w_eco47439, w_eco47440, w_eco47441, w_eco47442, w_eco47443, w_eco47444, w_eco47445, w_eco47446, w_eco47447, w_eco47448, w_eco47449, w_eco47450, w_eco47451, w_eco47452, w_eco47453, w_eco47454, w_eco47455, w_eco47456, w_eco47457, w_eco47458, w_eco47459, w_eco47460, w_eco47461, w_eco47462, w_eco47463, w_eco47464, w_eco47465, w_eco47466, w_eco47467, w_eco47468, w_eco47469, w_eco47470, w_eco47471, w_eco47472, w_eco47473, w_eco47474, w_eco47475, w_eco47476, w_eco47477, w_eco47478, w_eco47479, w_eco47480, w_eco47481, w_eco47482, w_eco47483, w_eco47484, w_eco47485, w_eco47486, w_eco47487, w_eco47488, w_eco47489, w_eco47490, w_eco47491, w_eco47492, w_eco47493, w_eco47494, w_eco47495, w_eco47496, w_eco47497, w_eco47498, w_eco47499, w_eco47500, w_eco47501, w_eco47502, w_eco47503, w_eco47504, w_eco47505, w_eco47506, w_eco47507, w_eco47508, w_eco47509, w_eco47510, w_eco47511, w_eco47512, w_eco47513, w_eco47514, w_eco47515, w_eco47516, w_eco47517, w_eco47518, w_eco47519, w_eco47520, w_eco47521, w_eco47522, w_eco47523, w_eco47524, w_eco47525, w_eco47526, w_eco47527, w_eco47528, w_eco47529, w_eco47530, w_eco47531, w_eco47532, w_eco47533, w_eco47534, w_eco47535, w_eco47536, w_eco47537, w_eco47538, w_eco47539, w_eco47540, w_eco47541, w_eco47542, w_eco47543, w_eco47544, w_eco47545, w_eco47546, w_eco47547, w_eco47548, w_eco47549, w_eco47550, w_eco47551, w_eco47552, w_eco47553, w_eco47554, w_eco47555, w_eco47556, w_eco47557, w_eco47558, w_eco47559, w_eco47560, w_eco47561, w_eco47562, w_eco47563, w_eco47564, w_eco47565, w_eco47566, w_eco47567, w_eco47568, w_eco47569, w_eco47570, w_eco47571, w_eco47572, w_eco47573, w_eco47574, w_eco47575, w_eco47576, w_eco47577, w_eco47578, w_eco47579, w_eco47580, w_eco47581, w_eco47582, w_eco47583, w_eco47584, w_eco47585, w_eco47586, w_eco47587, w_eco47588, w_eco47589, w_eco47590, w_eco47591, w_eco47592, w_eco47593, w_eco47594, w_eco47595, w_eco47596, w_eco47597, w_eco47598, w_eco47599, w_eco47600, w_eco47601, w_eco47602, w_eco47603, w_eco47604, w_eco47605, w_eco47606, w_eco47607, w_eco47608, w_eco47609, w_eco47610, w_eco47611, w_eco47612, w_eco47613, w_eco47614, w_eco47615, w_eco47616, w_eco47617, w_eco47618, w_eco47619, w_eco47620, w_eco47621, w_eco47622, w_eco47623, w_eco47624, w_eco47625, w_eco47626, w_eco47627, w_eco47628, w_eco47629, w_eco47630, w_eco47631, w_eco47632, w_eco47633, w_eco47634, w_eco47635, w_eco47636, w_eco47637, w_eco47638, w_eco47639, w_eco47640, w_eco47641, w_eco47642, w_eco47643, w_eco47644, w_eco47645, w_eco47646, w_eco47647, w_eco47648, w_eco47649, w_eco47650, w_eco47651, w_eco47652, w_eco47653, w_eco47654, w_eco47655, w_eco47656, w_eco47657, w_eco47658, w_eco47659, w_eco47660, w_eco47661, w_eco47662, w_eco47663, w_eco47664, w_eco47665, w_eco47666, w_eco47667, w_eco47668, w_eco47669, w_eco47670, w_eco47671, w_eco47672, w_eco47673, w_eco47674, w_eco47675, w_eco47676, w_eco47677, w_eco47678, w_eco47679, w_eco47680, w_eco47681, w_eco47682, w_eco47683, w_eco47684, w_eco47685, w_eco47686, w_eco47687, w_eco47688, w_eco47689, w_eco47690, w_eco47691, w_eco47692, w_eco47693, w_eco47694, w_eco47695, w_eco47696, w_eco47697, w_eco47698, w_eco47699, w_eco47700, w_eco47701, w_eco47702, w_eco47703, w_eco47704, w_eco47705, w_eco47706, w_eco47707, w_eco47708, w_eco47709, w_eco47710, w_eco47711, w_eco47712, w_eco47713, w_eco47714, w_eco47715, w_eco47716, w_eco47717, w_eco47718, w_eco47719, w_eco47720, w_eco47721, w_eco47722, w_eco47723, w_eco47724, w_eco47725, w_eco47726, w_eco47727, w_eco47728, w_eco47729, w_eco47730, w_eco47731, w_eco47732, w_eco47733, w_eco47734, w_eco47735, w_eco47736, w_eco47737, w_eco47738, w_eco47739, w_eco47740, w_eco47741, w_eco47742, w_eco47743, w_eco47744, w_eco47745, w_eco47746, w_eco47747, w_eco47748, w_eco47749, w_eco47750, w_eco47751, w_eco47752, w_eco47753, w_eco47754, w_eco47755, w_eco47756, w_eco47757, w_eco47758, w_eco47759, w_eco47760, w_eco47761, w_eco47762, w_eco47763, w_eco47764, w_eco47765, w_eco47766, w_eco47767, w_eco47768, w_eco47769, w_eco47770, w_eco47771, w_eco47772, w_eco47773, w_eco47774, w_eco47775, w_eco47776, w_eco47777, w_eco47778, w_eco47779, w_eco47780, w_eco47781, w_eco47782, w_eco47783, w_eco47784, w_eco47785, w_eco47786, w_eco47787, w_eco47788, w_eco47789, w_eco47790, w_eco47791, w_eco47792, w_eco47793, w_eco47794, w_eco47795, w_eco47796, w_eco47797, w_eco47798, w_eco47799, w_eco47800, w_eco47801, w_eco47802, w_eco47803, w_eco47804, w_eco47805, w_eco47806, w_eco47807, w_eco47808, w_eco47809, w_eco47810, w_eco47811, w_eco47812, w_eco47813, w_eco47814, w_eco47815, w_eco47816, w_eco47817, w_eco47818, w_eco47819, w_eco47820, w_eco47821, w_eco47822, w_eco47823, w_eco47824, w_eco47825, w_eco47826, w_eco47827, w_eco47828, w_eco47829, w_eco47830, w_eco47831, w_eco47832, w_eco47833, w_eco47834, w_eco47835, w_eco47836, w_eco47837, w_eco47838, w_eco47839, w_eco47840, w_eco47841, w_eco47842, w_eco47843, w_eco47844, w_eco47845, w_eco47846, w_eco47847, w_eco47848, w_eco47849, w_eco47850, w_eco47851, w_eco47852, w_eco47853, w_eco47854, w_eco47855, w_eco47856, w_eco47857, w_eco47858, w_eco47859, w_eco47860, w_eco47861, w_eco47862, w_eco47863, w_eco47864, w_eco47865, w_eco47866, w_eco47867, w_eco47868, w_eco47869, w_eco47870, w_eco47871, w_eco47872, w_eco47873, w_eco47874, w_eco47875, w_eco47876, w_eco47877, w_eco47878, w_eco47879, w_eco47880, w_eco47881, w_eco47882, w_eco47883, w_eco47884, w_eco47885, w_eco47886, w_eco47887, w_eco47888, w_eco47889, w_eco47890, w_eco47891, w_eco47892, w_eco47893, w_eco47894, w_eco47895, w_eco47896, w_eco47897, w_eco47898, w_eco47899, w_eco47900, w_eco47901, w_eco47902, w_eco47903, w_eco47904, w_eco47905, w_eco47906, w_eco47907, w_eco47908, w_eco47909, w_eco47910, w_eco47911, w_eco47912, w_eco47913, w_eco47914, w_eco47915, w_eco47916, w_eco47917, w_eco47918, w_eco47919, w_eco47920, w_eco47921, w_eco47922, w_eco47923, w_eco47924, w_eco47925, w_eco47926, w_eco47927, w_eco47928, w_eco47929, w_eco47930, w_eco47931, w_eco47932, w_eco47933, w_eco47934, w_eco47935, w_eco47936, w_eco47937, w_eco47938, w_eco47939, w_eco47940, w_eco47941, w_eco47942, w_eco47943, w_eco47944, w_eco47945, w_eco47946, w_eco47947, w_eco47948, w_eco47949, w_eco47950, w_eco47951, w_eco47952, w_eco47953, w_eco47954, w_eco47955, w_eco47956, w_eco47957, w_eco47958, w_eco47959, w_eco47960, w_eco47961, w_eco47962, w_eco47963, w_eco47964, w_eco47965, w_eco47966, w_eco47967, w_eco47968, w_eco47969, w_eco47970, w_eco47971, w_eco47972, w_eco47973, w_eco47974, w_eco47975, w_eco47976, w_eco47977, w_eco47978, w_eco47979, w_eco47980, w_eco47981, w_eco47982, w_eco47983, w_eco47984, w_eco47985, w_eco47986, w_eco47987, w_eco47988, w_eco47989, w_eco47990, w_eco47991, w_eco47992, w_eco47993, w_eco47994, w_eco47995, w_eco47996, w_eco47997, w_eco47998, w_eco47999, w_eco48000, w_eco48001, w_eco48002, w_eco48003, w_eco48004, w_eco48005, w_eco48006, w_eco48007, w_eco48008, w_eco48009, w_eco48010, w_eco48011, w_eco48012, w_eco48013, w_eco48014, w_eco48015, w_eco48016, w_eco48017, w_eco48018, w_eco48019, w_eco48020, w_eco48021, w_eco48022, w_eco48023, w_eco48024, w_eco48025, w_eco48026, w_eco48027, w_eco48028, w_eco48029, w_eco48030, w_eco48031, w_eco48032, w_eco48033, w_eco48034, w_eco48035, w_eco48036, w_eco48037, w_eco48038, w_eco48039, w_eco48040, w_eco48041, w_eco48042, w_eco48043, w_eco48044, w_eco48045, w_eco48046, w_eco48047, w_eco48048, w_eco48049, w_eco48050, w_eco48051, w_eco48052, w_eco48053, w_eco48054, w_eco48055, w_eco48056, w_eco48057, w_eco48058, w_eco48059, w_eco48060, w_eco48061, w_eco48062, w_eco48063, w_eco48064, w_eco48065, w_eco48066, w_eco48067, w_eco48068, w_eco48069, w_eco48070, w_eco48071, w_eco48072, w_eco48073, w_eco48074, w_eco48075, w_eco48076, w_eco48077, w_eco48078, w_eco48079, w_eco48080, w_eco48081, w_eco48082, w_eco48083, w_eco48084, w_eco48085, w_eco48086, w_eco48087, w_eco48088, w_eco48089, w_eco48090, w_eco48091, w_eco48092, w_eco48093, w_eco48094, w_eco48095, w_eco48096, w_eco48097, w_eco48098, w_eco48099, w_eco48100, w_eco48101, w_eco48102, w_eco48103, w_eco48104, w_eco48105, w_eco48106, w_eco48107, w_eco48108, w_eco48109, w_eco48110, w_eco48111, w_eco48112, w_eco48113, w_eco48114, w_eco48115, w_eco48116, w_eco48117, w_eco48118, w_eco48119, w_eco48120, w_eco48121, w_eco48122, w_eco48123, w_eco48124, w_eco48125, w_eco48126, w_eco48127, w_eco48128, w_eco48129, w_eco48130, w_eco48131, w_eco48132, w_eco48133, w_eco48134, w_eco48135, w_eco48136, w_eco48137, w_eco48138, w_eco48139, w_eco48140, w_eco48141, w_eco48142, w_eco48143, w_eco48144, w_eco48145, w_eco48146, w_eco48147, w_eco48148, w_eco48149, w_eco48150, w_eco48151, w_eco48152, w_eco48153, w_eco48154, w_eco48155, w_eco48156, w_eco48157, w_eco48158, w_eco48159, w_eco48160, w_eco48161, w_eco48162, w_eco48163, w_eco48164, w_eco48165, w_eco48166, w_eco48167, w_eco48168, w_eco48169, w_eco48170, w_eco48171, w_eco48172, w_eco48173, w_eco48174, w_eco48175, w_eco48176, w_eco48177, w_eco48178, w_eco48179, w_eco48180, w_eco48181, w_eco48182, w_eco48183, w_eco48184, w_eco48185, w_eco48186, w_eco48187, w_eco48188, w_eco48189, w_eco48190, w_eco48191, w_eco48192, w_eco48193, w_eco48194, w_eco48195, w_eco48196, w_eco48197, w_eco48198, w_eco48199, w_eco48200, w_eco48201, w_eco48202, w_eco48203, w_eco48204, w_eco48205, w_eco48206, w_eco48207, w_eco48208, w_eco48209, w_eco48210, w_eco48211, w_eco48212, w_eco48213, w_eco48214, w_eco48215, w_eco48216, w_eco48217, w_eco48218, w_eco48219, w_eco48220, w_eco48221, w_eco48222, w_eco48223, w_eco48224, w_eco48225, w_eco48226, w_eco48227, w_eco48228, w_eco48229, w_eco48230, w_eco48231, w_eco48232, w_eco48233, w_eco48234, w_eco48235, w_eco48236, w_eco48237, w_eco48238, w_eco48239, w_eco48240, w_eco48241, w_eco48242, w_eco48243, w_eco48244, w_eco48245, w_eco48246, w_eco48247, w_eco48248, w_eco48249, w_eco48250, w_eco48251, w_eco48252, w_eco48253, w_eco48254, w_eco48255, w_eco48256, w_eco48257, w_eco48258, w_eco48259, w_eco48260, w_eco48261, w_eco48262, w_eco48263, w_eco48264, w_eco48265, w_eco48266, w_eco48267, w_eco48268, w_eco48269, w_eco48270, w_eco48271, w_eco48272, w_eco48273, w_eco48274, w_eco48275, w_eco48276, w_eco48277, w_eco48278, w_eco48279, w_eco48280, w_eco48281, w_eco48282, w_eco48283, w_eco48284, w_eco48285, w_eco48286, w_eco48287, w_eco48288, w_eco48289, w_eco48290, w_eco48291, w_eco48292, w_eco48293, w_eco48294, w_eco48295, w_eco48296, w_eco48297, w_eco48298, w_eco48299, w_eco48300, w_eco48301, w_eco48302, w_eco48303, w_eco48304, w_eco48305, w_eco48306, w_eco48307, w_eco48308, w_eco48309, w_eco48310, w_eco48311, w_eco48312, w_eco48313, w_eco48314, w_eco48315, w_eco48316, w_eco48317, w_eco48318, w_eco48319, w_eco48320, w_eco48321, w_eco48322, w_eco48323, w_eco48324, w_eco48325, w_eco48326, w_eco48327, w_eco48328, w_eco48329, w_eco48330, w_eco48331, w_eco48332, w_eco48333, w_eco48334, w_eco48335, w_eco48336, w_eco48337, w_eco48338, w_eco48339, w_eco48340, w_eco48341, w_eco48342, w_eco48343, w_eco48344, w_eco48345, w_eco48346, w_eco48347, w_eco48348, w_eco48349, w_eco48350, w_eco48351, w_eco48352, w_eco48353, w_eco48354, w_eco48355, w_eco48356, w_eco48357, w_eco48358, w_eco48359, w_eco48360, w_eco48361, w_eco48362, w_eco48363, w_eco48364, w_eco48365, w_eco48366, w_eco48367, w_eco48368, w_eco48369, w_eco48370, w_eco48371, w_eco48372, w_eco48373, w_eco48374, w_eco48375, w_eco48376, w_eco48377, w_eco48378, w_eco48379, w_eco48380, w_eco48381, w_eco48382, w_eco48383, w_eco48384, w_eco48385, w_eco48386, w_eco48387, w_eco48388, w_eco48389, w_eco48390, w_eco48391, w_eco48392, w_eco48393, w_eco48394, w_eco48395, w_eco48396, w_eco48397, w_eco48398, w_eco48399, w_eco48400, w_eco48401, w_eco48402, w_eco48403, w_eco48404, w_eco48405, w_eco48406, w_eco48407, w_eco48408, w_eco48409, w_eco48410, w_eco48411, w_eco48412, w_eco48413, w_eco48414, w_eco48415, w_eco48416, w_eco48417, w_eco48418, w_eco48419, w_eco48420, w_eco48421, w_eco48422, w_eco48423, w_eco48424, w_eco48425, w_eco48426, w_eco48427, w_eco48428, w_eco48429, w_eco48430, w_eco48431, w_eco48432, w_eco48433, w_eco48434, w_eco48435, w_eco48436, w_eco48437, w_eco48438, w_eco48439, w_eco48440, w_eco48441, w_eco48442, w_eco48443, w_eco48444, w_eco48445, w_eco48446, w_eco48447, w_eco48448, w_eco48449, w_eco48450, w_eco48451, w_eco48452, w_eco48453, w_eco48454, w_eco48455, w_eco48456, w_eco48457, w_eco48458, w_eco48459, w_eco48460, w_eco48461, w_eco48462, w_eco48463, w_eco48464, w_eco48465, w_eco48466, w_eco48467, w_eco48468, w_eco48469, w_eco48470, w_eco48471, w_eco48472, w_eco48473, w_eco48474, w_eco48475, w_eco48476, w_eco48477, w_eco48478, w_eco48479, w_eco48480, w_eco48481, w_eco48482, w_eco48483, w_eco48484, w_eco48485, w_eco48486, w_eco48487, w_eco48488, w_eco48489, w_eco48490, w_eco48491, w_eco48492, w_eco48493, w_eco48494, w_eco48495, w_eco48496, w_eco48497, w_eco48498, w_eco48499, w_eco48500, w_eco48501, w_eco48502, w_eco48503, w_eco48504, w_eco48505, w_eco48506, w_eco48507, w_eco48508, w_eco48509, w_eco48510, w_eco48511, w_eco48512, w_eco48513, w_eco48514, w_eco48515, w_eco48516, w_eco48517, w_eco48518, w_eco48519, w_eco48520, w_eco48521, w_eco48522, w_eco48523, w_eco48524, w_eco48525, w_eco48526, w_eco48527, w_eco48528, w_eco48529, w_eco48530, w_eco48531, w_eco48532, w_eco48533, w_eco48534, w_eco48535, w_eco48536, w_eco48537, w_eco48538, w_eco48539, w_eco48540, w_eco48541, w_eco48542, w_eco48543, w_eco48544, w_eco48545, w_eco48546, w_eco48547, w_eco48548, w_eco48549, w_eco48550, w_eco48551, w_eco48552, w_eco48553, w_eco48554, w_eco48555, w_eco48556, w_eco48557, w_eco48558, w_eco48559, w_eco48560, w_eco48561, w_eco48562, w_eco48563, w_eco48564, w_eco48565, w_eco48566, w_eco48567, w_eco48568, w_eco48569, w_eco48570, w_eco48571, w_eco48572, w_eco48573, w_eco48574, w_eco48575, w_eco48576, w_eco48577, w_eco48578, w_eco48579, w_eco48580, w_eco48581, w_eco48582, w_eco48583, w_eco48584, w_eco48585, w_eco48586, w_eco48587, w_eco48588, w_eco48589, w_eco48590, w_eco48591, w_eco48592, w_eco48593, w_eco48594, w_eco48595, w_eco48596, w_eco48597, w_eco48598, w_eco48599, w_eco48600, w_eco48601, w_eco48602, w_eco48603, w_eco48604, w_eco48605, w_eco48606, w_eco48607, w_eco48608, w_eco48609, w_eco48610, w_eco48611, w_eco48612, w_eco48613, w_eco48614, w_eco48615, w_eco48616, w_eco48617, w_eco48618, w_eco48619, w_eco48620, w_eco48621, w_eco48622, w_eco48623, w_eco48624, w_eco48625, w_eco48626, w_eco48627, w_eco48628, w_eco48629, w_eco48630, w_eco48631, w_eco48632, w_eco48633, w_eco48634, w_eco48635, w_eco48636, w_eco48637, w_eco48638, w_eco48639, w_eco48640, w_eco48641, w_eco48642, w_eco48643, w_eco48644, w_eco48645, w_eco48646, w_eco48647, w_eco48648, w_eco48649, w_eco48650, w_eco48651, w_eco48652, w_eco48653, w_eco48654, w_eco48655, w_eco48656, w_eco48657, w_eco48658, w_eco48659, w_eco48660, w_eco48661, w_eco48662, w_eco48663, w_eco48664, w_eco48665, w_eco48666, w_eco48667, w_eco48668, w_eco48669, w_eco48670, w_eco48671, w_eco48672, w_eco48673, w_eco48674, w_eco48675, w_eco48676, w_eco48677, w_eco48678, w_eco48679, w_eco48680, w_eco48681, w_eco48682, w_eco48683, w_eco48684, w_eco48685, w_eco48686, w_eco48687, w_eco48688, w_eco48689, w_eco48690, w_eco48691, w_eco48692, w_eco48693, w_eco48694, w_eco48695, w_eco48696, w_eco48697, w_eco48698, w_eco48699, w_eco48700, w_eco48701, w_eco48702, w_eco48703, w_eco48704, w_eco48705, w_eco48706, w_eco48707, w_eco48708, w_eco48709, w_eco48710, w_eco48711, w_eco48712, w_eco48713, w_eco48714, w_eco48715, w_eco48716, w_eco48717, w_eco48718, w_eco48719, w_eco48720, w_eco48721, w_eco48722, w_eco48723, w_eco48724, w_eco48725, w_eco48726, w_eco48727, w_eco48728, w_eco48729, w_eco48730, w_eco48731, w_eco48732, w_eco48733, w_eco48734, w_eco48735, w_eco48736, w_eco48737, w_eco48738, w_eco48739, w_eco48740, w_eco48741, w_eco48742, w_eco48743, w_eco48744, w_eco48745, w_eco48746, w_eco48747, w_eco48748, w_eco48749, w_eco48750, w_eco48751, w_eco48752, w_eco48753, w_eco48754, w_eco48755, w_eco48756, w_eco48757, w_eco48758, w_eco48759, w_eco48760, w_eco48761, w_eco48762, w_eco48763, w_eco48764, w_eco48765, w_eco48766, w_eco48767, w_eco48768, w_eco48769, w_eco48770, w_eco48771, w_eco48772, w_eco48773, w_eco48774, w_eco48775, w_eco48776, w_eco48777, w_eco48778, w_eco48779, w_eco48780, w_eco48781, w_eco48782, w_eco48783, w_eco48784, w_eco48785, w_eco48786, w_eco48787, w_eco48788, w_eco48789, w_eco48790, w_eco48791, w_eco48792, w_eco48793, w_eco48794, w_eco48795, w_eco48796, w_eco48797, w_eco48798, w_eco48799, w_eco48800, w_eco48801, w_eco48802, w_eco48803, w_eco48804, w_eco48805, w_eco48806, w_eco48807, w_eco48808, w_eco48809, w_eco48810, w_eco48811, w_eco48812, w_eco48813, w_eco48814, w_eco48815, w_eco48816, w_eco48817, w_eco48818, w_eco48819, w_eco48820, w_eco48821, w_eco48822, w_eco48823, w_eco48824, w_eco48825, w_eco48826, w_eco48827, w_eco48828, w_eco48829, w_eco48830, w_eco48831, w_eco48832, w_eco48833, w_eco48834, w_eco48835, w_eco48836, w_eco48837, w_eco48838, w_eco48839, w_eco48840, w_eco48841, w_eco48842, w_eco48843, w_eco48844, w_eco48845, w_eco48846, w_eco48847, w_eco48848, w_eco48849, w_eco48850, w_eco48851, w_eco48852, w_eco48853, w_eco48854, w_eco48855, w_eco48856, w_eco48857, w_eco48858, w_eco48859, w_eco48860, w_eco48861, w_eco48862, w_eco48863, w_eco48864, w_eco48865, w_eco48866, w_eco48867, w_eco48868, w_eco48869, w_eco48870, w_eco48871, w_eco48872, w_eco48873, w_eco48874, w_eco48875, w_eco48876, w_eco48877, w_eco48878, w_eco48879, w_eco48880, w_eco48881, w_eco48882, w_eco48883, w_eco48884, w_eco48885, w_eco48886, w_eco48887, w_eco48888, w_eco48889, w_eco48890, w_eco48891, w_eco48892, w_eco48893, w_eco48894, w_eco48895, w_eco48896, w_eco48897, w_eco48898, w_eco48899, w_eco48900, w_eco48901, w_eco48902, w_eco48903, w_eco48904, w_eco48905, w_eco48906, w_eco48907, w_eco48908, w_eco48909, w_eco48910, w_eco48911, w_eco48912, w_eco48913, w_eco48914, w_eco48915, w_eco48916, w_eco48917, w_eco48918, w_eco48919, w_eco48920, w_eco48921, w_eco48922, w_eco48923, w_eco48924, w_eco48925, w_eco48926, w_eco48927, w_eco48928, w_eco48929, w_eco48930, w_eco48931, w_eco48932, w_eco48933, w_eco48934, w_eco48935, w_eco48936, w_eco48937, w_eco48938, w_eco48939, w_eco48940, w_eco48941, w_eco48942, w_eco48943, w_eco48944, w_eco48945, w_eco48946, w_eco48947, w_eco48948, w_eco48949, w_eco48950, w_eco48951, w_eco48952, w_eco48953, w_eco48954, w_eco48955, w_eco48956, w_eco48957, w_eco48958, w_eco48959, w_eco48960, w_eco48961, w_eco48962, w_eco48963, w_eco48964, w_eco48965, w_eco48966, w_eco48967, w_eco48968, w_eco48969, w_eco48970, w_eco48971, w_eco48972, w_eco48973, w_eco48974, w_eco48975, w_eco48976, w_eco48977, w_eco48978, w_eco48979, w_eco48980, w_eco48981, w_eco48982, w_eco48983, w_eco48984, w_eco48985, w_eco48986, w_eco48987, w_eco48988, w_eco48989, w_eco48990, w_eco48991, w_eco48992, w_eco48993, w_eco48994, w_eco48995, w_eco48996, w_eco48997, w_eco48998, w_eco48999, w_eco49000, w_eco49001, w_eco49002, w_eco49003, w_eco49004, w_eco49005, w_eco49006, w_eco49007, w_eco49008, w_eco49009, w_eco49010, w_eco49011, w_eco49012, w_eco49013, w_eco49014, w_eco49015, w_eco49016, w_eco49017, w_eco49018, w_eco49019, w_eco49020, w_eco49021, w_eco49022, w_eco49023, w_eco49024, w_eco49025, w_eco49026, w_eco49027, w_eco49028, w_eco49029, w_eco49030, w_eco49031, w_eco49032, w_eco49033, w_eco49034, w_eco49035, w_eco49036, w_eco49037, w_eco49038, w_eco49039, w_eco49040, w_eco49041, w_eco49042, w_eco49043, w_eco49044, w_eco49045, w_eco49046, w_eco49047, w_eco49048, w_eco49049, w_eco49050, w_eco49051, w_eco49052, w_eco49053, w_eco49054, w_eco49055, w_eco49056, w_eco49057, w_eco49058, w_eco49059, w_eco49060, w_eco49061, w_eco49062, w_eco49063, w_eco49064, w_eco49065, w_eco49066, w_eco49067, w_eco49068, w_eco49069, w_eco49070, w_eco49071, w_eco49072, w_eco49073, w_eco49074, w_eco49075, w_eco49076, w_eco49077, w_eco49078, w_eco49079, w_eco49080, w_eco49081, w_eco49082, w_eco49083, w_eco49084, w_eco49085, w_eco49086, w_eco49087, w_eco49088, w_eco49089, w_eco49090, w_eco49091, w_eco49092, w_eco49093, w_eco49094, w_eco49095, w_eco49096, w_eco49097, w_eco49098, w_eco49099, w_eco49100, w_eco49101, w_eco49102, w_eco49103, w_eco49104, w_eco49105, w_eco49106, w_eco49107, w_eco49108, w_eco49109, w_eco49110, w_eco49111, w_eco49112, w_eco49113, w_eco49114, w_eco49115, w_eco49116, w_eco49117, w_eco49118, w_eco49119, w_eco49120, w_eco49121, w_eco49122, w_eco49123, w_eco49124, w_eco49125, w_eco49126, w_eco49127, w_eco49128, w_eco49129, w_eco49130, w_eco49131, w_eco49132, w_eco49133, w_eco49134, w_eco49135, w_eco49136, w_eco49137, w_eco49138, w_eco49139, w_eco49140, w_eco49141, w_eco49142, w_eco49143, w_eco49144, w_eco49145, w_eco49146, w_eco49147, w_eco49148, w_eco49149, w_eco49150, w_eco49151, w_eco49152, w_eco49153, w_eco49154, w_eco49155, w_eco49156, w_eco49157, w_eco49158, w_eco49159, w_eco49160, w_eco49161, w_eco49162, w_eco49163, w_eco49164, w_eco49165, w_eco49166, w_eco49167, w_eco49168, w_eco49169, w_eco49170, w_eco49171, w_eco49172, w_eco49173, w_eco49174, w_eco49175, w_eco49176, w_eco49177, w_eco49178, w_eco49179, w_eco49180, w_eco49181, w_eco49182, w_eco49183, w_eco49184, w_eco49185, w_eco49186, w_eco49187, w_eco49188, w_eco49189, w_eco49190, w_eco49191, w_eco49192, w_eco49193, w_eco49194, w_eco49195, w_eco49196, w_eco49197, w_eco49198, w_eco49199, w_eco49200, w_eco49201, w_eco49202, w_eco49203, w_eco49204, w_eco49205, w_eco49206, w_eco49207, w_eco49208, w_eco49209, w_eco49210, w_eco49211, w_eco49212, w_eco49213, w_eco49214, w_eco49215, w_eco49216, w_eco49217, w_eco49218, w_eco49219, w_eco49220, w_eco49221, w_eco49222, w_eco49223, w_eco49224, w_eco49225, w_eco49226, w_eco49227, w_eco49228, w_eco49229, w_eco49230, w_eco49231, w_eco49232, w_eco49233, w_eco49234, w_eco49235, w_eco49236, w_eco49237, w_eco49238, w_eco49239, w_eco49240, w_eco49241, w_eco49242, w_eco49243, w_eco49244, w_eco49245, w_eco49246, w_eco49247, w_eco49248, w_eco49249, w_eco49250, w_eco49251, w_eco49252, w_eco49253, w_eco49254, w_eco49255, w_eco49256, w_eco49257, w_eco49258, w_eco49259, w_eco49260, w_eco49261, w_eco49262, w_eco49263, w_eco49264, w_eco49265, w_eco49266, w_eco49267, w_eco49268, w_eco49269, w_eco49270, w_eco49271, w_eco49272, w_eco49273, w_eco49274, w_eco49275, w_eco49276, w_eco49277, w_eco49278, w_eco49279, w_eco49280, w_eco49281, w_eco49282, w_eco49283, w_eco49284, w_eco49285, w_eco49286, w_eco49287, w_eco49288, w_eco49289, w_eco49290, w_eco49291, w_eco49292, w_eco49293, w_eco49294, w_eco49295, w_eco49296, w_eco49297, w_eco49298, w_eco49299, w_eco49300, w_eco49301, w_eco49302, w_eco49303, w_eco49304, w_eco49305, w_eco49306, w_eco49307, w_eco49308, w_eco49309, w_eco49310, w_eco49311, w_eco49312, w_eco49313, w_eco49314, w_eco49315, w_eco49316, w_eco49317, w_eco49318, w_eco49319, w_eco49320, w_eco49321, w_eco49322, w_eco49323, w_eco49324, w_eco49325, w_eco49326, w_eco49327, w_eco49328, w_eco49329, w_eco49330, w_eco49331, w_eco49332, w_eco49333, w_eco49334, w_eco49335, w_eco49336, w_eco49337, w_eco49338, w_eco49339, w_eco49340, w_eco49341, w_eco49342, w_eco49343, w_eco49344, w_eco49345, w_eco49346, w_eco49347, w_eco49348, w_eco49349, w_eco49350, w_eco49351, w_eco49352, w_eco49353, w_eco49354, w_eco49355, w_eco49356, w_eco49357, w_eco49358, w_eco49359, w_eco49360, w_eco49361, w_eco49362, w_eco49363, w_eco49364, w_eco49365, w_eco49366, w_eco49367, w_eco49368, w_eco49369, w_eco49370, w_eco49371, w_eco49372, w_eco49373, w_eco49374, w_eco49375, w_eco49376, w_eco49377, w_eco49378, w_eco49379, w_eco49380, w_eco49381, w_eco49382, w_eco49383, w_eco49384, w_eco49385, w_eco49386, w_eco49387, w_eco49388, w_eco49389, w_eco49390, w_eco49391, w_eco49392, w_eco49393, w_eco49394, w_eco49395, w_eco49396, w_eco49397, w_eco49398, w_eco49399, w_eco49400, w_eco49401, w_eco49402, w_eco49403, w_eco49404, w_eco49405, w_eco49406, w_eco49407, w_eco49408, w_eco49409, w_eco49410, w_eco49411, w_eco49412, w_eco49413, w_eco49414, w_eco49415, w_eco49416, w_eco49417, w_eco49418, w_eco49419, w_eco49420, w_eco49421, w_eco49422, w_eco49423, w_eco49424, w_eco49425, w_eco49426, w_eco49427, w_eco49428, w_eco49429, w_eco49430, w_eco49431, w_eco49432, w_eco49433, w_eco49434, w_eco49435, w_eco49436, w_eco49437, w_eco49438, w_eco49439, w_eco49440, w_eco49441, w_eco49442, w_eco49443, w_eco49444, w_eco49445, w_eco49446, w_eco49447, w_eco49448, w_eco49449, w_eco49450, w_eco49451, w_eco49452, w_eco49453, w_eco49454, w_eco49455, w_eco49456, w_eco49457, w_eco49458, w_eco49459, w_eco49460, w_eco49461, w_eco49462, w_eco49463, w_eco49464, w_eco49465, w_eco49466, w_eco49467, w_eco49468, w_eco49469, w_eco49470, w_eco49471, w_eco49472, w_eco49473, w_eco49474, w_eco49475, w_eco49476, w_eco49477, w_eco49478, w_eco49479, w_eco49480, w_eco49481, w_eco49482, w_eco49483, w_eco49484, w_eco49485, w_eco49486, w_eco49487, w_eco49488, w_eco49489, w_eco49490, w_eco49491, w_eco49492, w_eco49493, w_eco49494, w_eco49495, w_eco49496, w_eco49497, w_eco49498, w_eco49499, w_eco49500, w_eco49501, w_eco49502, w_eco49503, w_eco49504, w_eco49505, w_eco49506, w_eco49507, w_eco49508, w_eco49509, w_eco49510, w_eco49511, w_eco49512, w_eco49513, w_eco49514, w_eco49515, w_eco49516, w_eco49517, w_eco49518, w_eco49519, w_eco49520, w_eco49521, w_eco49522, w_eco49523, w_eco49524, w_eco49525, w_eco49526, w_eco49527, w_eco49528, w_eco49529, w_eco49530, w_eco49531, w_eco49532, w_eco49533, w_eco49534, w_eco49535, w_eco49536, w_eco49537, w_eco49538, w_eco49539, w_eco49540, w_eco49541, w_eco49542, w_eco49543, w_eco49544, w_eco49545, w_eco49546, w_eco49547, w_eco49548, w_eco49549, w_eco49550, w_eco49551, w_eco49552, w_eco49553, w_eco49554, w_eco49555, w_eco49556, w_eco49557, w_eco49558, w_eco49559, w_eco49560, w_eco49561, w_eco49562, w_eco49563, w_eco49564, w_eco49565, w_eco49566, w_eco49567, w_eco49568, w_eco49569, w_eco49570, w_eco49571, w_eco49572, w_eco49573, w_eco49574, w_eco49575, w_eco49576, w_eco49577, w_eco49578, w_eco49579, w_eco49580, w_eco49581, w_eco49582, w_eco49583, w_eco49584, w_eco49585, w_eco49586, w_eco49587, w_eco49588, w_eco49589, w_eco49590, w_eco49591, w_eco49592, w_eco49593, w_eco49594, w_eco49595, w_eco49596, w_eco49597, w_eco49598, w_eco49599, w_eco49600, w_eco49601, w_eco49602, w_eco49603, w_eco49604, w_eco49605, w_eco49606, w_eco49607, w_eco49608, w_eco49609, w_eco49610, w_eco49611, w_eco49612, w_eco49613, w_eco49614, w_eco49615, w_eco49616, w_eco49617, w_eco49618, w_eco49619, w_eco49620, w_eco49621, w_eco49622, w_eco49623, w_eco49624, w_eco49625, w_eco49626, w_eco49627, w_eco49628, w_eco49629, w_eco49630, w_eco49631, w_eco49632, w_eco49633, w_eco49634, w_eco49635, w_eco49636, w_eco49637, w_eco49638, w_eco49639, w_eco49640, w_eco49641, w_eco49642, w_eco49643, w_eco49644, w_eco49645, w_eco49646, w_eco49647, w_eco49648, w_eco49649, w_eco49650, w_eco49651, w_eco49652, w_eco49653, w_eco49654, w_eco49655, w_eco49656, w_eco49657, w_eco49658, w_eco49659, w_eco49660, w_eco49661, w_eco49662, w_eco49663, w_eco49664, w_eco49665, w_eco49666, w_eco49667, w_eco49668, w_eco49669, w_eco49670, w_eco49671, w_eco49672, w_eco49673, w_eco49674, w_eco49675, w_eco49676, w_eco49677, w_eco49678, w_eco49679, w_eco49680, w_eco49681, w_eco49682, w_eco49683, w_eco49684, w_eco49685, w_eco49686, w_eco49687, w_eco49688, w_eco49689, w_eco49690, w_eco49691, w_eco49692, w_eco49693, w_eco49694, w_eco49695, w_eco49696, w_eco49697, w_eco49698, w_eco49699, w_eco49700, w_eco49701, w_eco49702, w_eco49703, w_eco49704, w_eco49705, w_eco49706, w_eco49707, w_eco49708, w_eco49709, w_eco49710, w_eco49711, w_eco49712, w_eco49713, w_eco49714, w_eco49715, w_eco49716, w_eco49717, w_eco49718, w_eco49719, w_eco49720, w_eco49721, w_eco49722, w_eco49723, w_eco49724, w_eco49725, w_eco49726, w_eco49727, w_eco49728, w_eco49729, w_eco49730, w_eco49731, w_eco49732, w_eco49733, w_eco49734, w_eco49735, w_eco49736, w_eco49737, w_eco49738, w_eco49739, w_eco49740, w_eco49741, w_eco49742, w_eco49743, w_eco49744, w_eco49745, w_eco49746, w_eco49747, w_eco49748, w_eco49749, w_eco49750, w_eco49751, w_eco49752, w_eco49753, w_eco49754, w_eco49755, w_eco49756, w_eco49757, w_eco49758, w_eco49759, w_eco49760, w_eco49761, w_eco49762, w_eco49763, w_eco49764, w_eco49765, w_eco49766, w_eco49767, w_eco49768, w_eco49769, w_eco49770, w_eco49771, w_eco49772, w_eco49773, w_eco49774, w_eco49775, w_eco49776, w_eco49777, w_eco49778, w_eco49779, w_eco49780, w_eco49781, w_eco49782, w_eco49783, w_eco49784, w_eco49785, w_eco49786, w_eco49787, w_eco49788, w_eco49789, w_eco49790, w_eco49791, w_eco49792, w_eco49793, w_eco49794, w_eco49795, w_eco49796, w_eco49797, w_eco49798, w_eco49799, w_eco49800, w_eco49801, w_eco49802, w_eco49803, w_eco49804, w_eco49805, w_eco49806, w_eco49807, w_eco49808, w_eco49809, w_eco49810, w_eco49811, w_eco49812, w_eco49813, w_eco49814, w_eco49815, w_eco49816, w_eco49817, w_eco49818, w_eco49819, w_eco49820, w_eco49821, w_eco49822, w_eco49823, w_eco49824, w_eco49825, w_eco49826, w_eco49827, w_eco49828, w_eco49829, w_eco49830, w_eco49831, w_eco49832, w_eco49833, w_eco49834, w_eco49835, w_eco49836, w_eco49837, w_eco49838, w_eco49839, w_eco49840, w_eco49841, w_eco49842, w_eco49843, w_eco49844, w_eco49845, w_eco49846, w_eco49847, w_eco49848, w_eco49849, w_eco49850, w_eco49851, w_eco49852, w_eco49853, w_eco49854, w_eco49855, w_eco49856, w_eco49857, w_eco49858, w_eco49859, w_eco49860, w_eco49861, w_eco49862, w_eco49863, w_eco49864, w_eco49865, w_eco49866, w_eco49867, w_eco49868, w_eco49869, w_eco49870, w_eco49871, w_eco49872, w_eco49873, w_eco49874, w_eco49875, w_eco49876, w_eco49877, w_eco49878, w_eco49879, w_eco49880, w_eco49881, w_eco49882, w_eco49883, w_eco49884, w_eco49885, w_eco49886, w_eco49887, w_eco49888, w_eco49889, w_eco49890, w_eco49891, w_eco49892, w_eco49893, w_eco49894, w_eco49895, w_eco49896, w_eco49897, w_eco49898, w_eco49899, w_eco49900, w_eco49901, w_eco49902, w_eco49903, w_eco49904, w_eco49905, w_eco49906, w_eco49907, w_eco49908, w_eco49909, w_eco49910, w_eco49911, w_eco49912, w_eco49913, w_eco49914, w_eco49915, w_eco49916, w_eco49917, w_eco49918, w_eco49919, w_eco49920, w_eco49921, w_eco49922, w_eco49923, w_eco49924, w_eco49925, w_eco49926, w_eco49927, w_eco49928, w_eco49929, w_eco49930, w_eco49931, w_eco49932, w_eco49933, w_eco49934, w_eco49935, w_eco49936, w_eco49937, w_eco49938, w_eco49939, w_eco49940, w_eco49941, w_eco49942, w_eco49943, w_eco49944, w_eco49945, w_eco49946, w_eco49947, w_eco49948, w_eco49949, w_eco49950, w_eco49951, w_eco49952, w_eco49953, w_eco49954, w_eco49955, w_eco49956, w_eco49957, w_eco49958, w_eco49959, w_eco49960, w_eco49961, w_eco49962, w_eco49963, w_eco49964, w_eco49965, w_eco49966, w_eco49967, w_eco49968, w_eco49969, w_eco49970, w_eco49971, w_eco49972, w_eco49973, w_eco49974, w_eco49975, w_eco49976, w_eco49977, w_eco49978, w_eco49979, w_eco49980, w_eco49981, w_eco49982, w_eco49983, w_eco49984, w_eco49985, w_eco49986, w_eco49987, w_eco49988, w_eco49989, w_eco49990, w_eco49991, w_eco49992, w_eco49993, w_eco49994, w_eco49995, w_eco49996, w_eco49997, w_eco49998, w_eco49999, w_eco50000, w_eco50001, w_eco50002, w_eco50003, w_eco50004, w_eco50005, w_eco50006, w_eco50007, w_eco50008, w_eco50009, w_eco50010, w_eco50011, w_eco50012, w_eco50013, w_eco50014, w_eco50015, w_eco50016, w_eco50017, w_eco50018, w_eco50019, w_eco50020, w_eco50021, w_eco50022, w_eco50023, w_eco50024, w_eco50025, w_eco50026, w_eco50027, w_eco50028, w_eco50029, w_eco50030, w_eco50031, w_eco50032, w_eco50033, w_eco50034, w_eco50035, w_eco50036, w_eco50037, w_eco50038, w_eco50039, w_eco50040, w_eco50041, w_eco50042, w_eco50043, w_eco50044, w_eco50045, w_eco50046, w_eco50047, w_eco50048, w_eco50049, w_eco50050, w_eco50051, w_eco50052, w_eco50053, w_eco50054, w_eco50055, w_eco50056, w_eco50057, w_eco50058, w_eco50059, w_eco50060, w_eco50061, w_eco50062, w_eco50063, w_eco50064, w_eco50065, w_eco50066, w_eco50067, w_eco50068, w_eco50069, w_eco50070, w_eco50071, w_eco50072, w_eco50073, w_eco50074, w_eco50075, w_eco50076, w_eco50077, w_eco50078, w_eco50079, w_eco50080, w_eco50081, w_eco50082, w_eco50083, w_eco50084, w_eco50085, w_eco50086, w_eco50087, w_eco50088, w_eco50089, w_eco50090, w_eco50091, w_eco50092, w_eco50093, w_eco50094, w_eco50095, w_eco50096, w_eco50097, w_eco50098, w_eco50099, w_eco50100, w_eco50101, w_eco50102, w_eco50103, w_eco50104, w_eco50105, w_eco50106, w_eco50107, w_eco50108, w_eco50109, w_eco50110, w_eco50111, w_eco50112, w_eco50113, w_eco50114, w_eco50115, w_eco50116, w_eco50117, w_eco50118, w_eco50119, w_eco50120, w_eco50121, w_eco50122, w_eco50123, w_eco50124, w_eco50125, w_eco50126, w_eco50127, w_eco50128, w_eco50129, w_eco50130, w_eco50131, w_eco50132, w_eco50133, w_eco50134, w_eco50135, w_eco50136, w_eco50137, w_eco50138, w_eco50139, w_eco50140, w_eco50141, w_eco50142, w_eco50143, w_eco50144, w_eco50145, w_eco50146, w_eco50147, w_eco50148, w_eco50149, w_eco50150, w_eco50151, w_eco50152, w_eco50153, w_eco50154, w_eco50155, w_eco50156, w_eco50157, w_eco50158, w_eco50159, w_eco50160, w_eco50161, w_eco50162, w_eco50163, w_eco50164, w_eco50165, w_eco50166, w_eco50167, w_eco50168, w_eco50169, w_eco50170, w_eco50171, w_eco50172, w_eco50173, w_eco50174, w_eco50175, w_eco50176, w_eco50177, w_eco50178, w_eco50179, w_eco50180, w_eco50181, w_eco50182, w_eco50183, w_eco50184, w_eco50185, w_eco50186, w_eco50187, w_eco50188, w_eco50189, w_eco50190, w_eco50191, w_eco50192, w_eco50193, w_eco50194, w_eco50195, w_eco50196, w_eco50197, w_eco50198, w_eco50199, w_eco50200, w_eco50201, w_eco50202, w_eco50203, w_eco50204, w_eco50205, w_eco50206, w_eco50207, w_eco50208, w_eco50209, w_eco50210, w_eco50211, w_eco50212, w_eco50213, w_eco50214, w_eco50215, w_eco50216, w_eco50217, w_eco50218, w_eco50219, w_eco50220, w_eco50221, w_eco50222, w_eco50223, w_eco50224, w_eco50225, w_eco50226, w_eco50227, w_eco50228, w_eco50229, w_eco50230, w_eco50231, w_eco50232, w_eco50233, w_eco50234, w_eco50235, w_eco50236, w_eco50237, w_eco50238, w_eco50239, w_eco50240, w_eco50241, w_eco50242, w_eco50243, w_eco50244, w_eco50245, w_eco50246, w_eco50247, w_eco50248, w_eco50249, w_eco50250, w_eco50251, w_eco50252, w_eco50253, w_eco50254, w_eco50255, w_eco50256, w_eco50257, w_eco50258, w_eco50259, w_eco50260, w_eco50261, w_eco50262, w_eco50263, w_eco50264, w_eco50265, w_eco50266, w_eco50267, w_eco50268, w_eco50269, w_eco50270, w_eco50271, w_eco50272, w_eco50273, w_eco50274, w_eco50275, w_eco50276, w_eco50277, w_eco50278, w_eco50279, w_eco50280, w_eco50281, w_eco50282, w_eco50283, w_eco50284, w_eco50285, w_eco50286, w_eco50287, w_eco50288, w_eco50289, w_eco50290, w_eco50291, w_eco50292, w_eco50293, w_eco50294, w_eco50295, w_eco50296, w_eco50297, w_eco50298, w_eco50299, w_eco50300, w_eco50301, w_eco50302, w_eco50303, w_eco50304, w_eco50305, w_eco50306, w_eco50307, w_eco50308, w_eco50309, w_eco50310, w_eco50311, w_eco50312, w_eco50313, w_eco50314, w_eco50315, w_eco50316, w_eco50317, w_eco50318, w_eco50319, w_eco50320, w_eco50321, w_eco50322, w_eco50323, w_eco50324, w_eco50325, w_eco50326, w_eco50327, w_eco50328, w_eco50329, w_eco50330, w_eco50331, w_eco50332, w_eco50333, w_eco50334, w_eco50335, w_eco50336, w_eco50337, w_eco50338, w_eco50339, w_eco50340, w_eco50341, w_eco50342, w_eco50343, w_eco50344, w_eco50345, w_eco50346, w_eco50347, w_eco50348, w_eco50349, w_eco50350, w_eco50351, w_eco50352, w_eco50353, w_eco50354, w_eco50355, w_eco50356, w_eco50357, w_eco50358, w_eco50359, w_eco50360, w_eco50361, w_eco50362, w_eco50363, w_eco50364, w_eco50365, w_eco50366, w_eco50367, w_eco50368, w_eco50369, w_eco50370, w_eco50371, w_eco50372, w_eco50373, w_eco50374, w_eco50375, w_eco50376, w_eco50377, w_eco50378, w_eco50379, w_eco50380, w_eco50381, w_eco50382, w_eco50383, w_eco50384, w_eco50385, w_eco50386, w_eco50387, w_eco50388, w_eco50389, w_eco50390, w_eco50391, w_eco50392, w_eco50393, w_eco50394, w_eco50395, w_eco50396, w_eco50397, w_eco50398, w_eco50399, w_eco50400, w_eco50401, w_eco50402, w_eco50403, w_eco50404, w_eco50405, w_eco50406, w_eco50407, w_eco50408, w_eco50409, w_eco50410, w_eco50411, w_eco50412, w_eco50413, w_eco50414, w_eco50415, w_eco50416, w_eco50417, w_eco50418, w_eco50419, w_eco50420, w_eco50421, w_eco50422, w_eco50423, w_eco50424, w_eco50425, w_eco50426, w_eco50427, w_eco50428, w_eco50429, w_eco50430, w_eco50431, w_eco50432, w_eco50433, w_eco50434, w_eco50435, w_eco50436, w_eco50437, w_eco50438, w_eco50439, w_eco50440, w_eco50441, w_eco50442, w_eco50443, w_eco50444, w_eco50445, w_eco50446, w_eco50447, w_eco50448, w_eco50449, w_eco50450, w_eco50451, w_eco50452, w_eco50453, w_eco50454, w_eco50455, w_eco50456, w_eco50457, w_eco50458, w_eco50459, w_eco50460, w_eco50461, w_eco50462, w_eco50463, w_eco50464, w_eco50465, w_eco50466, w_eco50467, w_eco50468, w_eco50469, w_eco50470, w_eco50471, w_eco50472, w_eco50473, w_eco50474, w_eco50475, w_eco50476, w_eco50477, w_eco50478, w_eco50479, w_eco50480, w_eco50481, w_eco50482, w_eco50483, w_eco50484, w_eco50485, w_eco50486, w_eco50487, w_eco50488, w_eco50489, w_eco50490, w_eco50491, w_eco50492, w_eco50493, w_eco50494, w_eco50495, w_eco50496, w_eco50497, w_eco50498, w_eco50499, w_eco50500, w_eco50501, w_eco50502, w_eco50503, w_eco50504, w_eco50505, w_eco50506, w_eco50507, w_eco50508, w_eco50509, w_eco50510, w_eco50511, w_eco50512, w_eco50513, w_eco50514, w_eco50515, w_eco50516, w_eco50517, w_eco50518, w_eco50519, w_eco50520, w_eco50521, w_eco50522, w_eco50523, w_eco50524, w_eco50525, w_eco50526, w_eco50527, w_eco50528, w_eco50529, w_eco50530, w_eco50531, w_eco50532, w_eco50533, w_eco50534, w_eco50535, w_eco50536, w_eco50537, w_eco50538, w_eco50539, w_eco50540, w_eco50541, w_eco50542, w_eco50543, w_eco50544, w_eco50545, w_eco50546, w_eco50547, w_eco50548, w_eco50549, w_eco50550, w_eco50551, w_eco50552, w_eco50553, w_eco50554, w_eco50555, w_eco50556, w_eco50557, w_eco50558, w_eco50559, w_eco50560, w_eco50561, w_eco50562, w_eco50563, w_eco50564, w_eco50565, w_eco50566, w_eco50567, w_eco50568, w_eco50569, w_eco50570, w_eco50571, w_eco50572, w_eco50573, w_eco50574, w_eco50575, w_eco50576, w_eco50577, w_eco50578, w_eco50579, w_eco50580, w_eco50581, w_eco50582, w_eco50583, w_eco50584, w_eco50585, w_eco50586, w_eco50587, w_eco50588, w_eco50589, w_eco50590, w_eco50591, w_eco50592, w_eco50593, w_eco50594, w_eco50595, w_eco50596, w_eco50597, w_eco50598, w_eco50599, w_eco50600, w_eco50601, w_eco50602, w_eco50603, w_eco50604, w_eco50605, w_eco50606, w_eco50607, w_eco50608, w_eco50609, w_eco50610, w_eco50611, w_eco50612, w_eco50613, w_eco50614, w_eco50615, w_eco50616, w_eco50617, w_eco50618, w_eco50619, w_eco50620, w_eco50621, w_eco50622, w_eco50623, w_eco50624, w_eco50625, w_eco50626, w_eco50627, w_eco50628, w_eco50629, w_eco50630, w_eco50631, w_eco50632, w_eco50633, w_eco50634, w_eco50635, w_eco50636, w_eco50637, w_eco50638, w_eco50639, w_eco50640, w_eco50641, w_eco50642, w_eco50643, w_eco50644, w_eco50645, w_eco50646, w_eco50647, w_eco50648, w_eco50649, w_eco50650, w_eco50651, w_eco50652, w_eco50653, w_eco50654, w_eco50655, w_eco50656, w_eco50657, w_eco50658, w_eco50659, w_eco50660, w_eco50661, w_eco50662, w_eco50663, w_eco50664, w_eco50665, w_eco50666, w_eco50667, w_eco50668, w_eco50669, w_eco50670, w_eco50671, w_eco50672, w_eco50673, w_eco50674, w_eco50675, w_eco50676, w_eco50677, w_eco50678, w_eco50679, w_eco50680, w_eco50681, w_eco50682, w_eco50683, w_eco50684, w_eco50685, w_eco50686, w_eco50687, w_eco50688, w_eco50689, w_eco50690, w_eco50691, w_eco50692, w_eco50693, w_eco50694, w_eco50695, w_eco50696, w_eco50697, w_eco50698, w_eco50699, w_eco50700, w_eco50701, w_eco50702, w_eco50703, w_eco50704, w_eco50705, w_eco50706, w_eco50707, w_eco50708, w_eco50709, w_eco50710, w_eco50711, w_eco50712, w_eco50713, w_eco50714, w_eco50715, w_eco50716, w_eco50717, w_eco50718, w_eco50719, w_eco50720, w_eco50721, w_eco50722, w_eco50723, w_eco50724, w_eco50725, w_eco50726, w_eco50727, w_eco50728, w_eco50729, w_eco50730, w_eco50731, w_eco50732, w_eco50733, w_eco50734, w_eco50735, w_eco50736, w_eco50737, w_eco50738, w_eco50739, w_eco50740, w_eco50741, w_eco50742, w_eco50743, w_eco50744, w_eco50745, w_eco50746, w_eco50747, w_eco50748, w_eco50749, w_eco50750, w_eco50751, w_eco50752, w_eco50753, w_eco50754, w_eco50755, w_eco50756, w_eco50757, w_eco50758, w_eco50759, w_eco50760, w_eco50761, w_eco50762, w_eco50763, w_eco50764, w_eco50765, w_eco50766, w_eco50767, w_eco50768, w_eco50769, w_eco50770, w_eco50771, w_eco50772, w_eco50773, w_eco50774, w_eco50775, w_eco50776, w_eco50777, w_eco50778, w_eco50779, w_eco50780, w_eco50781, w_eco50782, w_eco50783, w_eco50784, w_eco50785, w_eco50786, w_eco50787, w_eco50788, w_eco50789, w_eco50790, w_eco50791, w_eco50792, w_eco50793, w_eco50794, w_eco50795, w_eco50796, w_eco50797, w_eco50798, w_eco50799, w_eco50800, w_eco50801, w_eco50802, w_eco50803, w_eco50804, w_eco50805, w_eco50806, w_eco50807, w_eco50808, w_eco50809, w_eco50810, w_eco50811, w_eco50812, w_eco50813, w_eco50814, w_eco50815, w_eco50816, w_eco50817, w_eco50818, w_eco50819, w_eco50820, w_eco50821, w_eco50822, w_eco50823, w_eco50824, w_eco50825, w_eco50826, w_eco50827, w_eco50828, w_eco50829, w_eco50830, w_eco50831, w_eco50832, w_eco50833, w_eco50834, w_eco50835, w_eco50836, w_eco50837, w_eco50838, w_eco50839, w_eco50840, w_eco50841, w_eco50842, w_eco50843, w_eco50844, w_eco50845, w_eco50846, w_eco50847, w_eco50848, w_eco50849, w_eco50850, w_eco50851, w_eco50852, w_eco50853, w_eco50854, w_eco50855, w_eco50856, w_eco50857, w_eco50858, w_eco50859, w_eco50860, w_eco50861, w_eco50862, w_eco50863, w_eco50864, w_eco50865, w_eco50866, w_eco50867, w_eco50868, w_eco50869, w_eco50870, w_eco50871, w_eco50872, w_eco50873, w_eco50874, w_eco50875, w_eco50876, w_eco50877, w_eco50878, w_eco50879, w_eco50880, w_eco50881, w_eco50882, w_eco50883, w_eco50884, w_eco50885, w_eco50886, w_eco50887, w_eco50888, w_eco50889, w_eco50890, w_eco50891, w_eco50892, w_eco50893, w_eco50894, w_eco50895, w_eco50896, w_eco50897, w_eco50898, w_eco50899, w_eco50900, w_eco50901, w_eco50902, w_eco50903, w_eco50904, w_eco50905, w_eco50906, w_eco50907, w_eco50908, w_eco50909, w_eco50910, w_eco50911, w_eco50912, w_eco50913, w_eco50914, w_eco50915, w_eco50916, w_eco50917, w_eco50918, w_eco50919, w_eco50920, w_eco50921, w_eco50922, w_eco50923, w_eco50924, w_eco50925, w_eco50926, w_eco50927, w_eco50928, w_eco50929, w_eco50930, w_eco50931, w_eco50932, w_eco50933, w_eco50934, w_eco50935, w_eco50936, w_eco50937, w_eco50938, w_eco50939, w_eco50940, w_eco50941, w_eco50942, w_eco50943, w_eco50944, w_eco50945, w_eco50946, w_eco50947, w_eco50948, w_eco50949, w_eco50950, w_eco50951, w_eco50952, w_eco50953, w_eco50954, w_eco50955, w_eco50956, w_eco50957, w_eco50958, w_eco50959, w_eco50960, w_eco50961, w_eco50962, w_eco50963, w_eco50964, w_eco50965, w_eco50966, w_eco50967, w_eco50968, w_eco50969, w_eco50970, w_eco50971, w_eco50972, w_eco50973, w_eco50974, w_eco50975, w_eco50976, w_eco50977, w_eco50978, w_eco50979, w_eco50980, w_eco50981, w_eco50982, w_eco50983, w_eco50984, w_eco50985, w_eco50986, w_eco50987, w_eco50988, w_eco50989, w_eco50990, w_eco50991, w_eco50992, w_eco50993, w_eco50994, w_eco50995, w_eco50996, w_eco50997, w_eco50998, w_eco50999, w_eco51000, w_eco51001, w_eco51002, w_eco51003, w_eco51004, w_eco51005, w_eco51006, w_eco51007, w_eco51008, w_eco51009, w_eco51010, w_eco51011, w_eco51012, w_eco51013, w_eco51014, w_eco51015, w_eco51016, w_eco51017, w_eco51018, w_eco51019, w_eco51020, w_eco51021, w_eco51022, w_eco51023, w_eco51024, w_eco51025, w_eco51026, w_eco51027, w_eco51028, w_eco51029, w_eco51030, w_eco51031, w_eco51032, w_eco51033, w_eco51034, w_eco51035, w_eco51036, w_eco51037, w_eco51038, w_eco51039, w_eco51040, w_eco51041, w_eco51042, w_eco51043, w_eco51044, w_eco51045, w_eco51046, w_eco51047, w_eco51048, w_eco51049, w_eco51050, w_eco51051, w_eco51052, w_eco51053, w_eco51054, w_eco51055, w_eco51056, w_eco51057, w_eco51058, w_eco51059, w_eco51060, w_eco51061, w_eco51062, w_eco51063, w_eco51064, w_eco51065, w_eco51066, w_eco51067, w_eco51068, w_eco51069, w_eco51070, w_eco51071, w_eco51072, w_eco51073, w_eco51074, w_eco51075, w_eco51076, w_eco51077, w_eco51078, w_eco51079, w_eco51080, w_eco51081, w_eco51082, w_eco51083, w_eco51084, w_eco51085, w_eco51086, w_eco51087, w_eco51088, w_eco51089, w_eco51090, w_eco51091, w_eco51092, w_eco51093, w_eco51094, w_eco51095, w_eco51096, w_eco51097, w_eco51098, w_eco51099, w_eco51100, w_eco51101, w_eco51102, w_eco51103, w_eco51104, w_eco51105, w_eco51106, w_eco51107, w_eco51108, w_eco51109, w_eco51110, w_eco51111, w_eco51112, w_eco51113, w_eco51114, w_eco51115, w_eco51116, w_eco51117, w_eco51118, w_eco51119, w_eco51120, w_eco51121, w_eco51122, w_eco51123, w_eco51124, w_eco51125, w_eco51126, w_eco51127, w_eco51128, w_eco51129, w_eco51130, w_eco51131, w_eco51132, w_eco51133, w_eco51134, w_eco51135, w_eco51136, w_eco51137, w_eco51138, w_eco51139, w_eco51140, w_eco51141, w_eco51142, w_eco51143, w_eco51144, w_eco51145, w_eco51146, w_eco51147, w_eco51148, w_eco51149, w_eco51150, w_eco51151, w_eco51152, w_eco51153, w_eco51154, w_eco51155, w_eco51156, w_eco51157, w_eco51158, w_eco51159, w_eco51160, w_eco51161, w_eco51162, w_eco51163, w_eco51164, w_eco51165, w_eco51166, w_eco51167, w_eco51168, w_eco51169, w_eco51170, w_eco51171, w_eco51172, w_eco51173, w_eco51174, w_eco51175, w_eco51176, w_eco51177, w_eco51178, w_eco51179, w_eco51180, w_eco51181, w_eco51182, w_eco51183, w_eco51184, w_eco51185, w_eco51186, w_eco51187, w_eco51188, w_eco51189, w_eco51190, w_eco51191, w_eco51192, w_eco51193, w_eco51194, w_eco51195, w_eco51196, w_eco51197, w_eco51198, w_eco51199, w_eco51200, w_eco51201, w_eco51202, w_eco51203, w_eco51204, w_eco51205, w_eco51206, w_eco51207, w_eco51208, w_eco51209, w_eco51210, w_eco51211, w_eco51212, w_eco51213, w_eco51214, w_eco51215, w_eco51216, w_eco51217, w_eco51218, w_eco51219, w_eco51220, w_eco51221, w_eco51222, w_eco51223, w_eco51224, w_eco51225, w_eco51226, w_eco51227, w_eco51228, w_eco51229, w_eco51230, w_eco51231, w_eco51232, w_eco51233, w_eco51234, w_eco51235, w_eco51236, w_eco51237, w_eco51238, w_eco51239, w_eco51240, w_eco51241, w_eco51242, w_eco51243, w_eco51244, w_eco51245, w_eco51246, w_eco51247, w_eco51248, w_eco51249, w_eco51250, w_eco51251, w_eco51252, w_eco51253, w_eco51254, w_eco51255, w_eco51256, w_eco51257, w_eco51258, w_eco51259, w_eco51260, w_eco51261, w_eco51262, w_eco51263, w_eco51264, w_eco51265, w_eco51266, w_eco51267, w_eco51268, w_eco51269, w_eco51270, w_eco51271, w_eco51272, w_eco51273, w_eco51274, w_eco51275, w_eco51276, w_eco51277, w_eco51278, w_eco51279, w_eco51280, w_eco51281, w_eco51282, w_eco51283, w_eco51284, w_eco51285, w_eco51286, w_eco51287, w_eco51288, w_eco51289, w_eco51290, w_eco51291, w_eco51292, w_eco51293, w_eco51294, w_eco51295, w_eco51296, w_eco51297, w_eco51298, w_eco51299, w_eco51300, w_eco51301, w_eco51302, w_eco51303, w_eco51304, w_eco51305, w_eco51306, w_eco51307, w_eco51308, w_eco51309, w_eco51310, w_eco51311, w_eco51312, w_eco51313, w_eco51314, w_eco51315, w_eco51316, w_eco51317, w_eco51318, w_eco51319, w_eco51320, w_eco51321, w_eco51322, w_eco51323, w_eco51324, w_eco51325, w_eco51326, w_eco51327, w_eco51328, w_eco51329, w_eco51330, w_eco51331, w_eco51332, w_eco51333, w_eco51334, w_eco51335, w_eco51336, w_eco51337, w_eco51338, w_eco51339, w_eco51340, w_eco51341, w_eco51342, w_eco51343, w_eco51344, w_eco51345, w_eco51346, w_eco51347, w_eco51348, w_eco51349, w_eco51350, w_eco51351, w_eco51352, w_eco51353, w_eco51354, w_eco51355, w_eco51356, w_eco51357, w_eco51358, w_eco51359, w_eco51360, w_eco51361, w_eco51362, w_eco51363, w_eco51364, w_eco51365, w_eco51366, w_eco51367, w_eco51368, w_eco51369, w_eco51370, w_eco51371, w_eco51372, w_eco51373, w_eco51374, w_eco51375, w_eco51376, w_eco51377, w_eco51378, w_eco51379, w_eco51380, w_eco51381, w_eco51382, w_eco51383, w_eco51384, w_eco51385, w_eco51386, w_eco51387, w_eco51388, w_eco51389, w_eco51390, w_eco51391, w_eco51392, w_eco51393, w_eco51394, w_eco51395, w_eco51396, w_eco51397, w_eco51398, w_eco51399, w_eco51400, w_eco51401, w_eco51402, w_eco51403, w_eco51404, w_eco51405, w_eco51406, w_eco51407, w_eco51408, w_eco51409, w_eco51410, w_eco51411, w_eco51412, w_eco51413, w_eco51414, w_eco51415, w_eco51416, w_eco51417, w_eco51418, w_eco51419, w_eco51420, w_eco51421, w_eco51422, w_eco51423, w_eco51424, w_eco51425, w_eco51426, w_eco51427, w_eco51428, w_eco51429, w_eco51430, w_eco51431, w_eco51432, w_eco51433, w_eco51434, w_eco51435, w_eco51436, w_eco51437, w_eco51438, w_eco51439, w_eco51440, w_eco51441, w_eco51442, w_eco51443, w_eco51444, w_eco51445, w_eco51446, w_eco51447, w_eco51448, w_eco51449, w_eco51450, w_eco51451, w_eco51452, w_eco51453, w_eco51454, w_eco51455, w_eco51456, w_eco51457, w_eco51458, w_eco51459, w_eco51460, w_eco51461, w_eco51462, w_eco51463, w_eco51464, w_eco51465, w_eco51466, w_eco51467, w_eco51468, w_eco51469, w_eco51470, w_eco51471, w_eco51472, w_eco51473, w_eco51474, w_eco51475, w_eco51476, w_eco51477, w_eco51478, w_eco51479, w_eco51480, w_eco51481, w_eco51482, w_eco51483, w_eco51484, w_eco51485, w_eco51486, w_eco51487, w_eco51488, w_eco51489, w_eco51490, w_eco51491, w_eco51492, w_eco51493, w_eco51494, w_eco51495, w_eco51496, w_eco51497, w_eco51498, w_eco51499, w_eco51500, w_eco51501, w_eco51502, w_eco51503, w_eco51504, w_eco51505, w_eco51506, w_eco51507, w_eco51508, w_eco51509, w_eco51510, w_eco51511, w_eco51512, w_eco51513, w_eco51514, w_eco51515, w_eco51516, w_eco51517, w_eco51518, w_eco51519, w_eco51520, w_eco51521, w_eco51522, w_eco51523, w_eco51524, w_eco51525, w_eco51526, w_eco51527, w_eco51528, w_eco51529, w_eco51530, w_eco51531, w_eco51532, w_eco51533, w_eco51534, w_eco51535, w_eco51536, w_eco51537, w_eco51538, w_eco51539, w_eco51540, w_eco51541, w_eco51542, w_eco51543, w_eco51544, w_eco51545, w_eco51546, w_eco51547, w_eco51548, w_eco51549, w_eco51550, w_eco51551, w_eco51552, w_eco51553, w_eco51554, w_eco51555, w_eco51556, w_eco51557, w_eco51558, w_eco51559, w_eco51560, w_eco51561, w_eco51562, w_eco51563, w_eco51564, w_eco51565, w_eco51566, w_eco51567, w_eco51568, w_eco51569, w_eco51570, w_eco51571, w_eco51572, w_eco51573, w_eco51574, w_eco51575, w_eco51576, w_eco51577, w_eco51578, w_eco51579, w_eco51580, w_eco51581, w_eco51582, w_eco51583, w_eco51584, w_eco51585, w_eco51586, w_eco51587, w_eco51588, w_eco51589, w_eco51590, w_eco51591, w_eco51592, w_eco51593, w_eco51594, w_eco51595, w_eco51596, w_eco51597, w_eco51598, w_eco51599, w_eco51600, w_eco51601, w_eco51602, w_eco51603, w_eco51604, w_eco51605, w_eco51606, w_eco51607, w_eco51608, w_eco51609, w_eco51610, w_eco51611, w_eco51612, w_eco51613, w_eco51614, w_eco51615, w_eco51616, w_eco51617, w_eco51618, w_eco51619, w_eco51620, w_eco51621, w_eco51622, w_eco51623, w_eco51624, w_eco51625, w_eco51626, w_eco51627, w_eco51628, w_eco51629, w_eco51630, w_eco51631, w_eco51632, w_eco51633, w_eco51634, w_eco51635, w_eco51636, w_eco51637, w_eco51638, w_eco51639, w_eco51640, w_eco51641, w_eco51642, w_eco51643, w_eco51644, w_eco51645, w_eco51646, w_eco51647, w_eco51648, w_eco51649, w_eco51650, w_eco51651, w_eco51652, w_eco51653, w_eco51654, w_eco51655, w_eco51656, w_eco51657, w_eco51658, w_eco51659, w_eco51660, w_eco51661, w_eco51662, w_eco51663, w_eco51664, w_eco51665, w_eco51666, w_eco51667, w_eco51668, w_eco51669, w_eco51670, w_eco51671, w_eco51672, w_eco51673, w_eco51674, w_eco51675, w_eco51676, w_eco51677, w_eco51678, w_eco51679, w_eco51680, w_eco51681, w_eco51682, w_eco51683, w_eco51684, w_eco51685, w_eco51686, w_eco51687, w_eco51688, w_eco51689, w_eco51690, w_eco51691, w_eco51692, w_eco51693, w_eco51694, w_eco51695, w_eco51696, w_eco51697, w_eco51698, w_eco51699, w_eco51700, w_eco51701, w_eco51702, w_eco51703, w_eco51704, w_eco51705, w_eco51706, w_eco51707, w_eco51708, w_eco51709, w_eco51710, w_eco51711, w_eco51712, w_eco51713, w_eco51714, w_eco51715, w_eco51716, w_eco51717, w_eco51718, w_eco51719, w_eco51720, w_eco51721, w_eco51722, w_eco51723, w_eco51724, w_eco51725, w_eco51726, w_eco51727, w_eco51728, w_eco51729, w_eco51730, w_eco51731, w_eco51732, w_eco51733, w_eco51734, w_eco51735, w_eco51736, w_eco51737, w_eco51738, w_eco51739, w_eco51740, w_eco51741, w_eco51742, w_eco51743, w_eco51744, w_eco51745, w_eco51746, w_eco51747, w_eco51748, w_eco51749, w_eco51750, w_eco51751, w_eco51752, w_eco51753, w_eco51754, w_eco51755, w_eco51756, w_eco51757, w_eco51758, w_eco51759, w_eco51760, w_eco51761, w_eco51762, w_eco51763, w_eco51764, w_eco51765, w_eco51766, w_eco51767, w_eco51768, w_eco51769, w_eco51770, w_eco51771, w_eco51772, w_eco51773, w_eco51774, w_eco51775, w_eco51776, w_eco51777, w_eco51778, w_eco51779, w_eco51780, w_eco51781, w_eco51782, w_eco51783, w_eco51784, w_eco51785, w_eco51786, w_eco51787, w_eco51788, w_eco51789, w_eco51790, w_eco51791, w_eco51792, w_eco51793, w_eco51794, w_eco51795, w_eco51796, w_eco51797, w_eco51798, w_eco51799, w_eco51800, w_eco51801, w_eco51802, w_eco51803, w_eco51804, w_eco51805, w_eco51806, w_eco51807, w_eco51808, w_eco51809, w_eco51810, w_eco51811, w_eco51812, w_eco51813, w_eco51814, w_eco51815, w_eco51816, w_eco51817, w_eco51818, w_eco51819, w_eco51820, w_eco51821, w_eco51822, w_eco51823, w_eco51824, w_eco51825, w_eco51826, w_eco51827, w_eco51828, w_eco51829, w_eco51830, w_eco51831, w_eco51832, w_eco51833, w_eco51834, w_eco51835, w_eco51836, w_eco51837, w_eco51838, w_eco51839, w_eco51840, w_eco51841, w_eco51842, w_eco51843, w_eco51844, w_eco51845, w_eco51846, w_eco51847, w_eco51848, w_eco51849, w_eco51850, w_eco51851, w_eco51852, w_eco51853, w_eco51854, w_eco51855, w_eco51856, w_eco51857, w_eco51858, w_eco51859, w_eco51860, w_eco51861, w_eco51862, w_eco51863, w_eco51864, w_eco51865, w_eco51866, w_eco51867, w_eco51868, w_eco51869, w_eco51870, w_eco51871, w_eco51872, w_eco51873, w_eco51874, w_eco51875, w_eco51876, w_eco51877, w_eco51878, w_eco51879, w_eco51880, w_eco51881, w_eco51882, w_eco51883, w_eco51884, w_eco51885, w_eco51886, w_eco51887, w_eco51888, w_eco51889, w_eco51890, w_eco51891, w_eco51892, w_eco51893, w_eco51894, w_eco51895, w_eco51896, w_eco51897, w_eco51898, w_eco51899, w_eco51900, w_eco51901, w_eco51902, w_eco51903, w_eco51904, w_eco51905, w_eco51906, w_eco51907, w_eco51908, w_eco51909, w_eco51910, w_eco51911, w_eco51912, w_eco51913, w_eco51914, w_eco51915, w_eco51916, w_eco51917, w_eco51918, w_eco51919, w_eco51920, w_eco51921, w_eco51922, w_eco51923, w_eco51924, w_eco51925, w_eco51926, w_eco51927, w_eco51928, w_eco51929, w_eco51930, w_eco51931, w_eco51932, w_eco51933, w_eco51934, w_eco51935, w_eco51936, w_eco51937, w_eco51938, w_eco51939, w_eco51940, w_eco51941, w_eco51942, w_eco51943, w_eco51944, w_eco51945, w_eco51946, w_eco51947, w_eco51948, w_eco51949, w_eco51950, w_eco51951, w_eco51952, w_eco51953, w_eco51954, w_eco51955, w_eco51956, w_eco51957, w_eco51958, w_eco51959, w_eco51960, w_eco51961, w_eco51962, w_eco51963, w_eco51964, w_eco51965, w_eco51966, w_eco51967, w_eco51968, w_eco51969, w_eco51970, w_eco51971, w_eco51972, w_eco51973, w_eco51974, w_eco51975, w_eco51976, w_eco51977, w_eco51978, w_eco51979, w_eco51980, w_eco51981, w_eco51982, w_eco51983, w_eco51984, w_eco51985, w_eco51986, w_eco51987, w_eco51988, w_eco51989, w_eco51990, w_eco51991, w_eco51992, w_eco51993, w_eco51994, w_eco51995, w_eco51996, w_eco51997, w_eco51998, w_eco51999, w_eco52000, w_eco52001, w_eco52002, w_eco52003, w_eco52004, w_eco52005, w_eco52006, w_eco52007, w_eco52008, w_eco52009, w_eco52010, w_eco52011, w_eco52012, w_eco52013, w_eco52014, w_eco52015, w_eco52016, w_eco52017, w_eco52018, w_eco52019, w_eco52020, w_eco52021, w_eco52022, w_eco52023, w_eco52024, w_eco52025, w_eco52026, w_eco52027, w_eco52028, w_eco52029, w_eco52030, w_eco52031, w_eco52032, w_eco52033, w_eco52034, w_eco52035, w_eco52036, w_eco52037, w_eco52038, w_eco52039, w_eco52040, w_eco52041, w_eco52042, w_eco52043, w_eco52044, w_eco52045, w_eco52046, w_eco52047, w_eco52048, w_eco52049, w_eco52050, w_eco52051, w_eco52052, w_eco52053, w_eco52054, w_eco52055, w_eco52056, w_eco52057, w_eco52058, w_eco52059, w_eco52060, w_eco52061, w_eco52062, w_eco52063, w_eco52064, w_eco52065, w_eco52066, w_eco52067, w_eco52068, w_eco52069, w_eco52070, w_eco52071, w_eco52072, w_eco52073, w_eco52074, w_eco52075, w_eco52076, w_eco52077, w_eco52078, w_eco52079, w_eco52080, w_eco52081, w_eco52082, w_eco52083, w_eco52084, w_eco52085, w_eco52086, w_eco52087, w_eco52088, w_eco52089, w_eco52090, w_eco52091, w_eco52092, w_eco52093, w_eco52094, w_eco52095, w_eco52096, w_eco52097, w_eco52098, w_eco52099, w_eco52100, w_eco52101, w_eco52102, w_eco52103, w_eco52104, w_eco52105, w_eco52106, w_eco52107, w_eco52108, w_eco52109, w_eco52110, w_eco52111, w_eco52112, w_eco52113, w_eco52114, w_eco52115, w_eco52116, w_eco52117, w_eco52118, w_eco52119, w_eco52120, w_eco52121, w_eco52122, w_eco52123, w_eco52124, w_eco52125, w_eco52126, w_eco52127, w_eco52128, w_eco52129, w_eco52130, w_eco52131, w_eco52132, w_eco52133, w_eco52134, w_eco52135, w_eco52136, w_eco52137, w_eco52138, w_eco52139, w_eco52140, w_eco52141, w_eco52142, w_eco52143, w_eco52144, w_eco52145, w_eco52146, w_eco52147, w_eco52148, w_eco52149, w_eco52150, w_eco52151, w_eco52152, w_eco52153, w_eco52154, w_eco52155, w_eco52156, w_eco52157, w_eco52158, w_eco52159, w_eco52160, w_eco52161, w_eco52162, w_eco52163, w_eco52164, w_eco52165, w_eco52166, w_eco52167, w_eco52168, w_eco52169, w_eco52170, w_eco52171, w_eco52172, w_eco52173, w_eco52174, w_eco52175, w_eco52176, w_eco52177, w_eco52178, w_eco52179, w_eco52180, w_eco52181, w_eco52182, w_eco52183, w_eco52184, w_eco52185, w_eco52186, w_eco52187, w_eco52188, w_eco52189, w_eco52190, w_eco52191, w_eco52192, w_eco52193, w_eco52194, w_eco52195, w_eco52196, w_eco52197, w_eco52198, w_eco52199, w_eco52200, w_eco52201, w_eco52202, w_eco52203, w_eco52204, w_eco52205, w_eco52206, w_eco52207, w_eco52208, w_eco52209, w_eco52210, w_eco52211, w_eco52212, w_eco52213, w_eco52214, w_eco52215, w_eco52216, w_eco52217, w_eco52218, w_eco52219, w_eco52220, w_eco52221, w_eco52222, w_eco52223, w_eco52224, w_eco52225, w_eco52226, w_eco52227, w_eco52228, w_eco52229, w_eco52230, w_eco52231, w_eco52232, w_eco52233, w_eco52234, w_eco52235, w_eco52236, w_eco52237, w_eco52238, w_eco52239, w_eco52240, w_eco52241, w_eco52242, w_eco52243, w_eco52244, w_eco52245, w_eco52246, w_eco52247, w_eco52248, w_eco52249, w_eco52250, w_eco52251, w_eco52252, w_eco52253, w_eco52254, w_eco52255, w_eco52256, w_eco52257, w_eco52258, w_eco52259, w_eco52260, w_eco52261, w_eco52262, w_eco52263, w_eco52264, w_eco52265, w_eco52266, w_eco52267, w_eco52268, w_eco52269, w_eco52270, w_eco52271, w_eco52272, w_eco52273, w_eco52274, w_eco52275, w_eco52276, w_eco52277, w_eco52278, w_eco52279, w_eco52280, w_eco52281, w_eco52282, w_eco52283, w_eco52284, w_eco52285, w_eco52286, w_eco52287, w_eco52288, w_eco52289, w_eco52290, w_eco52291, w_eco52292, w_eco52293, w_eco52294, w_eco52295, w_eco52296, w_eco52297, w_eco52298, w_eco52299, w_eco52300, w_eco52301, w_eco52302, w_eco52303, w_eco52304, w_eco52305, w_eco52306, w_eco52307, w_eco52308, w_eco52309, w_eco52310, w_eco52311, w_eco52312, w_eco52313, w_eco52314, w_eco52315, w_eco52316, w_eco52317, w_eco52318, w_eco52319, w_eco52320, w_eco52321, w_eco52322, w_eco52323, w_eco52324, w_eco52325, w_eco52326, w_eco52327, w_eco52328, w_eco52329, w_eco52330, w_eco52331, w_eco52332, w_eco52333, w_eco52334, w_eco52335, w_eco52336, w_eco52337, w_eco52338, w_eco52339, w_eco52340, w_eco52341, w_eco52342, w_eco52343, w_eco52344, w_eco52345, w_eco52346, w_eco52347, w_eco52348, w_eco52349, w_eco52350, w_eco52351, w_eco52352, w_eco52353, w_eco52354, w_eco52355, w_eco52356, w_eco52357, w_eco52358, w_eco52359, w_eco52360, w_eco52361, w_eco52362, w_eco52363, w_eco52364, w_eco52365, w_eco52366, w_eco52367, w_eco52368, w_eco52369, w_eco52370, w_eco52371, w_eco52372, w_eco52373, w_eco52374, w_eco52375, w_eco52376, w_eco52377, w_eco52378, w_eco52379, w_eco52380, w_eco52381, w_eco52382, w_eco52383, w_eco52384, w_eco52385, w_eco52386, w_eco52387, w_eco52388, w_eco52389, w_eco52390, w_eco52391, w_eco52392, w_eco52393, w_eco52394, w_eco52395, w_eco52396, w_eco52397, w_eco52398, w_eco52399, w_eco52400, w_eco52401, w_eco52402, w_eco52403, w_eco52404, w_eco52405, w_eco52406, w_eco52407, w_eco52408, w_eco52409, w_eco52410, w_eco52411, w_eco52412, w_eco52413, w_eco52414, w_eco52415, w_eco52416, w_eco52417, w_eco52418, w_eco52419, w_eco52420, w_eco52421, w_eco52422, w_eco52423, w_eco52424, w_eco52425, w_eco52426, w_eco52427, w_eco52428, w_eco52429, w_eco52430, w_eco52431, w_eco52432, w_eco52433, w_eco52434, w_eco52435, w_eco52436, w_eco52437, w_eco52438, w_eco52439, w_eco52440, w_eco52441, w_eco52442, w_eco52443, w_eco52444, w_eco52445, w_eco52446, w_eco52447, w_eco52448, w_eco52449, w_eco52450, w_eco52451, w_eco52452, w_eco52453, w_eco52454, w_eco52455, w_eco52456, w_eco52457, w_eco52458, w_eco52459, w_eco52460, w_eco52461, w_eco52462, w_eco52463, w_eco52464, w_eco52465, w_eco52466, w_eco52467, w_eco52468, w_eco52469, w_eco52470, w_eco52471, w_eco52472, w_eco52473, w_eco52474, w_eco52475, w_eco52476, w_eco52477, w_eco52478, w_eco52479, w_eco52480, w_eco52481, w_eco52482, w_eco52483, w_eco52484, w_eco52485, w_eco52486, w_eco52487, w_eco52488, w_eco52489, w_eco52490, w_eco52491, w_eco52492, w_eco52493, w_eco52494, w_eco52495, w_eco52496, w_eco52497, w_eco52498, w_eco52499, w_eco52500, w_eco52501, w_eco52502, w_eco52503, w_eco52504, w_eco52505, w_eco52506, w_eco52507, w_eco52508, w_eco52509, w_eco52510, w_eco52511, w_eco52512, w_eco52513, w_eco52514, w_eco52515, w_eco52516, w_eco52517, w_eco52518, w_eco52519, w_eco52520, w_eco52521, w_eco52522, w_eco52523, w_eco52524, w_eco52525, w_eco52526, w_eco52527, w_eco52528, w_eco52529, w_eco52530, w_eco52531, w_eco52532, w_eco52533, w_eco52534, w_eco52535, w_eco52536, w_eco52537, w_eco52538, w_eco52539, w_eco52540, w_eco52541, w_eco52542, w_eco52543, w_eco52544, w_eco52545, w_eco52546, w_eco52547, w_eco52548, w_eco52549, w_eco52550, w_eco52551, w_eco52552, w_eco52553, w_eco52554, w_eco52555, w_eco52556, w_eco52557, w_eco52558, w_eco52559, w_eco52560, w_eco52561, w_eco52562, w_eco52563, w_eco52564, w_eco52565, w_eco52566, w_eco52567, w_eco52568, w_eco52569, w_eco52570, w_eco52571, w_eco52572, w_eco52573, w_eco52574, w_eco52575, w_eco52576, w_eco52577, w_eco52578, w_eco52579, w_eco52580, w_eco52581, w_eco52582, w_eco52583, w_eco52584, w_eco52585, w_eco52586, w_eco52587, w_eco52588, w_eco52589, w_eco52590, w_eco52591, w_eco52592, w_eco52593, w_eco52594, w_eco52595, w_eco52596, w_eco52597, w_eco52598, w_eco52599, w_eco52600, w_eco52601, w_eco52602, w_eco52603, w_eco52604, w_eco52605, w_eco52606, w_eco52607, w_eco52608, w_eco52609, w_eco52610, w_eco52611, w_eco52612, w_eco52613, w_eco52614, w_eco52615, w_eco52616, w_eco52617, w_eco52618, w_eco52619, w_eco52620, w_eco52621, w_eco52622, w_eco52623, w_eco52624, w_eco52625, w_eco52626, w_eco52627, w_eco52628, w_eco52629, w_eco52630, w_eco52631, w_eco52632, w_eco52633, w_eco52634, w_eco52635, w_eco52636, w_eco52637, w_eco52638, w_eco52639, w_eco52640, w_eco52641, w_eco52642, w_eco52643, w_eco52644, w_eco52645, w_eco52646, w_eco52647, w_eco52648, w_eco52649, w_eco52650, w_eco52651, w_eco52652, w_eco52653, w_eco52654, w_eco52655, w_eco52656, w_eco52657, w_eco52658, w_eco52659, w_eco52660, w_eco52661, w_eco52662, w_eco52663, w_eco52664, w_eco52665, w_eco52666, w_eco52667, w_eco52668, w_eco52669, w_eco52670, w_eco52671, w_eco52672, w_eco52673, w_eco52674, w_eco52675, w_eco52676, w_eco52677, w_eco52678, w_eco52679, w_eco52680, w_eco52681, w_eco52682, w_eco52683, w_eco52684, w_eco52685, w_eco52686, w_eco52687, w_eco52688, w_eco52689, w_eco52690, w_eco52691, w_eco52692, w_eco52693, w_eco52694, w_eco52695, w_eco52696, w_eco52697, w_eco52698, w_eco52699, w_eco52700, w_eco52701, w_eco52702, w_eco52703, w_eco52704, w_eco52705, w_eco52706, w_eco52707, w_eco52708, w_eco52709, w_eco52710, w_eco52711, w_eco52712, w_eco52713, w_eco52714, w_eco52715, w_eco52716, w_eco52717, w_eco52718, w_eco52719, w_eco52720, w_eco52721, w_eco52722, w_eco52723, w_eco52724, w_eco52725, w_eco52726, w_eco52727, w_eco52728, w_eco52729, w_eco52730, w_eco52731, w_eco52732, w_eco52733, w_eco52734, w_eco52735, w_eco52736, w_eco52737, w_eco52738, w_eco52739, w_eco52740, w_eco52741, w_eco52742, w_eco52743, w_eco52744, w_eco52745, w_eco52746, w_eco52747, w_eco52748, w_eco52749, w_eco52750, w_eco52751, w_eco52752, w_eco52753, w_eco52754, w_eco52755, w_eco52756, w_eco52757, w_eco52758, w_eco52759, w_eco52760, w_eco52761, w_eco52762, w_eco52763, w_eco52764, w_eco52765, w_eco52766, w_eco52767, w_eco52768, w_eco52769, w_eco52770, w_eco52771, w_eco52772, w_eco52773, w_eco52774, w_eco52775, w_eco52776, w_eco52777, w_eco52778, w_eco52779, w_eco52780, w_eco52781, w_eco52782, w_eco52783, w_eco52784, w_eco52785, w_eco52786, w_eco52787, w_eco52788, w_eco52789, w_eco52790, w_eco52791, w_eco52792, w_eco52793, w_eco52794, w_eco52795, w_eco52796, w_eco52797, w_eco52798, w_eco52799, w_eco52800, w_eco52801, w_eco52802, w_eco52803, w_eco52804, w_eco52805, w_eco52806, w_eco52807, w_eco52808, w_eco52809, w_eco52810, w_eco52811, w_eco52812, w_eco52813, w_eco52814, w_eco52815, w_eco52816, w_eco52817, w_eco52818, w_eco52819, w_eco52820, w_eco52821, w_eco52822, w_eco52823, w_eco52824, w_eco52825, w_eco52826, w_eco52827, w_eco52828, w_eco52829, w_eco52830, w_eco52831, w_eco52832, w_eco52833, w_eco52834, w_eco52835, w_eco52836, w_eco52837, w_eco52838, w_eco52839, w_eco52840, w_eco52841, w_eco52842, w_eco52843, w_eco52844, w_eco52845, w_eco52846, w_eco52847, w_eco52848, w_eco52849, w_eco52850, w_eco52851, w_eco52852, w_eco52853, w_eco52854, w_eco52855, w_eco52856, w_eco52857, w_eco52858, w_eco52859, w_eco52860, w_eco52861, w_eco52862, w_eco52863, w_eco52864, w_eco52865, w_eco52866, w_eco52867, w_eco52868, w_eco52869, w_eco52870, w_eco52871, w_eco52872, w_eco52873, w_eco52874, w_eco52875, w_eco52876, w_eco52877, w_eco52878, w_eco52879, w_eco52880, w_eco52881, w_eco52882, w_eco52883, w_eco52884, w_eco52885, w_eco52886, w_eco52887, w_eco52888, w_eco52889, w_eco52890, w_eco52891, w_eco52892, w_eco52893, w_eco52894, w_eco52895, w_eco52896, w_eco52897, w_eco52898, w_eco52899, w_eco52900, w_eco52901, w_eco52902, w_eco52903, w_eco52904, w_eco52905, w_eco52906, w_eco52907, w_eco52908, w_eco52909, w_eco52910, w_eco52911, w_eco52912, w_eco52913, w_eco52914, w_eco52915, w_eco52916, w_eco52917, w_eco52918, w_eco52919, w_eco52920, w_eco52921, w_eco52922, w_eco52923, w_eco52924, w_eco52925, w_eco52926, w_eco52927, w_eco52928, w_eco52929, w_eco52930, w_eco52931, w_eco52932, w_eco52933, w_eco52934, w_eco52935, w_eco52936, w_eco52937, w_eco52938, w_eco52939, w_eco52940, w_eco52941, w_eco52942, w_eco52943, w_eco52944, w_eco52945, w_eco52946, w_eco52947, w_eco52948, w_eco52949, w_eco52950, w_eco52951, w_eco52952, w_eco52953, w_eco52954, w_eco52955, w_eco52956, w_eco52957, w_eco52958, w_eco52959, w_eco52960, w_eco52961, w_eco52962, w_eco52963, w_eco52964, w_eco52965, w_eco52966, w_eco52967, w_eco52968, w_eco52969, w_eco52970, w_eco52971, w_eco52972, w_eco52973, w_eco52974, w_eco52975, w_eco52976, w_eco52977, w_eco52978, w_eco52979, w_eco52980, w_eco52981, w_eco52982, w_eco52983, w_eco52984, w_eco52985, w_eco52986, w_eco52987, w_eco52988, w_eco52989, w_eco52990, w_eco52991, w_eco52992, w_eco52993, w_eco52994, w_eco52995, w_eco52996, w_eco52997, w_eco52998, w_eco52999, w_eco53000, w_eco53001, w_eco53002, w_eco53003, w_eco53004, w_eco53005, w_eco53006, w_eco53007, w_eco53008, w_eco53009, w_eco53010, w_eco53011, w_eco53012, w_eco53013, w_eco53014, w_eco53015, w_eco53016, w_eco53017, w_eco53018, w_eco53019, w_eco53020, w_eco53021, w_eco53022, w_eco53023, w_eco53024, w_eco53025, w_eco53026, w_eco53027, w_eco53028, w_eco53029, w_eco53030, w_eco53031, w_eco53032, w_eco53033, w_eco53034, w_eco53035, w_eco53036, w_eco53037, w_eco53038, w_eco53039, w_eco53040, w_eco53041, w_eco53042, w_eco53043, w_eco53044, w_eco53045, w_eco53046, w_eco53047, w_eco53048, w_eco53049, w_eco53050, w_eco53051, w_eco53052, w_eco53053, w_eco53054, w_eco53055, w_eco53056, w_eco53057, w_eco53058, w_eco53059, w_eco53060, w_eco53061, w_eco53062, w_eco53063, w_eco53064, w_eco53065, w_eco53066, w_eco53067, w_eco53068, w_eco53069, w_eco53070, w_eco53071, w_eco53072, w_eco53073, w_eco53074, w_eco53075, w_eco53076, w_eco53077, w_eco53078, w_eco53079, w_eco53080, w_eco53081, w_eco53082, w_eco53083, w_eco53084, w_eco53085, w_eco53086, w_eco53087, w_eco53088, w_eco53089, w_eco53090, w_eco53091, w_eco53092, w_eco53093, w_eco53094, w_eco53095, w_eco53096, w_eco53097, w_eco53098, w_eco53099, w_eco53100, w_eco53101, w_eco53102, w_eco53103, w_eco53104, w_eco53105, w_eco53106, w_eco53107, w_eco53108, w_eco53109, w_eco53110, w_eco53111, w_eco53112, w_eco53113, w_eco53114, w_eco53115, w_eco53116, w_eco53117, w_eco53118, w_eco53119, w_eco53120, w_eco53121, w_eco53122, w_eco53123, w_eco53124, w_eco53125, w_eco53126, w_eco53127, w_eco53128, w_eco53129, w_eco53130, w_eco53131, w_eco53132, w_eco53133, w_eco53134, w_eco53135, w_eco53136, w_eco53137, w_eco53138, w_eco53139, w_eco53140, w_eco53141, w_eco53142, w_eco53143, w_eco53144, w_eco53145, w_eco53146, w_eco53147, w_eco53148, w_eco53149, w_eco53150, w_eco53151, w_eco53152, w_eco53153, w_eco53154, w_eco53155, w_eco53156, w_eco53157, w_eco53158, w_eco53159, w_eco53160, w_eco53161, w_eco53162, w_eco53163, w_eco53164, w_eco53165, w_eco53166, w_eco53167, w_eco53168, w_eco53169, w_eco53170, w_eco53171, w_eco53172, w_eco53173, w_eco53174, w_eco53175, w_eco53176, w_eco53177, w_eco53178, w_eco53179, w_eco53180, w_eco53181, w_eco53182, w_eco53183, w_eco53184, w_eco53185, w_eco53186, w_eco53187, w_eco53188, w_eco53189, w_eco53190, w_eco53191, w_eco53192, w_eco53193, w_eco53194, w_eco53195, w_eco53196, w_eco53197, w_eco53198, w_eco53199, w_eco53200, w_eco53201, w_eco53202, w_eco53203, w_eco53204, w_eco53205, w_eco53206, w_eco53207, w_eco53208, w_eco53209, w_eco53210, w_eco53211, w_eco53212, w_eco53213, w_eco53214, w_eco53215, w_eco53216, w_eco53217, w_eco53218, w_eco53219, w_eco53220, w_eco53221, w_eco53222, w_eco53223, w_eco53224, w_eco53225, w_eco53226, w_eco53227, w_eco53228, w_eco53229, w_eco53230, w_eco53231, w_eco53232, w_eco53233, w_eco53234, w_eco53235, w_eco53236, w_eco53237, w_eco53238, w_eco53239, w_eco53240, w_eco53241, w_eco53242, w_eco53243, w_eco53244, w_eco53245, w_eco53246, w_eco53247, w_eco53248, w_eco53249, w_eco53250, w_eco53251, w_eco53252, w_eco53253, w_eco53254, w_eco53255, w_eco53256, w_eco53257, w_eco53258, w_eco53259, w_eco53260, w_eco53261, w_eco53262, w_eco53263, w_eco53264, w_eco53265, w_eco53266, w_eco53267, w_eco53268, w_eco53269, w_eco53270, w_eco53271, w_eco53272, w_eco53273, w_eco53274, w_eco53275, w_eco53276, w_eco53277, w_eco53278, w_eco53279, w_eco53280, w_eco53281, w_eco53282, w_eco53283, w_eco53284, w_eco53285, w_eco53286, w_eco53287, w_eco53288, w_eco53289, w_eco53290, w_eco53291, w_eco53292, w_eco53293, w_eco53294, w_eco53295, w_eco53296, w_eco53297, w_eco53298, w_eco53299, w_eco53300, w_eco53301, w_eco53302, w_eco53303, w_eco53304, w_eco53305, w_eco53306, w_eco53307, w_eco53308, w_eco53309, w_eco53310, w_eco53311, w_eco53312, w_eco53313, w_eco53314, w_eco53315, w_eco53316, w_eco53317, w_eco53318, w_eco53319, w_eco53320, w_eco53321, w_eco53322, w_eco53323, w_eco53324, w_eco53325, w_eco53326, w_eco53327, w_eco53328, w_eco53329, w_eco53330, w_eco53331, w_eco53332, w_eco53333, w_eco53334, w_eco53335, w_eco53336, w_eco53337, w_eco53338, w_eco53339, w_eco53340, w_eco53341, w_eco53342, w_eco53343, w_eco53344, w_eco53345, w_eco53346, w_eco53347, w_eco53348, w_eco53349, w_eco53350, w_eco53351, w_eco53352, w_eco53353, w_eco53354, w_eco53355, w_eco53356, w_eco53357, w_eco53358, w_eco53359, w_eco53360, w_eco53361, w_eco53362, w_eco53363, w_eco53364, w_eco53365, w_eco53366, w_eco53367, w_eco53368, w_eco53369, w_eco53370, w_eco53371, w_eco53372, w_eco53373, w_eco53374, w_eco53375, w_eco53376, w_eco53377, w_eco53378, w_eco53379, w_eco53380, w_eco53381, w_eco53382, w_eco53383, w_eco53384, w_eco53385, w_eco53386, w_eco53387, w_eco53388, w_eco53389, w_eco53390, w_eco53391, w_eco53392, w_eco53393, w_eco53394, w_eco53395, w_eco53396, w_eco53397, w_eco53398, w_eco53399, w_eco53400, w_eco53401, w_eco53402, w_eco53403, w_eco53404, w_eco53405, w_eco53406, w_eco53407, w_eco53408, w_eco53409, w_eco53410, w_eco53411, w_eco53412, w_eco53413, w_eco53414, w_eco53415, w_eco53416, w_eco53417, w_eco53418, w_eco53419, w_eco53420, w_eco53421, w_eco53422, w_eco53423, w_eco53424, w_eco53425, w_eco53426, w_eco53427, w_eco53428, w_eco53429, w_eco53430, w_eco53431, w_eco53432, w_eco53433, w_eco53434, w_eco53435, w_eco53436, w_eco53437, w_eco53438, w_eco53439, w_eco53440, w_eco53441, w_eco53442, w_eco53443, w_eco53444, w_eco53445, w_eco53446, w_eco53447, w_eco53448, w_eco53449, w_eco53450, w_eco53451, w_eco53452, w_eco53453, w_eco53454, w_eco53455, w_eco53456, w_eco53457, w_eco53458, w_eco53459, w_eco53460, w_eco53461, w_eco53462, w_eco53463, w_eco53464, w_eco53465, w_eco53466, w_eco53467, w_eco53468, w_eco53469, w_eco53470, w_eco53471, w_eco53472, w_eco53473, w_eco53474, w_eco53475, w_eco53476, w_eco53477, w_eco53478, w_eco53479, w_eco53480, w_eco53481, w_eco53482, w_eco53483, w_eco53484, w_eco53485, w_eco53486, w_eco53487, w_eco53488, w_eco53489, w_eco53490, w_eco53491, w_eco53492, w_eco53493, w_eco53494, w_eco53495, w_eco53496, w_eco53497, w_eco53498, w_eco53499, w_eco53500, w_eco53501, w_eco53502, w_eco53503, w_eco53504, w_eco53505, w_eco53506, w_eco53507, w_eco53508, w_eco53509, w_eco53510, w_eco53511, w_eco53512, w_eco53513, w_eco53514, w_eco53515, w_eco53516, w_eco53517, w_eco53518, w_eco53519, w_eco53520, w_eco53521, w_eco53522, w_eco53523, w_eco53524, w_eco53525, w_eco53526, w_eco53527, w_eco53528, w_eco53529, w_eco53530, w_eco53531, w_eco53532, w_eco53533, w_eco53534, w_eco53535, w_eco53536, w_eco53537, w_eco53538, w_eco53539, w_eco53540, w_eco53541, w_eco53542, w_eco53543, w_eco53544, w_eco53545, w_eco53546, w_eco53547, w_eco53548, w_eco53549, w_eco53550, w_eco53551, w_eco53552, w_eco53553, w_eco53554, w_eco53555, w_eco53556, w_eco53557, w_eco53558, w_eco53559, w_eco53560, w_eco53561, w_eco53562, w_eco53563, w_eco53564, w_eco53565, w_eco53566, w_eco53567, w_eco53568, w_eco53569, w_eco53570, w_eco53571, w_eco53572, w_eco53573, w_eco53574, w_eco53575, w_eco53576, w_eco53577, w_eco53578, w_eco53579, w_eco53580, w_eco53581, w_eco53582, w_eco53583, w_eco53584, w_eco53585, w_eco53586, w_eco53587, w_eco53588, w_eco53589, w_eco53590, w_eco53591, w_eco53592, w_eco53593, w_eco53594, w_eco53595, w_eco53596, w_eco53597, w_eco53598, w_eco53599, w_eco53600, w_eco53601, w_eco53602, w_eco53603, w_eco53604, w_eco53605, w_eco53606, w_eco53607, w_eco53608, w_eco53609, w_eco53610, w_eco53611, w_eco53612, w_eco53613, w_eco53614, w_eco53615, w_eco53616, w_eco53617, w_eco53618, w_eco53619, w_eco53620, w_eco53621, w_eco53622, w_eco53623, w_eco53624, w_eco53625, w_eco53626, w_eco53627, w_eco53628, w_eco53629, w_eco53630, w_eco53631, w_eco53632, w_eco53633, w_eco53634, w_eco53635, w_eco53636, w_eco53637, w_eco53638, w_eco53639, w_eco53640, w_eco53641, w_eco53642, w_eco53643, w_eco53644, w_eco53645, w_eco53646, w_eco53647, w_eco53648, w_eco53649, w_eco53650, w_eco53651, w_eco53652, w_eco53653, w_eco53654, w_eco53655, w_eco53656, w_eco53657, w_eco53658, w_eco53659, w_eco53660, w_eco53661, w_eco53662, w_eco53663, w_eco53664, w_eco53665, w_eco53666, w_eco53667, w_eco53668, w_eco53669, w_eco53670, w_eco53671, w_eco53672, w_eco53673, w_eco53674, w_eco53675, w_eco53676, w_eco53677, w_eco53678, w_eco53679, w_eco53680, w_eco53681, w_eco53682, w_eco53683, w_eco53684, w_eco53685, w_eco53686, w_eco53687, w_eco53688, w_eco53689, w_eco53690, w_eco53691, w_eco53692, w_eco53693, w_eco53694, w_eco53695, w_eco53696, w_eco53697, w_eco53698, w_eco53699, w_eco53700, w_eco53701, w_eco53702, w_eco53703, w_eco53704, w_eco53705, w_eco53706, w_eco53707, w_eco53708, w_eco53709, w_eco53710, w_eco53711, w_eco53712, w_eco53713, w_eco53714, w_eco53715, w_eco53716, w_eco53717, w_eco53718, w_eco53719, w_eco53720, w_eco53721, w_eco53722, w_eco53723, w_eco53724, w_eco53725, w_eco53726, w_eco53727, w_eco53728, w_eco53729, w_eco53730, w_eco53731, w_eco53732, w_eco53733, w_eco53734, w_eco53735, w_eco53736, w_eco53737, w_eco53738, w_eco53739, w_eco53740, w_eco53741, w_eco53742, w_eco53743, w_eco53744, w_eco53745, w_eco53746, w_eco53747, w_eco53748, w_eco53749, w_eco53750, w_eco53751, w_eco53752, w_eco53753, w_eco53754, w_eco53755, w_eco53756, w_eco53757, w_eco53758, w_eco53759, w_eco53760, w_eco53761, w_eco53762, w_eco53763, w_eco53764, w_eco53765, w_eco53766, w_eco53767, w_eco53768, w_eco53769, w_eco53770, w_eco53771, w_eco53772, w_eco53773, w_eco53774, w_eco53775, w_eco53776, w_eco53777, w_eco53778, w_eco53779, w_eco53780, w_eco53781, w_eco53782, w_eco53783, w_eco53784, w_eco53785, w_eco53786, w_eco53787, w_eco53788, w_eco53789, w_eco53790, w_eco53791, w_eco53792, w_eco53793, w_eco53794, w_eco53795, w_eco53796, w_eco53797, w_eco53798, w_eco53799, w_eco53800, w_eco53801, w_eco53802, w_eco53803, w_eco53804, w_eco53805, w_eco53806, w_eco53807, w_eco53808, w_eco53809, w_eco53810, w_eco53811, w_eco53812, w_eco53813, w_eco53814, w_eco53815, w_eco53816, w_eco53817, w_eco53818, w_eco53819, w_eco53820, w_eco53821, w_eco53822, w_eco53823, w_eco53824, w_eco53825, w_eco53826, w_eco53827, w_eco53828, w_eco53829, w_eco53830, w_eco53831, w_eco53832, w_eco53833, w_eco53834, w_eco53835, w_eco53836, w_eco53837, w_eco53838, w_eco53839, w_eco53840, w_eco53841, w_eco53842, w_eco53843, w_eco53844, w_eco53845, w_eco53846, w_eco53847, w_eco53848, w_eco53849, w_eco53850, w_eco53851, w_eco53852, w_eco53853, w_eco53854, w_eco53855, w_eco53856, w_eco53857, w_eco53858, w_eco53859, w_eco53860, w_eco53861, w_eco53862, w_eco53863, w_eco53864, w_eco53865, w_eco53866, w_eco53867, w_eco53868, w_eco53869, w_eco53870, w_eco53871, w_eco53872, w_eco53873, w_eco53874, w_eco53875, w_eco53876, w_eco53877, w_eco53878, w_eco53879, w_eco53880, w_eco53881, w_eco53882, w_eco53883, w_eco53884, w_eco53885, w_eco53886, w_eco53887, w_eco53888, w_eco53889, w_eco53890, w_eco53891, w_eco53892, w_eco53893, w_eco53894, w_eco53895, w_eco53896, w_eco53897, w_eco53898, w_eco53899, w_eco53900, w_eco53901, w_eco53902, w_eco53903, w_eco53904, w_eco53905, w_eco53906, w_eco53907, w_eco53908, w_eco53909, w_eco53910, w_eco53911, w_eco53912, w_eco53913, w_eco53914, w_eco53915, w_eco53916, w_eco53917, w_eco53918, w_eco53919, w_eco53920, w_eco53921, w_eco53922, w_eco53923, w_eco53924, w_eco53925, w_eco53926, w_eco53927, w_eco53928, w_eco53929, w_eco53930, w_eco53931, w_eco53932, w_eco53933, w_eco53934, w_eco53935, w_eco53936, w_eco53937, w_eco53938, w_eco53939, w_eco53940, w_eco53941, w_eco53942, w_eco53943, w_eco53944, w_eco53945, w_eco53946, w_eco53947, w_eco53948, w_eco53949, w_eco53950, w_eco53951, w_eco53952, w_eco53953, w_eco53954, w_eco53955, w_eco53956, w_eco53957, w_eco53958, w_eco53959, w_eco53960, w_eco53961, w_eco53962, w_eco53963, w_eco53964, w_eco53965, w_eco53966, w_eco53967, w_eco53968, w_eco53969, w_eco53970, w_eco53971, w_eco53972, w_eco53973, w_eco53974, w_eco53975, w_eco53976, w_eco53977, w_eco53978, w_eco53979, w_eco53980, w_eco53981, w_eco53982, w_eco53983, w_eco53984, w_eco53985, w_eco53986, w_eco53987, w_eco53988, w_eco53989, w_eco53990, w_eco53991, w_eco53992, w_eco53993, w_eco53994, w_eco53995, w_eco53996, w_eco53997, w_eco53998, w_eco53999, w_eco54000, w_eco54001, w_eco54002, w_eco54003, w_eco54004, w_eco54005, w_eco54006, w_eco54007, w_eco54008, w_eco54009, w_eco54010, w_eco54011, w_eco54012, w_eco54013, w_eco54014, w_eco54015, w_eco54016, w_eco54017, w_eco54018, w_eco54019, w_eco54020, w_eco54021, w_eco54022, w_eco54023, w_eco54024, w_eco54025, w_eco54026, w_eco54027, w_eco54028, w_eco54029, w_eco54030, w_eco54031, w_eco54032, w_eco54033, w_eco54034, w_eco54035, w_eco54036, w_eco54037, w_eco54038, w_eco54039, w_eco54040, w_eco54041, w_eco54042, w_eco54043, w_eco54044, w_eco54045, w_eco54046, w_eco54047, w_eco54048, w_eco54049, w_eco54050, w_eco54051, w_eco54052, w_eco54053, w_eco54054, w_eco54055, w_eco54056, w_eco54057, w_eco54058, w_eco54059, w_eco54060, w_eco54061, w_eco54062, w_eco54063, w_eco54064, w_eco54065, w_eco54066, w_eco54067, w_eco54068, w_eco54069, w_eco54070, w_eco54071, w_eco54072, w_eco54073, w_eco54074, w_eco54075, w_eco54076, w_eco54077, w_eco54078, w_eco54079, w_eco54080, w_eco54081, w_eco54082, w_eco54083, w_eco54084, w_eco54085, w_eco54086, w_eco54087, w_eco54088, w_eco54089, w_eco54090, w_eco54091, w_eco54092, w_eco54093, w_eco54094, w_eco54095, w_eco54096, w_eco54097, w_eco54098, w_eco54099, w_eco54100, w_eco54101, w_eco54102, w_eco54103, w_eco54104, w_eco54105, w_eco54106, w_eco54107, w_eco54108, w_eco54109, w_eco54110, w_eco54111, w_eco54112, w_eco54113, w_eco54114, w_eco54115, w_eco54116, w_eco54117, w_eco54118, w_eco54119, w_eco54120, w_eco54121, w_eco54122, w_eco54123, w_eco54124, w_eco54125, w_eco54126, w_eco54127, w_eco54128, w_eco54129, w_eco54130, w_eco54131, w_eco54132, w_eco54133, w_eco54134, w_eco54135, w_eco54136, w_eco54137, w_eco54138, w_eco54139, w_eco54140, w_eco54141, w_eco54142, w_eco54143, w_eco54144, w_eco54145, w_eco54146, w_eco54147, w_eco54148, w_eco54149, w_eco54150, w_eco54151, w_eco54152, w_eco54153, w_eco54154, w_eco54155, w_eco54156, w_eco54157, w_eco54158, w_eco54159, w_eco54160, w_eco54161, w_eco54162, w_eco54163, w_eco54164, w_eco54165, w_eco54166, w_eco54167, w_eco54168, w_eco54169, w_eco54170, w_eco54171, w_eco54172, w_eco54173, w_eco54174, w_eco54175, w_eco54176, w_eco54177, w_eco54178, w_eco54179, w_eco54180, w_eco54181, w_eco54182, w_eco54183, w_eco54184, w_eco54185, w_eco54186, w_eco54187, w_eco54188, w_eco54189, w_eco54190, w_eco54191, w_eco54192, w_eco54193, w_eco54194, w_eco54195, w_eco54196, w_eco54197, w_eco54198, w_eco54199, w_eco54200, w_eco54201, w_eco54202, w_eco54203, w_eco54204, w_eco54205, w_eco54206, w_eco54207, w_eco54208, w_eco54209, w_eco54210, w_eco54211, w_eco54212, w_eco54213, w_eco54214, w_eco54215, w_eco54216, w_eco54217, w_eco54218, w_eco54219, w_eco54220, w_eco54221, w_eco54222, w_eco54223, w_eco54224, w_eco54225, w_eco54226, w_eco54227, w_eco54228, w_eco54229, w_eco54230, w_eco54231, w_eco54232, w_eco54233, w_eco54234, w_eco54235, w_eco54236, w_eco54237, w_eco54238, w_eco54239, w_eco54240, w_eco54241, w_eco54242, w_eco54243, w_eco54244, w_eco54245, w_eco54246, w_eco54247, w_eco54248, w_eco54249, w_eco54250, w_eco54251, w_eco54252, w_eco54253, w_eco54254, w_eco54255, w_eco54256, w_eco54257, w_eco54258, w_eco54259, w_eco54260, w_eco54261, w_eco54262, w_eco54263, w_eco54264, w_eco54265, w_eco54266, w_eco54267, w_eco54268, w_eco54269, w_eco54270, w_eco54271, w_eco54272, w_eco54273, w_eco54274, w_eco54275, w_eco54276, w_eco54277, w_eco54278, w_eco54279, w_eco54280, w_eco54281, w_eco54282, w_eco54283, w_eco54284, w_eco54285, w_eco54286, w_eco54287, w_eco54288, w_eco54289, w_eco54290, w_eco54291, w_eco54292, w_eco54293, w_eco54294, w_eco54295, w_eco54296, w_eco54297, w_eco54298, w_eco54299, w_eco54300, w_eco54301, w_eco54302, w_eco54303, w_eco54304, w_eco54305, w_eco54306, w_eco54307, w_eco54308, w_eco54309, w_eco54310, w_eco54311, w_eco54312, w_eco54313, w_eco54314, w_eco54315, w_eco54316, w_eco54317, w_eco54318, w_eco54319, w_eco54320, w_eco54321, w_eco54322, w_eco54323, w_eco54324, w_eco54325, w_eco54326, w_eco54327, w_eco54328, w_eco54329, w_eco54330, w_eco54331, w_eco54332, w_eco54333, w_eco54334, w_eco54335, w_eco54336, w_eco54337, w_eco54338, w_eco54339, w_eco54340, w_eco54341, w_eco54342, w_eco54343, w_eco54344, w_eco54345, w_eco54346, w_eco54347, w_eco54348, w_eco54349, w_eco54350, w_eco54351, w_eco54352, w_eco54353, w_eco54354, w_eco54355, w_eco54356, w_eco54357, w_eco54358, w_eco54359, w_eco54360, w_eco54361, w_eco54362, w_eco54363, w_eco54364, w_eco54365, w_eco54366, w_eco54367, w_eco54368, w_eco54369, w_eco54370, w_eco54371, w_eco54372, w_eco54373, w_eco54374, w_eco54375, w_eco54376, w_eco54377, w_eco54378, w_eco54379, w_eco54380, w_eco54381, w_eco54382, w_eco54383, w_eco54384, w_eco54385, w_eco54386, w_eco54387, w_eco54388, w_eco54389, w_eco54390, w_eco54391, w_eco54392, w_eco54393, w_eco54394, w_eco54395, w_eco54396, w_eco54397, w_eco54398, w_eco54399, w_eco54400, w_eco54401, w_eco54402, w_eco54403, w_eco54404, w_eco54405, w_eco54406, w_eco54407, w_eco54408, w_eco54409, w_eco54410, w_eco54411, w_eco54412, w_eco54413, w_eco54414, w_eco54415, w_eco54416, w_eco54417, w_eco54418, w_eco54419, w_eco54420, w_eco54421, w_eco54422, w_eco54423, w_eco54424, w_eco54425, w_eco54426, w_eco54427, w_eco54428, w_eco54429, w_eco54430, w_eco54431, w_eco54432, w_eco54433, w_eco54434, w_eco54435, w_eco54436, w_eco54437, w_eco54438, w_eco54439, w_eco54440, w_eco54441, w_eco54442, w_eco54443, w_eco54444, w_eco54445, w_eco54446, w_eco54447, w_eco54448, w_eco54449, w_eco54450, w_eco54451, w_eco54452, w_eco54453, w_eco54454, w_eco54455, w_eco54456, w_eco54457, w_eco54458, w_eco54459, w_eco54460, w_eco54461, w_eco54462, w_eco54463, w_eco54464, w_eco54465, w_eco54466, w_eco54467, w_eco54468, w_eco54469, w_eco54470, w_eco54471, w_eco54472, w_eco54473, w_eco54474, w_eco54475, w_eco54476, w_eco54477, w_eco54478, w_eco54479, w_eco54480, w_eco54481, w_eco54482, w_eco54483, w_eco54484, w_eco54485, w_eco54486, w_eco54487, w_eco54488, w_eco54489, w_eco54490, w_eco54491, w_eco54492, w_eco54493, w_eco54494, w_eco54495, w_eco54496, w_eco54497, w_eco54498, w_eco54499, w_eco54500, w_eco54501, w_eco54502, w_eco54503, w_eco54504, w_eco54505, w_eco54506, w_eco54507, w_eco54508, w_eco54509, w_eco54510, w_eco54511, w_eco54512, w_eco54513, w_eco54514, w_eco54515, w_eco54516, w_eco54517, w_eco54518, w_eco54519, w_eco54520, w_eco54521, w_eco54522, w_eco54523, w_eco54524, w_eco54525, w_eco54526, w_eco54527, w_eco54528, w_eco54529, w_eco54530, w_eco54531, w_eco54532, w_eco54533, w_eco54534, w_eco54535, w_eco54536, w_eco54537, w_eco54538, w_eco54539, w_eco54540, w_eco54541, w_eco54542, w_eco54543, w_eco54544, w_eco54545, w_eco54546, w_eco54547, w_eco54548, w_eco54549, w_eco54550, w_eco54551, w_eco54552, w_eco54553, w_eco54554, w_eco54555, w_eco54556, w_eco54557, w_eco54558, w_eco54559, w_eco54560, w_eco54561, w_eco54562, w_eco54563, w_eco54564, w_eco54565, w_eco54566, w_eco54567, w_eco54568, w_eco54569, w_eco54570, w_eco54571, w_eco54572, w_eco54573, w_eco54574, w_eco54575, w_eco54576, w_eco54577, w_eco54578, w_eco54579, w_eco54580, w_eco54581, w_eco54582, w_eco54583, w_eco54584, w_eco54585, w_eco54586, w_eco54587, w_eco54588, w_eco54589, w_eco54590, w_eco54591, w_eco54592, w_eco54593, w_eco54594, w_eco54595, w_eco54596, w_eco54597, w_eco54598, w_eco54599, w_eco54600, w_eco54601, w_eco54602, w_eco54603, w_eco54604, w_eco54605, w_eco54606, w_eco54607, w_eco54608, w_eco54609, w_eco54610, w_eco54611, w_eco54612, w_eco54613, w_eco54614, w_eco54615, w_eco54616, w_eco54617, w_eco54618, w_eco54619, w_eco54620, w_eco54621, w_eco54622, w_eco54623, w_eco54624, w_eco54625, w_eco54626, w_eco54627, w_eco54628, w_eco54629, w_eco54630, w_eco54631, w_eco54632, w_eco54633, w_eco54634, w_eco54635, w_eco54636, w_eco54637, w_eco54638, w_eco54639, w_eco54640, w_eco54641, w_eco54642, w_eco54643, w_eco54644, w_eco54645, w_eco54646, w_eco54647, w_eco54648, w_eco54649, w_eco54650, w_eco54651, w_eco54652, w_eco54653, w_eco54654, w_eco54655, w_eco54656, w_eco54657, w_eco54658, w_eco54659, w_eco54660, w_eco54661, w_eco54662, w_eco54663, w_eco54664, w_eco54665, w_eco54666, w_eco54667, w_eco54668, w_eco54669, w_eco54670, w_eco54671, w_eco54672, w_eco54673, w_eco54674, w_eco54675, w_eco54676, w_eco54677, w_eco54678, w_eco54679, w_eco54680, w_eco54681, w_eco54682, w_eco54683, w_eco54684, w_eco54685, w_eco54686, w_eco54687, w_eco54688, w_eco54689, w_eco54690, w_eco54691, w_eco54692, w_eco54693, w_eco54694, w_eco54695, w_eco54696, w_eco54697, w_eco54698, w_eco54699, w_eco54700, w_eco54701, w_eco54702, w_eco54703, w_eco54704, w_eco54705, w_eco54706, w_eco54707, w_eco54708, w_eco54709, w_eco54710, w_eco54711, w_eco54712, w_eco54713, w_eco54714, w_eco54715, w_eco54716, w_eco54717, w_eco54718, w_eco54719, w_eco54720, w_eco54721, w_eco54722, w_eco54723, w_eco54724, w_eco54725, w_eco54726, w_eco54727, w_eco54728, w_eco54729, w_eco54730, w_eco54731, w_eco54732, w_eco54733, w_eco54734, w_eco54735, w_eco54736, w_eco54737, w_eco54738, w_eco54739, w_eco54740, w_eco54741, w_eco54742, w_eco54743, w_eco54744, w_eco54745, w_eco54746, w_eco54747, w_eco54748, w_eco54749, w_eco54750, w_eco54751, w_eco54752, w_eco54753, w_eco54754, w_eco54755, w_eco54756, w_eco54757, w_eco54758, w_eco54759, w_eco54760, w_eco54761, w_eco54762, w_eco54763, w_eco54764, w_eco54765, w_eco54766, w_eco54767, w_eco54768, w_eco54769, w_eco54770, w_eco54771, w_eco54772, w_eco54773, w_eco54774, w_eco54775, w_eco54776, w_eco54777, w_eco54778, w_eco54779, w_eco54780, w_eco54781, w_eco54782, w_eco54783, w_eco54784, w_eco54785, w_eco54786, w_eco54787, w_eco54788, w_eco54789, w_eco54790, w_eco54791, w_eco54792, w_eco54793, w_eco54794, w_eco54795, w_eco54796, w_eco54797, w_eco54798, w_eco54799, w_eco54800, w_eco54801, w_eco54802, w_eco54803, w_eco54804, w_eco54805, w_eco54806, w_eco54807, w_eco54808, w_eco54809, w_eco54810, w_eco54811, w_eco54812, w_eco54813, w_eco54814, w_eco54815, w_eco54816, w_eco54817, w_eco54818, w_eco54819, w_eco54820, w_eco54821, w_eco54822, w_eco54823, w_eco54824, w_eco54825, w_eco54826, w_eco54827, w_eco54828, w_eco54829, w_eco54830, w_eco54831, w_eco54832, w_eco54833, w_eco54834, w_eco54835, w_eco54836, w_eco54837, w_eco54838, w_eco54839, w_eco54840, w_eco54841, w_eco54842, w_eco54843, w_eco54844, w_eco54845, w_eco54846, w_eco54847, w_eco54848, w_eco54849, w_eco54850, w_eco54851, w_eco54852, w_eco54853, w_eco54854, w_eco54855, w_eco54856, w_eco54857, w_eco54858, w_eco54859, w_eco54860, w_eco54861, w_eco54862, w_eco54863, w_eco54864, w_eco54865, w_eco54866, w_eco54867, w_eco54868, w_eco54869, w_eco54870, w_eco54871, w_eco54872, w_eco54873, w_eco54874, w_eco54875, w_eco54876, w_eco54877, w_eco54878, w_eco54879, w_eco54880, w_eco54881, w_eco54882, w_eco54883, w_eco54884, w_eco54885, w_eco54886, w_eco54887, w_eco54888, w_eco54889, w_eco54890, w_eco54891, w_eco54892, w_eco54893, w_eco54894, w_eco54895, w_eco54896, w_eco54897, w_eco54898, w_eco54899, w_eco54900, w_eco54901, w_eco54902, w_eco54903, w_eco54904, w_eco54905, w_eco54906, w_eco54907, w_eco54908, w_eco54909, w_eco54910, w_eco54911, w_eco54912, w_eco54913, w_eco54914, w_eco54915, w_eco54916, w_eco54917, w_eco54918, w_eco54919, w_eco54920, w_eco54921, w_eco54922, w_eco54923, w_eco54924, w_eco54925, w_eco54926, w_eco54927, w_eco54928, w_eco54929, w_eco54930, w_eco54931, w_eco54932, w_eco54933, w_eco54934, w_eco54935, w_eco54936, w_eco54937, w_eco54938, w_eco54939, w_eco54940, w_eco54941, w_eco54942, w_eco54943, w_eco54944, w_eco54945, w_eco54946, w_eco54947, w_eco54948, w_eco54949, w_eco54950, w_eco54951, w_eco54952, w_eco54953, w_eco54954, w_eco54955, w_eco54956, w_eco54957, w_eco54958, w_eco54959, w_eco54960, w_eco54961, w_eco54962, w_eco54963, w_eco54964, w_eco54965, w_eco54966, w_eco54967, w_eco54968, w_eco54969, w_eco54970, w_eco54971, w_eco54972, w_eco54973, w_eco54974, w_eco54975, w_eco54976, w_eco54977, w_eco54978, w_eco54979, w_eco54980, w_eco54981, w_eco54982, w_eco54983, w_eco54984, w_eco54985, w_eco54986, w_eco54987, w_eco54988, w_eco54989, w_eco54990, w_eco54991, w_eco54992, w_eco54993, w_eco54994, w_eco54995, w_eco54996, w_eco54997, w_eco54998, w_eco54999, w_eco55000, w_eco55001, w_eco55002, w_eco55003, w_eco55004, w_eco55005, w_eco55006, w_eco55007, w_eco55008, w_eco55009, w_eco55010, w_eco55011, w_eco55012, w_eco55013, w_eco55014, w_eco55015, w_eco55016, w_eco55017, w_eco55018, w_eco55019, w_eco55020, w_eco55021, w_eco55022, w_eco55023, w_eco55024, w_eco55025, w_eco55026, w_eco55027, w_eco55028, w_eco55029, w_eco55030, w_eco55031, w_eco55032, w_eco55033, w_eco55034, w_eco55035, w_eco55036, w_eco55037, w_eco55038, w_eco55039, w_eco55040, w_eco55041, w_eco55042, w_eco55043, w_eco55044, w_eco55045, w_eco55046, w_eco55047, w_eco55048, w_eco55049, w_eco55050, w_eco55051, w_eco55052, w_eco55053, w_eco55054, w_eco55055, w_eco55056, w_eco55057, w_eco55058, w_eco55059, w_eco55060, w_eco55061, w_eco55062, w_eco55063, w_eco55064, w_eco55065, w_eco55066, w_eco55067, w_eco55068, w_eco55069, w_eco55070, w_eco55071, w_eco55072, w_eco55073, w_eco55074, w_eco55075, w_eco55076, w_eco55077, w_eco55078, w_eco55079, w_eco55080, w_eco55081, w_eco55082, w_eco55083, w_eco55084, w_eco55085, w_eco55086, w_eco55087, w_eco55088, w_eco55089, w_eco55090, w_eco55091, w_eco55092, w_eco55093, w_eco55094, w_eco55095, w_eco55096, w_eco55097, w_eco55098, w_eco55099, w_eco55100, w_eco55101, w_eco55102, w_eco55103, w_eco55104, w_eco55105, w_eco55106, w_eco55107, w_eco55108, w_eco55109, w_eco55110, w_eco55111, w_eco55112, w_eco55113, w_eco55114, w_eco55115, w_eco55116, w_eco55117, w_eco55118, w_eco55119, w_eco55120, w_eco55121, w_eco55122, w_eco55123, w_eco55124, w_eco55125, w_eco55126, w_eco55127, w_eco55128, w_eco55129, w_eco55130, w_eco55131, w_eco55132, w_eco55133, w_eco55134, w_eco55135, w_eco55136, w_eco55137, w_eco55138, w_eco55139, w_eco55140, w_eco55141, w_eco55142, w_eco55143, w_eco55144, w_eco55145, w_eco55146, w_eco55147, w_eco55148, w_eco55149, w_eco55150, w_eco55151, w_eco55152, w_eco55153, w_eco55154, w_eco55155, w_eco55156, w_eco55157, w_eco55158, w_eco55159, w_eco55160, w_eco55161, w_eco55162, w_eco55163, w_eco55164, w_eco55165, w_eco55166, w_eco55167, w_eco55168, w_eco55169, w_eco55170, w_eco55171, w_eco55172, w_eco55173, w_eco55174, w_eco55175, w_eco55176, w_eco55177, w_eco55178, w_eco55179, w_eco55180, w_eco55181, w_eco55182, w_eco55183, w_eco55184, w_eco55185, w_eco55186, w_eco55187, w_eco55188, w_eco55189, w_eco55190, w_eco55191, w_eco55192, w_eco55193, w_eco55194, w_eco55195, w_eco55196, w_eco55197, w_eco55198, w_eco55199, w_eco55200, w_eco55201, w_eco55202, w_eco55203, w_eco55204, w_eco55205, w_eco55206, w_eco55207, w_eco55208, w_eco55209, w_eco55210, w_eco55211, w_eco55212, w_eco55213, w_eco55214, w_eco55215, w_eco55216, w_eco55217, w_eco55218, w_eco55219, w_eco55220, w_eco55221, w_eco55222, w_eco55223, w_eco55224, w_eco55225, w_eco55226, w_eco55227, w_eco55228, w_eco55229, w_eco55230, w_eco55231, w_eco55232, w_eco55233, w_eco55234, w_eco55235, w_eco55236, w_eco55237, w_eco55238, w_eco55239, w_eco55240, w_eco55241, w_eco55242, w_eco55243, w_eco55244, w_eco55245, w_eco55246, w_eco55247, w_eco55248, w_eco55249, w_eco55250, w_eco55251, w_eco55252, w_eco55253, w_eco55254, w_eco55255, w_eco55256, w_eco55257, w_eco55258, w_eco55259, w_eco55260, w_eco55261, w_eco55262, w_eco55263, w_eco55264, w_eco55265, w_eco55266, w_eco55267, w_eco55268, w_eco55269, w_eco55270, w_eco55271, w_eco55272, w_eco55273, w_eco55274, w_eco55275, w_eco55276, w_eco55277, w_eco55278, w_eco55279, w_eco55280, w_eco55281, w_eco55282, w_eco55283, w_eco55284, w_eco55285, w_eco55286, w_eco55287, w_eco55288, w_eco55289, w_eco55290, w_eco55291, w_eco55292, w_eco55293, w_eco55294, w_eco55295, w_eco55296, w_eco55297, w_eco55298, w_eco55299, w_eco55300, w_eco55301, w_eco55302, w_eco55303, w_eco55304, w_eco55305, w_eco55306, w_eco55307, w_eco55308, w_eco55309, w_eco55310, w_eco55311, w_eco55312, w_eco55313, w_eco55314, w_eco55315, w_eco55316, w_eco55317, w_eco55318, w_eco55319, w_eco55320, w_eco55321, w_eco55322, w_eco55323, w_eco55324, w_eco55325, w_eco55326, w_eco55327, w_eco55328, w_eco55329, w_eco55330, w_eco55331, w_eco55332, w_eco55333, w_eco55334, w_eco55335, w_eco55336, w_eco55337, w_eco55338, w_eco55339, w_eco55340, w_eco55341, w_eco55342, w_eco55343, w_eco55344, w_eco55345, w_eco55346, w_eco55347, w_eco55348, w_eco55349, w_eco55350, w_eco55351, w_eco55352, w_eco55353, w_eco55354, w_eco55355, w_eco55356, w_eco55357, w_eco55358, w_eco55359, w_eco55360, w_eco55361, w_eco55362, w_eco55363, w_eco55364, w_eco55365, w_eco55366, w_eco55367, w_eco55368, w_eco55369, w_eco55370, w_eco55371, w_eco55372, w_eco55373, w_eco55374, w_eco55375, w_eco55376, w_eco55377, w_eco55378, w_eco55379, w_eco55380, w_eco55381, w_eco55382, w_eco55383, w_eco55384, w_eco55385, w_eco55386, w_eco55387, w_eco55388, w_eco55389, w_eco55390, w_eco55391, w_eco55392, w_eco55393, w_eco55394, w_eco55395, w_eco55396, w_eco55397, w_eco55398, w_eco55399, w_eco55400, w_eco55401, w_eco55402, w_eco55403, w_eco55404, w_eco55405, w_eco55406, w_eco55407, w_eco55408, w_eco55409, w_eco55410, w_eco55411, w_eco55412, w_eco55413, w_eco55414, w_eco55415, w_eco55416, w_eco55417, w_eco55418, w_eco55419, w_eco55420, w_eco55421, w_eco55422, w_eco55423, w_eco55424, w_eco55425, w_eco55426, w_eco55427, w_eco55428, w_eco55429, w_eco55430, w_eco55431, w_eco55432, w_eco55433, w_eco55434, w_eco55435, w_eco55436, w_eco55437, w_eco55438, w_eco55439, w_eco55440, w_eco55441, w_eco55442, w_eco55443, w_eco55444, w_eco55445, w_eco55446, w_eco55447, w_eco55448, w_eco55449, w_eco55450, w_eco55451, w_eco55452, w_eco55453, w_eco55454, w_eco55455, w_eco55456, w_eco55457, w_eco55458, w_eco55459, w_eco55460, w_eco55461, w_eco55462, w_eco55463, w_eco55464, w_eco55465, w_eco55466, w_eco55467, w_eco55468, w_eco55469, w_eco55470, w_eco55471, w_eco55472, w_eco55473, w_eco55474, w_eco55475, w_eco55476, w_eco55477, w_eco55478, w_eco55479, w_eco55480, w_eco55481, w_eco55482, w_eco55483, w_eco55484, w_eco55485, w_eco55486, w_eco55487, w_eco55488, w_eco55489, w_eco55490, w_eco55491, w_eco55492, w_eco55493, w_eco55494, w_eco55495, w_eco55496, w_eco55497, w_eco55498, w_eco55499, w_eco55500, w_eco55501, w_eco55502, w_eco55503, w_eco55504, w_eco55505, w_eco55506, w_eco55507, w_eco55508, w_eco55509, w_eco55510, w_eco55511, w_eco55512, w_eco55513, w_eco55514, w_eco55515, w_eco55516, w_eco55517, w_eco55518, w_eco55519, w_eco55520, w_eco55521, w_eco55522, w_eco55523, w_eco55524, w_eco55525, w_eco55526, w_eco55527, w_eco55528, w_eco55529, w_eco55530, w_eco55531, w_eco55532, w_eco55533, w_eco55534, w_eco55535, w_eco55536, w_eco55537, w_eco55538, w_eco55539, w_eco55540, w_eco55541, w_eco55542, w_eco55543, w_eco55544, w_eco55545, w_eco55546, w_eco55547, w_eco55548, w_eco55549, w_eco55550, w_eco55551, w_eco55552, w_eco55553, w_eco55554, w_eco55555, w_eco55556, w_eco55557, w_eco55558, w_eco55559, w_eco55560, w_eco55561, w_eco55562, w_eco55563, w_eco55564, w_eco55565, w_eco55566, w_eco55567, w_eco55568, w_eco55569, w_eco55570, w_eco55571, w_eco55572, w_eco55573, w_eco55574, w_eco55575, w_eco55576, w_eco55577, w_eco55578, w_eco55579, w_eco55580, w_eco55581, w_eco55582, w_eco55583, w_eco55584, w_eco55585, w_eco55586, w_eco55587, w_eco55588, w_eco55589, w_eco55590, w_eco55591, w_eco55592, w_eco55593, w_eco55594, w_eco55595, w_eco55596, w_eco55597, w_eco55598, w_eco55599, w_eco55600, w_eco55601, w_eco55602, w_eco55603, w_eco55604, w_eco55605, w_eco55606, w_eco55607, w_eco55608, w_eco55609, w_eco55610, w_eco55611, w_eco55612, w_eco55613, w_eco55614, w_eco55615, w_eco55616, w_eco55617, w_eco55618, w_eco55619, w_eco55620, w_eco55621, w_eco55622, w_eco55623, w_eco55624, w_eco55625, w_eco55626, w_eco55627, w_eco55628, w_eco55629, w_eco55630, w_eco55631, w_eco55632, w_eco55633, w_eco55634, w_eco55635, w_eco55636, w_eco55637, w_eco55638, w_eco55639, w_eco55640, w_eco55641, w_eco55642, w_eco55643, w_eco55644, w_eco55645, w_eco55646, w_eco55647, w_eco55648, w_eco55649, w_eco55650, w_eco55651, w_eco55652, w_eco55653, w_eco55654, w_eco55655, w_eco55656, w_eco55657, w_eco55658, w_eco55659, w_eco55660, w_eco55661, w_eco55662, w_eco55663, w_eco55664, w_eco55665, w_eco55666, w_eco55667, w_eco55668, w_eco55669, w_eco55670, w_eco55671, w_eco55672, w_eco55673, w_eco55674, w_eco55675, w_eco55676, w_eco55677, w_eco55678, w_eco55679, w_eco55680, w_eco55681, w_eco55682, w_eco55683, w_eco55684, w_eco55685, w_eco55686, w_eco55687, w_eco55688, w_eco55689, w_eco55690, w_eco55691, w_eco55692, w_eco55693, w_eco55694, w_eco55695, w_eco55696, w_eco55697, w_eco55698, w_eco55699, w_eco55700, w_eco55701, w_eco55702, w_eco55703, w_eco55704, w_eco55705, w_eco55706, w_eco55707, w_eco55708, w_eco55709, w_eco55710, w_eco55711, w_eco55712, w_eco55713, w_eco55714, w_eco55715, w_eco55716, w_eco55717, w_eco55718, w_eco55719, w_eco55720, w_eco55721, w_eco55722, w_eco55723, w_eco55724, w_eco55725, w_eco55726, w_eco55727, w_eco55728, w_eco55729, w_eco55730, w_eco55731, w_eco55732, w_eco55733, w_eco55734, w_eco55735, w_eco55736, w_eco55737, w_eco55738, w_eco55739, w_eco55740, w_eco55741, w_eco55742, w_eco55743, w_eco55744, w_eco55745, w_eco55746, w_eco55747, w_eco55748, w_eco55749, w_eco55750, w_eco55751, w_eco55752, w_eco55753, w_eco55754, w_eco55755, w_eco55756, w_eco55757, w_eco55758, w_eco55759, w_eco55760, w_eco55761, w_eco55762, w_eco55763, w_eco55764, w_eco55765, w_eco55766, w_eco55767, w_eco55768, w_eco55769, w_eco55770, w_eco55771, w_eco55772, w_eco55773, w_eco55774, w_eco55775, w_eco55776, w_eco55777, w_eco55778, w_eco55779, w_eco55780, w_eco55781, w_eco55782, w_eco55783, w_eco55784, w_eco55785, w_eco55786, w_eco55787, w_eco55788, w_eco55789, w_eco55790, w_eco55791, w_eco55792, w_eco55793, w_eco55794, w_eco55795, w_eco55796, w_eco55797, w_eco55798, w_eco55799, w_eco55800, w_eco55801, w_eco55802, w_eco55803, w_eco55804, w_eco55805, w_eco55806, w_eco55807, w_eco55808, w_eco55809, w_eco55810, w_eco55811, w_eco55812, w_eco55813, w_eco55814, w_eco55815, w_eco55816, w_eco55817, w_eco55818, w_eco55819, w_eco55820, w_eco55821, w_eco55822, w_eco55823, w_eco55824, w_eco55825, w_eco55826, w_eco55827, w_eco55828, w_eco55829, w_eco55830, w_eco55831, w_eco55832, w_eco55833, w_eco55834, w_eco55835, w_eco55836, w_eco55837, w_eco55838, w_eco55839, w_eco55840, w_eco55841, w_eco55842, w_eco55843, w_eco55844, w_eco55845, w_eco55846, w_eco55847, w_eco55848, w_eco55849, w_eco55850, w_eco55851, w_eco55852, w_eco55853, w_eco55854, w_eco55855, w_eco55856, w_eco55857, w_eco55858, w_eco55859, w_eco55860, w_eco55861, w_eco55862, w_eco55863, w_eco55864, w_eco55865, w_eco55866, w_eco55867, w_eco55868, w_eco55869, w_eco55870, w_eco55871, w_eco55872, w_eco55873, w_eco55874, w_eco55875, w_eco55876, w_eco55877, w_eco55878, w_eco55879, w_eco55880, w_eco55881, w_eco55882, w_eco55883, w_eco55884, w_eco55885, w_eco55886, w_eco55887, w_eco55888, w_eco55889, w_eco55890, w_eco55891, w_eco55892, w_eco55893, w_eco55894, w_eco55895, w_eco55896, w_eco55897, w_eco55898, w_eco55899, w_eco55900, w_eco55901, w_eco55902, w_eco55903, w_eco55904, w_eco55905, w_eco55906, w_eco55907, w_eco55908, w_eco55909, w_eco55910, w_eco55911, w_eco55912, w_eco55913, w_eco55914, w_eco55915, w_eco55916, w_eco55917, w_eco55918, w_eco55919, w_eco55920, w_eco55921, w_eco55922, w_eco55923, w_eco55924, w_eco55925, w_eco55926, w_eco55927, w_eco55928, w_eco55929, w_eco55930, w_eco55931, w_eco55932, w_eco55933, w_eco55934, w_eco55935, w_eco55936, w_eco55937, w_eco55938, w_eco55939, w_eco55940, w_eco55941, w_eco55942, w_eco55943, w_eco55944, w_eco55945, w_eco55946, w_eco55947, w_eco55948, w_eco55949, w_eco55950, w_eco55951, w_eco55952, w_eco55953, w_eco55954, w_eco55955, w_eco55956, w_eco55957, w_eco55958, w_eco55959, w_eco55960, w_eco55961, w_eco55962, w_eco55963, w_eco55964, w_eco55965, w_eco55966, w_eco55967, w_eco55968, w_eco55969, w_eco55970, w_eco55971, w_eco55972, w_eco55973, w_eco55974, w_eco55975, w_eco55976, w_eco55977, w_eco55978, w_eco55979, w_eco55980, w_eco55981, w_eco55982, w_eco55983, w_eco55984, w_eco55985, w_eco55986, w_eco55987, w_eco55988, w_eco55989, w_eco55990, w_eco55991, w_eco55992, w_eco55993, w_eco55994, w_eco55995, w_eco55996, w_eco55997, w_eco55998, w_eco55999, w_eco56000, w_eco56001, w_eco56002, w_eco56003, w_eco56004, w_eco56005, w_eco56006, w_eco56007, w_eco56008, w_eco56009, w_eco56010, w_eco56011, w_eco56012, w_eco56013, w_eco56014, w_eco56015, w_eco56016, w_eco56017, w_eco56018, w_eco56019, w_eco56020, w_eco56021, w_eco56022, w_eco56023, w_eco56024, w_eco56025, w_eco56026, w_eco56027, w_eco56028, w_eco56029, w_eco56030, w_eco56031, w_eco56032, w_eco56033, w_eco56034, w_eco56035, w_eco56036, w_eco56037, w_eco56038, w_eco56039, w_eco56040, w_eco56041, w_eco56042, w_eco56043, w_eco56044, w_eco56045, w_eco56046, w_eco56047, w_eco56048, w_eco56049, w_eco56050, w_eco56051, w_eco56052, w_eco56053, w_eco56054, w_eco56055, w_eco56056, w_eco56057, w_eco56058, w_eco56059, w_eco56060, w_eco56061, w_eco56062, w_eco56063, w_eco56064, w_eco56065, w_eco56066, w_eco56067, w_eco56068, w_eco56069, w_eco56070, w_eco56071, w_eco56072, w_eco56073, w_eco56074, w_eco56075, w_eco56076, w_eco56077, w_eco56078, w_eco56079, w_eco56080, w_eco56081, w_eco56082, w_eco56083, w_eco56084, w_eco56085, w_eco56086, w_eco56087, w_eco56088, w_eco56089, w_eco56090, w_eco56091, w_eco56092, w_eco56093, w_eco56094, w_eco56095, w_eco56096, w_eco56097, w_eco56098, w_eco56099, w_eco56100, w_eco56101, w_eco56102, w_eco56103, w_eco56104, w_eco56105, w_eco56106, w_eco56107, w_eco56108, w_eco56109, w_eco56110, w_eco56111, w_eco56112, w_eco56113, w_eco56114, w_eco56115, w_eco56116, w_eco56117, w_eco56118, w_eco56119, w_eco56120, w_eco56121, w_eco56122, w_eco56123, w_eco56124, w_eco56125, w_eco56126, w_eco56127, w_eco56128, w_eco56129, w_eco56130, w_eco56131, w_eco56132, w_eco56133, w_eco56134, w_eco56135, w_eco56136, w_eco56137, w_eco56138, w_eco56139, w_eco56140, w_eco56141, w_eco56142, w_eco56143, w_eco56144, w_eco56145, w_eco56146, w_eco56147, w_eco56148, w_eco56149, w_eco56150, w_eco56151, w_eco56152, w_eco56153, w_eco56154, w_eco56155, w_eco56156, w_eco56157, w_eco56158, w_eco56159, w_eco56160, w_eco56161, w_eco56162, w_eco56163, w_eco56164, w_eco56165, w_eco56166, w_eco56167, w_eco56168, w_eco56169, w_eco56170, w_eco56171, w_eco56172, w_eco56173, w_eco56174, w_eco56175, w_eco56176, w_eco56177, w_eco56178, w_eco56179, w_eco56180, w_eco56181, w_eco56182, w_eco56183, w_eco56184, w_eco56185, w_eco56186, w_eco56187, w_eco56188, w_eco56189, w_eco56190, w_eco56191, w_eco56192, w_eco56193, w_eco56194, w_eco56195, w_eco56196, w_eco56197, w_eco56198, w_eco56199, w_eco56200, w_eco56201, w_eco56202, w_eco56203, w_eco56204, w_eco56205, w_eco56206, w_eco56207, w_eco56208, w_eco56209, w_eco56210, w_eco56211, w_eco56212, w_eco56213, w_eco56214, w_eco56215, w_eco56216, w_eco56217, w_eco56218, w_eco56219, w_eco56220, w_eco56221, w_eco56222, w_eco56223, w_eco56224, w_eco56225, w_eco56226, w_eco56227, w_eco56228, w_eco56229, w_eco56230, w_eco56231, w_eco56232, w_eco56233, w_eco56234, w_eco56235, w_eco56236, w_eco56237, w_eco56238, w_eco56239, w_eco56240, w_eco56241, w_eco56242, w_eco56243, w_eco56244, w_eco56245, w_eco56246, w_eco56247, w_eco56248, w_eco56249, w_eco56250, w_eco56251, w_eco56252, w_eco56253, w_eco56254, w_eco56255, w_eco56256, w_eco56257, w_eco56258, w_eco56259, w_eco56260, w_eco56261, w_eco56262, w_eco56263, w_eco56264, w_eco56265, w_eco56266, w_eco56267, w_eco56268, w_eco56269, w_eco56270, w_eco56271, w_eco56272, w_eco56273, w_eco56274, w_eco56275, w_eco56276, w_eco56277, w_eco56278, w_eco56279, w_eco56280, w_eco56281, w_eco56282, w_eco56283, w_eco56284, w_eco56285, w_eco56286, w_eco56287, w_eco56288, w_eco56289, w_eco56290, w_eco56291, w_eco56292, w_eco56293, w_eco56294, w_eco56295, w_eco56296, w_eco56297, w_eco56298, w_eco56299, w_eco56300, w_eco56301, w_eco56302, w_eco56303, w_eco56304, w_eco56305, w_eco56306, w_eco56307, w_eco56308, w_eco56309, w_eco56310, w_eco56311, w_eco56312, w_eco56313, w_eco56314, w_eco56315, w_eco56316, w_eco56317, w_eco56318, w_eco56319, w_eco56320, w_eco56321, w_eco56322, w_eco56323, w_eco56324, w_eco56325, w_eco56326, w_eco56327, w_eco56328, w_eco56329, w_eco56330, w_eco56331, w_eco56332, w_eco56333, w_eco56334, w_eco56335, w_eco56336, w_eco56337, w_eco56338, w_eco56339, w_eco56340, w_eco56341, w_eco56342, w_eco56343, w_eco56344, w_eco56345, w_eco56346, w_eco56347, w_eco56348, w_eco56349, w_eco56350, w_eco56351, w_eco56352, w_eco56353, w_eco56354, w_eco56355, w_eco56356, w_eco56357, w_eco56358, w_eco56359, w_eco56360, w_eco56361, w_eco56362, w_eco56363, w_eco56364, w_eco56365, w_eco56366, w_eco56367, w_eco56368, w_eco56369, w_eco56370, w_eco56371, w_eco56372, w_eco56373, w_eco56374, w_eco56375, w_eco56376, w_eco56377, w_eco56378, w_eco56379, w_eco56380, w_eco56381, w_eco56382, w_eco56383, w_eco56384, w_eco56385, w_eco56386, w_eco56387, w_eco56388, w_eco56389, w_eco56390, w_eco56391, w_eco56392, w_eco56393, w_eco56394, w_eco56395, w_eco56396, w_eco56397, w_eco56398, w_eco56399, w_eco56400, w_eco56401, w_eco56402, w_eco56403, w_eco56404, w_eco56405, w_eco56406, w_eco56407, w_eco56408, w_eco56409, w_eco56410, w_eco56411, w_eco56412, w_eco56413, w_eco56414, w_eco56415, w_eco56416, w_eco56417, w_eco56418, w_eco56419, w_eco56420, w_eco56421, w_eco56422, w_eco56423, w_eco56424, w_eco56425, w_eco56426, w_eco56427, w_eco56428, w_eco56429, w_eco56430, w_eco56431, w_eco56432, w_eco56433, w_eco56434, w_eco56435, w_eco56436, w_eco56437, w_eco56438, w_eco56439, w_eco56440, w_eco56441, w_eco56442, w_eco56443, w_eco56444, w_eco56445, w_eco56446, w_eco56447, w_eco56448, w_eco56449, w_eco56450, w_eco56451, w_eco56452, w_eco56453, w_eco56454, w_eco56455, w_eco56456, w_eco56457, w_eco56458, w_eco56459, w_eco56460, w_eco56461, w_eco56462, w_eco56463, w_eco56464, w_eco56465, w_eco56466, w_eco56467, w_eco56468, w_eco56469, w_eco56470, w_eco56471, w_eco56472, w_eco56473, w_eco56474, w_eco56475, w_eco56476, w_eco56477, w_eco56478, w_eco56479, w_eco56480, w_eco56481, w_eco56482, w_eco56483, w_eco56484, w_eco56485, w_eco56486, w_eco56487, w_eco56488, w_eco56489, w_eco56490, w_eco56491, w_eco56492, w_eco56493, w_eco56494, w_eco56495, w_eco56496, w_eco56497, w_eco56498, w_eco56499, w_eco56500, w_eco56501, w_eco56502, w_eco56503, w_eco56504, w_eco56505, w_eco56506, w_eco56507, w_eco56508, w_eco56509, w_eco56510, w_eco56511, w_eco56512, w_eco56513, w_eco56514, w_eco56515, w_eco56516, w_eco56517, w_eco56518, w_eco56519, w_eco56520, w_eco56521, w_eco56522, w_eco56523, w_eco56524, w_eco56525, w_eco56526, w_eco56527, w_eco56528, w_eco56529, w_eco56530, w_eco56531, w_eco56532, w_eco56533, w_eco56534, w_eco56535, w_eco56536, w_eco56537, w_eco56538, w_eco56539, w_eco56540, w_eco56541, w_eco56542, w_eco56543, w_eco56544, w_eco56545, w_eco56546, w_eco56547, w_eco56548, w_eco56549, w_eco56550, w_eco56551, w_eco56552, w_eco56553, w_eco56554, w_eco56555, w_eco56556, w_eco56557, w_eco56558, w_eco56559, w_eco56560, w_eco56561, w_eco56562, w_eco56563, w_eco56564, w_eco56565, w_eco56566, w_eco56567, w_eco56568, w_eco56569, w_eco56570, w_eco56571, w_eco56572, w_eco56573, w_eco56574, w_eco56575, w_eco56576, w_eco56577, w_eco56578, w_eco56579, w_eco56580, w_eco56581, w_eco56582, w_eco56583, w_eco56584, w_eco56585, w_eco56586, w_eco56587, w_eco56588, w_eco56589, w_eco56590, w_eco56591, w_eco56592, w_eco56593, w_eco56594, w_eco56595, w_eco56596, w_eco56597, w_eco56598, w_eco56599, w_eco56600, w_eco56601, w_eco56602, w_eco56603, w_eco56604, w_eco56605, w_eco56606, w_eco56607, w_eco56608, w_eco56609, w_eco56610, w_eco56611, w_eco56612, w_eco56613, w_eco56614, w_eco56615, w_eco56616, w_eco56617, w_eco56618, w_eco56619, w_eco56620, w_eco56621, w_eco56622, w_eco56623, w_eco56624, w_eco56625, w_eco56626, w_eco56627, w_eco56628, w_eco56629, w_eco56630, w_eco56631, w_eco56632, w_eco56633, w_eco56634, w_eco56635, w_eco56636, w_eco56637, w_eco56638, w_eco56639, w_eco56640, w_eco56641, w_eco56642, w_eco56643, w_eco56644, w_eco56645, w_eco56646, w_eco56647, w_eco56648, w_eco56649, w_eco56650, w_eco56651, w_eco56652, w_eco56653, w_eco56654, w_eco56655, w_eco56656, w_eco56657, w_eco56658, w_eco56659, w_eco56660, w_eco56661, w_eco56662, w_eco56663, w_eco56664, w_eco56665, w_eco56666, w_eco56667, w_eco56668, w_eco56669, w_eco56670, w_eco56671, w_eco56672, w_eco56673, w_eco56674, w_eco56675, w_eco56676, w_eco56677, w_eco56678, w_eco56679, w_eco56680, w_eco56681, w_eco56682, w_eco56683, w_eco56684, w_eco56685, w_eco56686, w_eco56687, w_eco56688, w_eco56689, w_eco56690, w_eco56691, w_eco56692, w_eco56693, w_eco56694, w_eco56695, w_eco56696, w_eco56697, w_eco56698, w_eco56699, w_eco56700, w_eco56701, w_eco56702, w_eco56703, w_eco56704, w_eco56705, w_eco56706, w_eco56707, w_eco56708, w_eco56709, w_eco56710, w_eco56711, w_eco56712, w_eco56713, w_eco56714, w_eco56715, w_eco56716, w_eco56717, w_eco56718, w_eco56719, w_eco56720, w_eco56721, w_eco56722, w_eco56723, w_eco56724, w_eco56725, w_eco56726, w_eco56727, w_eco56728, w_eco56729, w_eco56730, w_eco56731, w_eco56732, w_eco56733, w_eco56734, w_eco56735, w_eco56736, w_eco56737, w_eco56738, w_eco56739, w_eco56740, w_eco56741, w_eco56742, w_eco56743, w_eco56744, w_eco56745, w_eco56746, w_eco56747, w_eco56748, w_eco56749, w_eco56750, w_eco56751, w_eco56752, w_eco56753, w_eco56754, w_eco56755, w_eco56756, w_eco56757, w_eco56758, w_eco56759, w_eco56760, w_eco56761, w_eco56762, w_eco56763, w_eco56764, w_eco56765, w_eco56766, w_eco56767, w_eco56768, w_eco56769, w_eco56770, w_eco56771, w_eco56772, w_eco56773, w_eco56774, w_eco56775, w_eco56776, w_eco56777, w_eco56778, w_eco56779, w_eco56780, w_eco56781, w_eco56782, w_eco56783, w_eco56784, w_eco56785, w_eco56786, w_eco56787, w_eco56788, w_eco56789, w_eco56790, w_eco56791, w_eco56792, w_eco56793, w_eco56794, w_eco56795, w_eco56796, w_eco56797, w_eco56798, w_eco56799, w_eco56800, w_eco56801, w_eco56802, w_eco56803, w_eco56804, w_eco56805, w_eco56806, w_eco56807, w_eco56808, w_eco56809, w_eco56810, w_eco56811, w_eco56812, w_eco56813, w_eco56814, w_eco56815, w_eco56816, w_eco56817, w_eco56818, w_eco56819, w_eco56820, w_eco56821, w_eco56822, w_eco56823, w_eco56824, w_eco56825, w_eco56826, w_eco56827, w_eco56828, w_eco56829, w_eco56830, w_eco56831, w_eco56832, w_eco56833, w_eco56834, w_eco56835, w_eco56836, w_eco56837, w_eco56838, w_eco56839, w_eco56840, w_eco56841, w_eco56842, w_eco56843, w_eco56844, w_eco56845, w_eco56846, w_eco56847, w_eco56848, w_eco56849, w_eco56850, w_eco56851, w_eco56852, w_eco56853, w_eco56854, w_eco56855, w_eco56856, w_eco56857, w_eco56858, w_eco56859, w_eco56860, w_eco56861, w_eco56862, w_eco56863, w_eco56864, w_eco56865, w_eco56866, w_eco56867, w_eco56868, w_eco56869, w_eco56870, w_eco56871, w_eco56872, w_eco56873, w_eco56874, w_eco56875, w_eco56876, w_eco56877, w_eco56878, w_eco56879, w_eco56880, w_eco56881, w_eco56882, w_eco56883, w_eco56884, w_eco56885, w_eco56886, w_eco56887, w_eco56888, w_eco56889, w_eco56890, w_eco56891, w_eco56892, w_eco56893, w_eco56894, w_eco56895, w_eco56896, w_eco56897, w_eco56898, w_eco56899, w_eco56900, w_eco56901, w_eco56902, w_eco56903, w_eco56904, w_eco56905, w_eco56906, w_eco56907, w_eco56908, w_eco56909, w_eco56910, w_eco56911, w_eco56912, w_eco56913, w_eco56914, w_eco56915, w_eco56916, w_eco56917, w_eco56918, w_eco56919, w_eco56920, w_eco56921, w_eco56922, w_eco56923, w_eco56924, w_eco56925, w_eco56926, w_eco56927, w_eco56928, w_eco56929, w_eco56930, w_eco56931, w_eco56932, w_eco56933, w_eco56934, w_eco56935, w_eco56936, w_eco56937, w_eco56938, w_eco56939, w_eco56940, w_eco56941, w_eco56942, w_eco56943, w_eco56944, w_eco56945, w_eco56946, w_eco56947, w_eco56948, w_eco56949, w_eco56950, w_eco56951, w_eco56952, w_eco56953, w_eco56954, w_eco56955, w_eco56956, w_eco56957, w_eco56958, w_eco56959, w_eco56960, w_eco56961, w_eco56962, w_eco56963, w_eco56964, w_eco56965, w_eco56966, w_eco56967, w_eco56968, w_eco56969, w_eco56970, w_eco56971, w_eco56972, w_eco56973, w_eco56974, w_eco56975, w_eco56976, w_eco56977, w_eco56978, w_eco56979, w_eco56980, w_eco56981, w_eco56982, w_eco56983, w_eco56984, w_eco56985, w_eco56986, w_eco56987, w_eco56988, w_eco56989, w_eco56990, w_eco56991, w_eco56992, w_eco56993, w_eco56994, w_eco56995, w_eco56996, w_eco56997, w_eco56998, w_eco56999, w_eco57000, w_eco57001, w_eco57002, w_eco57003, w_eco57004, w_eco57005, w_eco57006, w_eco57007, w_eco57008, w_eco57009, w_eco57010, w_eco57011, w_eco57012, w_eco57013, w_eco57014, w_eco57015, w_eco57016, w_eco57017, w_eco57018, w_eco57019, w_eco57020, w_eco57021, w_eco57022, w_eco57023, w_eco57024, w_eco57025, w_eco57026, w_eco57027, w_eco57028, w_eco57029, w_eco57030, w_eco57031, w_eco57032, w_eco57033, w_eco57034, w_eco57035, w_eco57036, w_eco57037, w_eco57038, w_eco57039, w_eco57040, w_eco57041, w_eco57042, w_eco57043, w_eco57044, w_eco57045, w_eco57046, w_eco57047, w_eco57048, w_eco57049, w_eco57050, w_eco57051, w_eco57052, w_eco57053, w_eco57054, w_eco57055, w_eco57056, w_eco57057, w_eco57058, w_eco57059, w_eco57060, w_eco57061, w_eco57062, w_eco57063, w_eco57064, w_eco57065, w_eco57066, w_eco57067, w_eco57068, w_eco57069, w_eco57070, w_eco57071, w_eco57072, w_eco57073, w_eco57074, w_eco57075, w_eco57076, w_eco57077, w_eco57078, w_eco57079, w_eco57080, w_eco57081, w_eco57082, w_eco57083, w_eco57084, w_eco57085, w_eco57086, w_eco57087, w_eco57088, w_eco57089, w_eco57090, w_eco57091, w_eco57092, w_eco57093, w_eco57094, w_eco57095, w_eco57096, w_eco57097, w_eco57098, w_eco57099, w_eco57100, w_eco57101, w_eco57102, w_eco57103, w_eco57104, w_eco57105, w_eco57106, w_eco57107, w_eco57108, w_eco57109, w_eco57110, w_eco57111, w_eco57112, w_eco57113, w_eco57114, w_eco57115, w_eco57116, w_eco57117, w_eco57118, w_eco57119, w_eco57120, w_eco57121, w_eco57122, w_eco57123, w_eco57124, w_eco57125, w_eco57126, w_eco57127, w_eco57128, w_eco57129, w_eco57130, w_eco57131, w_eco57132, w_eco57133, w_eco57134, w_eco57135, w_eco57136, w_eco57137, w_eco57138, w_eco57139, w_eco57140, w_eco57141, w_eco57142, w_eco57143, w_eco57144, w_eco57145, w_eco57146, w_eco57147, w_eco57148, w_eco57149, w_eco57150, w_eco57151, w_eco57152, w_eco57153, w_eco57154, w_eco57155, w_eco57156, w_eco57157, w_eco57158, w_eco57159, w_eco57160, w_eco57161, w_eco57162, w_eco57163, w_eco57164, w_eco57165, w_eco57166, w_eco57167, w_eco57168, w_eco57169, w_eco57170, w_eco57171, w_eco57172, w_eco57173, w_eco57174, w_eco57175, w_eco57176, w_eco57177, w_eco57178, w_eco57179, w_eco57180, w_eco57181, w_eco57182, w_eco57183, w_eco57184, w_eco57185, w_eco57186, w_eco57187, w_eco57188, w_eco57189, w_eco57190, w_eco57191, w_eco57192, w_eco57193, w_eco57194, w_eco57195, w_eco57196, w_eco57197, w_eco57198, w_eco57199, w_eco57200, w_eco57201, w_eco57202, w_eco57203, w_eco57204, w_eco57205, w_eco57206, w_eco57207, w_eco57208, w_eco57209, w_eco57210, w_eco57211, w_eco57212, w_eco57213, w_eco57214, w_eco57215, w_eco57216, w_eco57217, w_eco57218, w_eco57219, w_eco57220, w_eco57221, w_eco57222, w_eco57223, w_eco57224, w_eco57225, w_eco57226, w_eco57227, w_eco57228, w_eco57229, w_eco57230, w_eco57231, w_eco57232, w_eco57233, w_eco57234, w_eco57235, w_eco57236, w_eco57237, w_eco57238, w_eco57239, w_eco57240, w_eco57241, w_eco57242, w_eco57243, w_eco57244, w_eco57245, w_eco57246, w_eco57247, w_eco57248, w_eco57249, w_eco57250, w_eco57251, w_eco57252, w_eco57253, w_eco57254, w_eco57255, w_eco57256, w_eco57257, w_eco57258, w_eco57259, w_eco57260, w_eco57261, w_eco57262, w_eco57263, w_eco57264, w_eco57265, w_eco57266, w_eco57267, w_eco57268, w_eco57269, w_eco57270, w_eco57271, w_eco57272, w_eco57273, w_eco57274, w_eco57275, w_eco57276, w_eco57277, w_eco57278, w_eco57279, w_eco57280, w_eco57281, w_eco57282, w_eco57283, w_eco57284, w_eco57285, w_eco57286, w_eco57287, w_eco57288, w_eco57289, w_eco57290, w_eco57291, w_eco57292, w_eco57293, w_eco57294, w_eco57295, w_eco57296, w_eco57297, w_eco57298, w_eco57299, w_eco57300, w_eco57301, w_eco57302, w_eco57303, w_eco57304, w_eco57305, w_eco57306, w_eco57307, w_eco57308, w_eco57309, w_eco57310, w_eco57311, w_eco57312, w_eco57313, w_eco57314, w_eco57315, w_eco57316, w_eco57317, w_eco57318, w_eco57319, w_eco57320, w_eco57321, w_eco57322, w_eco57323, w_eco57324, w_eco57325, w_eco57326, w_eco57327, w_eco57328, w_eco57329, w_eco57330, w_eco57331, w_eco57332, w_eco57333, w_eco57334, w_eco57335, w_eco57336, w_eco57337, w_eco57338, w_eco57339, w_eco57340, w_eco57341, w_eco57342, w_eco57343, w_eco57344, w_eco57345, w_eco57346, w_eco57347, w_eco57348, w_eco57349, w_eco57350, w_eco57351, w_eco57352, w_eco57353, w_eco57354, w_eco57355, w_eco57356, w_eco57357, w_eco57358, w_eco57359, w_eco57360, w_eco57361, w_eco57362, w_eco57363, w_eco57364, w_eco57365, w_eco57366, w_eco57367, w_eco57368, w_eco57369, w_eco57370, w_eco57371, w_eco57372, w_eco57373, w_eco57374, w_eco57375, w_eco57376, w_eco57377, w_eco57378, w_eco57379, w_eco57380, w_eco57381, w_eco57382, w_eco57383, w_eco57384, w_eco57385, w_eco57386, w_eco57387, w_eco57388, w_eco57389, w_eco57390, w_eco57391, w_eco57392, w_eco57393, w_eco57394, w_eco57395, w_eco57396, w_eco57397, w_eco57398, w_eco57399, w_eco57400, w_eco57401, w_eco57402, w_eco57403, w_eco57404, w_eco57405, w_eco57406, w_eco57407, w_eco57408, w_eco57409, w_eco57410, w_eco57411, w_eco57412, w_eco57413, w_eco57414, w_eco57415, w_eco57416, w_eco57417, w_eco57418, w_eco57419, w_eco57420, w_eco57421, w_eco57422, w_eco57423, w_eco57424, w_eco57425, w_eco57426, w_eco57427, w_eco57428, w_eco57429, w_eco57430, w_eco57431, w_eco57432, w_eco57433, w_eco57434, w_eco57435, w_eco57436, w_eco57437, w_eco57438, w_eco57439, w_eco57440, w_eco57441, w_eco57442, w_eco57443, w_eco57444, w_eco57445, w_eco57446, w_eco57447, w_eco57448, w_eco57449, w_eco57450, w_eco57451, w_eco57452, w_eco57453, w_eco57454, w_eco57455, w_eco57456, w_eco57457, w_eco57458, w_eco57459, w_eco57460, w_eco57461, w_eco57462, w_eco57463, w_eco57464, w_eco57465, w_eco57466, w_eco57467, w_eco57468, w_eco57469, w_eco57470, w_eco57471, w_eco57472, w_eco57473, w_eco57474, w_eco57475, w_eco57476, w_eco57477, w_eco57478, w_eco57479, w_eco57480, w_eco57481, w_eco57482, w_eco57483, w_eco57484, w_eco57485, w_eco57486, w_eco57487, w_eco57488, w_eco57489, w_eco57490, w_eco57491, w_eco57492, w_eco57493, w_eco57494, w_eco57495, w_eco57496, w_eco57497, w_eco57498, w_eco57499, w_eco57500, w_eco57501, w_eco57502, w_eco57503, w_eco57504, w_eco57505, w_eco57506, w_eco57507, w_eco57508, w_eco57509, w_eco57510, w_eco57511, w_eco57512, w_eco57513, w_eco57514, w_eco57515, w_eco57516, w_eco57517, w_eco57518, w_eco57519, w_eco57520, w_eco57521, w_eco57522, w_eco57523, w_eco57524, w_eco57525, w_eco57526, w_eco57527, w_eco57528, w_eco57529, w_eco57530, w_eco57531, w_eco57532, w_eco57533, w_eco57534, w_eco57535, w_eco57536, w_eco57537, w_eco57538, w_eco57539, w_eco57540, w_eco57541, w_eco57542, w_eco57543, w_eco57544, w_eco57545, w_eco57546, w_eco57547, w_eco57548, w_eco57549, w_eco57550, w_eco57551, w_eco57552, w_eco57553, w_eco57554, w_eco57555, w_eco57556, w_eco57557, w_eco57558, w_eco57559, w_eco57560, w_eco57561, w_eco57562, w_eco57563, w_eco57564, w_eco57565, w_eco57566, w_eco57567, w_eco57568, w_eco57569, w_eco57570, w_eco57571, w_eco57572, w_eco57573, w_eco57574, w_eco57575, w_eco57576, w_eco57577, w_eco57578, w_eco57579, w_eco57580, w_eco57581, w_eco57582, w_eco57583, w_eco57584, w_eco57585, w_eco57586, w_eco57587, w_eco57588, w_eco57589, w_eco57590, w_eco57591, w_eco57592, w_eco57593, w_eco57594, w_eco57595, w_eco57596, w_eco57597, w_eco57598, w_eco57599, w_eco57600, w_eco57601, w_eco57602, w_eco57603, w_eco57604, w_eco57605, w_eco57606, w_eco57607, w_eco57608, w_eco57609, w_eco57610, w_eco57611, w_eco57612, w_eco57613, w_eco57614, w_eco57615, w_eco57616, w_eco57617, w_eco57618, w_eco57619, w_eco57620, w_eco57621, w_eco57622, w_eco57623, w_eco57624, w_eco57625, w_eco57626, w_eco57627, w_eco57628, w_eco57629, w_eco57630, w_eco57631, w_eco57632, w_eco57633, w_eco57634, w_eco57635, w_eco57636, w_eco57637, w_eco57638, w_eco57639, w_eco57640, w_eco57641, w_eco57642, w_eco57643, w_eco57644, w_eco57645, w_eco57646, w_eco57647, w_eco57648, w_eco57649, w_eco57650, w_eco57651, w_eco57652, w_eco57653, w_eco57654, w_eco57655, w_eco57656, w_eco57657, w_eco57658, w_eco57659, w_eco57660, w_eco57661, w_eco57662, w_eco57663, w_eco57664, w_eco57665, w_eco57666, w_eco57667, w_eco57668, w_eco57669, w_eco57670, w_eco57671, w_eco57672, w_eco57673, w_eco57674, w_eco57675, w_eco57676, w_eco57677, w_eco57678, w_eco57679, w_eco57680, w_eco57681, w_eco57682, w_eco57683, w_eco57684, w_eco57685, w_eco57686, w_eco57687, w_eco57688, w_eco57689, w_eco57690, w_eco57691, w_eco57692, w_eco57693, w_eco57694, w_eco57695, w_eco57696, w_eco57697, w_eco57698, w_eco57699, w_eco57700, w_eco57701, w_eco57702, w_eco57703, w_eco57704, w_eco57705, w_eco57706, w_eco57707, w_eco57708, w_eco57709, w_eco57710, w_eco57711, w_eco57712, w_eco57713, w_eco57714, w_eco57715, w_eco57716, w_eco57717, w_eco57718, w_eco57719, w_eco57720, w_eco57721, w_eco57722, w_eco57723, w_eco57724, w_eco57725, w_eco57726, w_eco57727, w_eco57728, w_eco57729, w_eco57730, w_eco57731, w_eco57732, w_eco57733, w_eco57734, w_eco57735, w_eco57736, w_eco57737, w_eco57738, w_eco57739, w_eco57740, w_eco57741, w_eco57742, w_eco57743, w_eco57744, w_eco57745, w_eco57746, w_eco57747, w_eco57748, w_eco57749, w_eco57750, w_eco57751, w_eco57752, w_eco57753, w_eco57754, w_eco57755, w_eco57756, w_eco57757, w_eco57758, w_eco57759, w_eco57760, w_eco57761, w_eco57762, w_eco57763, w_eco57764, w_eco57765, w_eco57766, w_eco57767, w_eco57768, w_eco57769, w_eco57770, w_eco57771, w_eco57772, w_eco57773, w_eco57774, w_eco57775, w_eco57776, w_eco57777, w_eco57778, w_eco57779, w_eco57780, w_eco57781, w_eco57782, w_eco57783, w_eco57784, w_eco57785, w_eco57786, w_eco57787, w_eco57788, w_eco57789, w_eco57790, w_eco57791, w_eco57792, w_eco57793, w_eco57794, w_eco57795, w_eco57796, w_eco57797, w_eco57798, w_eco57799, w_eco57800, w_eco57801, w_eco57802, w_eco57803, w_eco57804, w_eco57805, w_eco57806, w_eco57807, w_eco57808, w_eco57809, w_eco57810, w_eco57811, w_eco57812, w_eco57813, w_eco57814, w_eco57815, w_eco57816, w_eco57817, w_eco57818, w_eco57819, w_eco57820, w_eco57821, w_eco57822, w_eco57823, w_eco57824, w_eco57825, w_eco57826, w_eco57827, w_eco57828, w_eco57829, w_eco57830, w_eco57831, w_eco57832, w_eco57833, w_eco57834, w_eco57835, w_eco57836, w_eco57837, w_eco57838, w_eco57839, w_eco57840, w_eco57841, w_eco57842, w_eco57843, w_eco57844, w_eco57845, w_eco57846, w_eco57847, w_eco57848, w_eco57849, w_eco57850, w_eco57851, w_eco57852, w_eco57853, w_eco57854, w_eco57855, w_eco57856, w_eco57857, w_eco57858, w_eco57859, w_eco57860, w_eco57861, w_eco57862, w_eco57863, w_eco57864, w_eco57865, w_eco57866, w_eco57867, w_eco57868, w_eco57869, w_eco57870, w_eco57871, w_eco57872, w_eco57873, w_eco57874, w_eco57875, w_eco57876, w_eco57877, w_eco57878, w_eco57879, w_eco57880, w_eco57881, w_eco57882, w_eco57883, w_eco57884, w_eco57885, w_eco57886, w_eco57887, w_eco57888, w_eco57889, w_eco57890, w_eco57891, w_eco57892, w_eco57893, w_eco57894, w_eco57895, w_eco57896, w_eco57897, w_eco57898, w_eco57899, w_eco57900, w_eco57901, w_eco57902, w_eco57903, w_eco57904, w_eco57905, w_eco57906, w_eco57907, w_eco57908, w_eco57909, w_eco57910, w_eco57911, w_eco57912, w_eco57913, w_eco57914, w_eco57915, w_eco57916, w_eco57917, w_eco57918, w_eco57919, w_eco57920, w_eco57921, w_eco57922, w_eco57923, w_eco57924, w_eco57925, w_eco57926, w_eco57927, w_eco57928, w_eco57929, w_eco57930, w_eco57931, w_eco57932, w_eco57933, w_eco57934, w_eco57935, w_eco57936, w_eco57937, w_eco57938, w_eco57939, w_eco57940, w_eco57941, w_eco57942, w_eco57943, w_eco57944, w_eco57945, w_eco57946, w_eco57947, w_eco57948, w_eco57949, w_eco57950, w_eco57951, w_eco57952, w_eco57953, w_eco57954, w_eco57955, w_eco57956, w_eco57957, w_eco57958, w_eco57959, w_eco57960, w_eco57961, w_eco57962, w_eco57963, w_eco57964, w_eco57965, w_eco57966, w_eco57967, w_eco57968, w_eco57969, w_eco57970, w_eco57971, w_eco57972, w_eco57973, w_eco57974, w_eco57975, w_eco57976, w_eco57977, w_eco57978, w_eco57979, w_eco57980, w_eco57981, w_eco57982, w_eco57983, w_eco57984, w_eco57985, w_eco57986, w_eco57987, w_eco57988, w_eco57989, w_eco57990, w_eco57991, w_eco57992, w_eco57993, w_eco57994, w_eco57995, w_eco57996, w_eco57997, w_eco57998, w_eco57999, w_eco58000, w_eco58001, w_eco58002, w_eco58003, w_eco58004, w_eco58005, w_eco58006, w_eco58007, w_eco58008, w_eco58009, w_eco58010, w_eco58011, w_eco58012, w_eco58013, w_eco58014, w_eco58015, w_eco58016, w_eco58017, w_eco58018, w_eco58019, w_eco58020, w_eco58021, w_eco58022, w_eco58023, w_eco58024, w_eco58025, w_eco58026, w_eco58027, w_eco58028, w_eco58029, w_eco58030, w_eco58031, w_eco58032, w_eco58033, w_eco58034, w_eco58035, w_eco58036, w_eco58037, w_eco58038, w_eco58039, w_eco58040, w_eco58041, w_eco58042, w_eco58043, w_eco58044, w_eco58045, w_eco58046, w_eco58047, w_eco58048, w_eco58049, w_eco58050, w_eco58051, w_eco58052, w_eco58053, w_eco58054, w_eco58055, w_eco58056, w_eco58057, w_eco58058, w_eco58059, w_eco58060, w_eco58061, w_eco58062, w_eco58063, w_eco58064, w_eco58065, w_eco58066, w_eco58067, w_eco58068, w_eco58069, w_eco58070, w_eco58071, w_eco58072, w_eco58073, w_eco58074, w_eco58075, w_eco58076, w_eco58077, w_eco58078, w_eco58079, w_eco58080, w_eco58081, w_eco58082, w_eco58083, w_eco58084, w_eco58085, w_eco58086, w_eco58087, w_eco58088, w_eco58089, w_eco58090, w_eco58091, w_eco58092, w_eco58093, w_eco58094, w_eco58095, w_eco58096, w_eco58097, w_eco58098, w_eco58099, w_eco58100, w_eco58101, w_eco58102, w_eco58103, w_eco58104, w_eco58105, w_eco58106, w_eco58107, w_eco58108, w_eco58109, w_eco58110, w_eco58111, w_eco58112, w_eco58113, w_eco58114, w_eco58115, w_eco58116, w_eco58117, w_eco58118, w_eco58119, w_eco58120, w_eco58121, w_eco58122, w_eco58123, w_eco58124, w_eco58125, w_eco58126, w_eco58127, w_eco58128, w_eco58129, w_eco58130, w_eco58131, w_eco58132, w_eco58133, w_eco58134, w_eco58135, w_eco58136, w_eco58137, w_eco58138, w_eco58139, w_eco58140, w_eco58141, w_eco58142, w_eco58143, w_eco58144, w_eco58145, w_eco58146, w_eco58147, w_eco58148, w_eco58149, w_eco58150, w_eco58151, w_eco58152, w_eco58153, w_eco58154, w_eco58155, w_eco58156, w_eco58157, w_eco58158, w_eco58159, w_eco58160, w_eco58161, w_eco58162, w_eco58163, w_eco58164, w_eco58165, w_eco58166, w_eco58167, w_eco58168, w_eco58169, w_eco58170, w_eco58171, w_eco58172, w_eco58173, w_eco58174, w_eco58175, w_eco58176, w_eco58177, w_eco58178, w_eco58179, w_eco58180, w_eco58181, w_eco58182, w_eco58183, w_eco58184, w_eco58185, w_eco58186, w_eco58187, w_eco58188, w_eco58189, w_eco58190, w_eco58191, w_eco58192, w_eco58193, w_eco58194, w_eco58195, w_eco58196, w_eco58197, w_eco58198, w_eco58199, w_eco58200, w_eco58201, w_eco58202, w_eco58203, w_eco58204, w_eco58205, w_eco58206, w_eco58207, w_eco58208, w_eco58209, w_eco58210, w_eco58211, w_eco58212, w_eco58213, w_eco58214, w_eco58215, w_eco58216, w_eco58217, w_eco58218, w_eco58219, w_eco58220, w_eco58221, w_eco58222, w_eco58223, w_eco58224, w_eco58225, w_eco58226, w_eco58227, w_eco58228, w_eco58229, w_eco58230, w_eco58231, w_eco58232, w_eco58233, w_eco58234, w_eco58235, w_eco58236, w_eco58237, w_eco58238, w_eco58239, w_eco58240, w_eco58241, w_eco58242, w_eco58243, w_eco58244, w_eco58245, w_eco58246, w_eco58247, w_eco58248, w_eco58249, w_eco58250, w_eco58251, w_eco58252, w_eco58253, w_eco58254, w_eco58255, w_eco58256, w_eco58257, w_eco58258, w_eco58259, w_eco58260, w_eco58261, w_eco58262, w_eco58263, w_eco58264, w_eco58265, w_eco58266, w_eco58267, w_eco58268, w_eco58269, w_eco58270, w_eco58271, w_eco58272, w_eco58273, w_eco58274, w_eco58275, w_eco58276, w_eco58277, w_eco58278, w_eco58279, w_eco58280, w_eco58281, w_eco58282, w_eco58283, w_eco58284, w_eco58285, w_eco58286, w_eco58287, w_eco58288, w_eco58289, w_eco58290, w_eco58291, w_eco58292, w_eco58293, w_eco58294, w_eco58295, w_eco58296, w_eco58297, w_eco58298, w_eco58299, w_eco58300, w_eco58301, w_eco58302, w_eco58303, w_eco58304, w_eco58305, w_eco58306, w_eco58307, w_eco58308, w_eco58309, w_eco58310, w_eco58311, w_eco58312, w_eco58313, w_eco58314, w_eco58315, w_eco58316, w_eco58317, w_eco58318, w_eco58319, w_eco58320, w_eco58321, w_eco58322, w_eco58323, w_eco58324, w_eco58325, w_eco58326, w_eco58327, w_eco58328, w_eco58329, w_eco58330, w_eco58331, w_eco58332, w_eco58333, w_eco58334, w_eco58335, w_eco58336, w_eco58337, w_eco58338, w_eco58339, w_eco58340, w_eco58341, w_eco58342, w_eco58343, w_eco58344, w_eco58345, w_eco58346, w_eco58347, w_eco58348, w_eco58349, w_eco58350, w_eco58351, w_eco58352, w_eco58353, w_eco58354, w_eco58355, w_eco58356, w_eco58357, w_eco58358, w_eco58359, w_eco58360, w_eco58361, w_eco58362, w_eco58363, w_eco58364, w_eco58365, w_eco58366, w_eco58367, w_eco58368, w_eco58369, w_eco58370, w_eco58371, w_eco58372, w_eco58373, w_eco58374, w_eco58375, w_eco58376, w_eco58377, w_eco58378, w_eco58379, w_eco58380, w_eco58381, w_eco58382, w_eco58383, w_eco58384, w_eco58385, w_eco58386, w_eco58387, w_eco58388, w_eco58389, w_eco58390, w_eco58391, w_eco58392, w_eco58393, w_eco58394, w_eco58395, w_eco58396, w_eco58397, w_eco58398, w_eco58399, w_eco58400, w_eco58401, w_eco58402, w_eco58403, w_eco58404, w_eco58405, w_eco58406, w_eco58407, w_eco58408, w_eco58409, w_eco58410, w_eco58411, w_eco58412, w_eco58413, w_eco58414, w_eco58415, w_eco58416, w_eco58417, w_eco58418, w_eco58419, w_eco58420, w_eco58421, w_eco58422, w_eco58423, w_eco58424, w_eco58425, w_eco58426, w_eco58427, w_eco58428, w_eco58429, w_eco58430, w_eco58431, w_eco58432, w_eco58433, w_eco58434, w_eco58435, w_eco58436, w_eco58437, w_eco58438, w_eco58439, w_eco58440, w_eco58441, w_eco58442, w_eco58443, w_eco58444, w_eco58445, w_eco58446, w_eco58447, w_eco58448, w_eco58449, w_eco58450, w_eco58451, w_eco58452, w_eco58453, w_eco58454, w_eco58455, w_eco58456, w_eco58457, w_eco58458, w_eco58459, w_eco58460, w_eco58461, w_eco58462, w_eco58463, w_eco58464, w_eco58465, w_eco58466, w_eco58467, w_eco58468, w_eco58469, w_eco58470, w_eco58471, w_eco58472, w_eco58473, w_eco58474, w_eco58475, w_eco58476, w_eco58477, w_eco58478, w_eco58479, w_eco58480, w_eco58481, w_eco58482, w_eco58483, w_eco58484, w_eco58485, w_eco58486, w_eco58487, w_eco58488, w_eco58489, w_eco58490, w_eco58491, w_eco58492, w_eco58493, w_eco58494, w_eco58495, w_eco58496, w_eco58497, w_eco58498, w_eco58499, w_eco58500, w_eco58501, w_eco58502, w_eco58503, w_eco58504, w_eco58505, w_eco58506, w_eco58507, w_eco58508, w_eco58509, w_eco58510, w_eco58511, w_eco58512, w_eco58513, w_eco58514, w_eco58515, w_eco58516, w_eco58517, w_eco58518, w_eco58519, w_eco58520, w_eco58521, w_eco58522, w_eco58523, w_eco58524, w_eco58525, w_eco58526, w_eco58527, w_eco58528, w_eco58529, w_eco58530, w_eco58531, w_eco58532, w_eco58533, w_eco58534, w_eco58535, w_eco58536, w_eco58537, w_eco58538, w_eco58539, w_eco58540, w_eco58541, w_eco58542, w_eco58543, w_eco58544, w_eco58545, w_eco58546, w_eco58547, w_eco58548, w_eco58549, w_eco58550, w_eco58551, w_eco58552, w_eco58553, w_eco58554, w_eco58555, w_eco58556, w_eco58557, w_eco58558, w_eco58559, w_eco58560, w_eco58561, w_eco58562, w_eco58563, w_eco58564, w_eco58565, w_eco58566, w_eco58567, w_eco58568, w_eco58569, w_eco58570, w_eco58571, w_eco58572, w_eco58573, w_eco58574, w_eco58575, w_eco58576, w_eco58577, w_eco58578, w_eco58579, w_eco58580, w_eco58581, w_eco58582, w_eco58583, w_eco58584, w_eco58585, w_eco58586, w_eco58587, w_eco58588, w_eco58589, w_eco58590, w_eco58591, w_eco58592, w_eco58593, w_eco58594, w_eco58595, w_eco58596, w_eco58597, w_eco58598, w_eco58599, w_eco58600, w_eco58601, w_eco58602, w_eco58603, w_eco58604, w_eco58605, w_eco58606, w_eco58607, w_eco58608, w_eco58609, w_eco58610, w_eco58611, w_eco58612, w_eco58613, w_eco58614, w_eco58615, w_eco58616, w_eco58617, w_eco58618, w_eco58619, w_eco58620, w_eco58621, w_eco58622, w_eco58623, w_eco58624, w_eco58625, w_eco58626, w_eco58627, w_eco58628, w_eco58629, w_eco58630, w_eco58631, w_eco58632, w_eco58633, w_eco58634, w_eco58635, w_eco58636, w_eco58637, w_eco58638, w_eco58639, w_eco58640, w_eco58641, w_eco58642, w_eco58643, w_eco58644, w_eco58645, w_eco58646, w_eco58647, w_eco58648, w_eco58649, w_eco58650, w_eco58651, w_eco58652, w_eco58653, w_eco58654, w_eco58655, w_eco58656, w_eco58657, w_eco58658, w_eco58659, w_eco58660, w_eco58661, w_eco58662, w_eco58663, w_eco58664, w_eco58665, w_eco58666, w_eco58667, w_eco58668, w_eco58669, w_eco58670, w_eco58671, w_eco58672, w_eco58673, w_eco58674, w_eco58675, w_eco58676, w_eco58677, w_eco58678, w_eco58679, w_eco58680, w_eco58681, w_eco58682, w_eco58683, w_eco58684, w_eco58685, w_eco58686, w_eco58687, w_eco58688, w_eco58689, w_eco58690, w_eco58691, w_eco58692, w_eco58693, w_eco58694, w_eco58695, w_eco58696, w_eco58697, w_eco58698, w_eco58699, w_eco58700, w_eco58701, w_eco58702, w_eco58703, w_eco58704, w_eco58705, w_eco58706, w_eco58707, w_eco58708, w_eco58709, w_eco58710, w_eco58711, w_eco58712, w_eco58713, w_eco58714, w_eco58715, w_eco58716, w_eco58717, w_eco58718, w_eco58719, w_eco58720, w_eco58721, w_eco58722, w_eco58723, w_eco58724, w_eco58725, w_eco58726, w_eco58727, w_eco58728, w_eco58729, w_eco58730, w_eco58731, w_eco58732, w_eco58733, w_eco58734, w_eco58735, w_eco58736, w_eco58737, w_eco58738, w_eco58739, w_eco58740, w_eco58741, w_eco58742, w_eco58743, w_eco58744, w_eco58745, w_eco58746, w_eco58747, w_eco58748, w_eco58749, w_eco58750, w_eco58751, w_eco58752, w_eco58753, w_eco58754, w_eco58755, w_eco58756, w_eco58757, w_eco58758, w_eco58759, w_eco58760, w_eco58761, w_eco58762, w_eco58763, w_eco58764, w_eco58765, w_eco58766, w_eco58767, w_eco58768, w_eco58769, w_eco58770, w_eco58771, w_eco58772, w_eco58773, w_eco58774, w_eco58775, w_eco58776, w_eco58777, w_eco58778, w_eco58779, w_eco58780, w_eco58781, w_eco58782, w_eco58783, w_eco58784, w_eco58785, w_eco58786, w_eco58787, w_eco58788, w_eco58789, w_eco58790, w_eco58791, w_eco58792, w_eco58793, w_eco58794, w_eco58795, w_eco58796, w_eco58797, w_eco58798, w_eco58799, w_eco58800, w_eco58801, w_eco58802, w_eco58803, w_eco58804, w_eco58805, w_eco58806, w_eco58807, w_eco58808, w_eco58809, w_eco58810, w_eco58811, w_eco58812, w_eco58813, w_eco58814, w_eco58815, w_eco58816, w_eco58817, w_eco58818, w_eco58819, w_eco58820, w_eco58821, w_eco58822, w_eco58823, w_eco58824, w_eco58825, w_eco58826, w_eco58827, w_eco58828, w_eco58829, w_eco58830, w_eco58831, w_eco58832, w_eco58833, w_eco58834, w_eco58835, w_eco58836, w_eco58837, w_eco58838, w_eco58839, w_eco58840, w_eco58841, w_eco58842, w_eco58843, w_eco58844, w_eco58845, w_eco58846, w_eco58847, w_eco58848, w_eco58849, w_eco58850, w_eco58851, w_eco58852, w_eco58853, w_eco58854, w_eco58855, w_eco58856, w_eco58857, w_eco58858, w_eco58859, w_eco58860, w_eco58861, w_eco58862, w_eco58863, w_eco58864, w_eco58865, w_eco58866, w_eco58867, w_eco58868, w_eco58869, w_eco58870, w_eco58871, w_eco58872, w_eco58873, w_eco58874, w_eco58875, w_eco58876, w_eco58877, w_eco58878, w_eco58879, w_eco58880, w_eco58881, w_eco58882, w_eco58883, w_eco58884, w_eco58885, w_eco58886, w_eco58887, w_eco58888, w_eco58889, w_eco58890, w_eco58891, w_eco58892, w_eco58893, w_eco58894, w_eco58895, w_eco58896, w_eco58897, w_eco58898, w_eco58899, w_eco58900, w_eco58901, w_eco58902, w_eco58903, w_eco58904, w_eco58905, w_eco58906, w_eco58907, w_eco58908, w_eco58909, w_eco58910, w_eco58911, w_eco58912, w_eco58913, w_eco58914, w_eco58915, w_eco58916, w_eco58917, w_eco58918, w_eco58919, w_eco58920, w_eco58921, w_eco58922, w_eco58923, w_eco58924, w_eco58925, w_eco58926, w_eco58927, w_eco58928, w_eco58929, w_eco58930, w_eco58931, w_eco58932, w_eco58933, w_eco58934, w_eco58935, w_eco58936, w_eco58937, w_eco58938, w_eco58939, w_eco58940, w_eco58941, w_eco58942, w_eco58943, w_eco58944, w_eco58945, w_eco58946, w_eco58947, w_eco58948, w_eco58949, w_eco58950, w_eco58951, w_eco58952, w_eco58953, w_eco58954, w_eco58955, w_eco58956, w_eco58957, w_eco58958, w_eco58959, w_eco58960, w_eco58961, w_eco58962, w_eco58963, w_eco58964, w_eco58965, w_eco58966, w_eco58967, w_eco58968, w_eco58969, w_eco58970, w_eco58971, w_eco58972, w_eco58973, w_eco58974, w_eco58975, w_eco58976, w_eco58977, w_eco58978, w_eco58979, w_eco58980, w_eco58981, w_eco58982, w_eco58983, w_eco58984, w_eco58985, w_eco58986, w_eco58987, w_eco58988, w_eco58989, w_eco58990, w_eco58991, w_eco58992, w_eco58993, w_eco58994, w_eco58995, w_eco58996, w_eco58997, w_eco58998, w_eco58999, w_eco59000, w_eco59001, w_eco59002, w_eco59003, w_eco59004, w_eco59005, w_eco59006, w_eco59007, w_eco59008, w_eco59009, w_eco59010, w_eco59011, w_eco59012, w_eco59013, w_eco59014, w_eco59015, w_eco59016, w_eco59017, w_eco59018, w_eco59019, w_eco59020, w_eco59021, w_eco59022, w_eco59023, w_eco59024, w_eco59025, w_eco59026, w_eco59027, w_eco59028, w_eco59029, w_eco59030, w_eco59031, w_eco59032, w_eco59033, w_eco59034, w_eco59035, w_eco59036, w_eco59037, w_eco59038, w_eco59039, w_eco59040, w_eco59041, w_eco59042, w_eco59043, w_eco59044, w_eco59045, w_eco59046, w_eco59047, w_eco59048, w_eco59049, w_eco59050, w_eco59051, w_eco59052, w_eco59053, w_eco59054, w_eco59055, w_eco59056, w_eco59057, w_eco59058, w_eco59059, w_eco59060, w_eco59061, w_eco59062, w_eco59063, w_eco59064, w_eco59065, w_eco59066, w_eco59067, w_eco59068, w_eco59069, w_eco59070, w_eco59071, w_eco59072, w_eco59073, w_eco59074, w_eco59075, w_eco59076, w_eco59077, w_eco59078, w_eco59079, w_eco59080, w_eco59081, w_eco59082, w_eco59083, w_eco59084, w_eco59085, w_eco59086, w_eco59087, w_eco59088, w_eco59089, w_eco59090, w_eco59091, w_eco59092, w_eco59093, w_eco59094, w_eco59095, w_eco59096, w_eco59097, w_eco59098, w_eco59099, w_eco59100, w_eco59101, w_eco59102, w_eco59103, w_eco59104, w_eco59105, w_eco59106, w_eco59107, w_eco59108, w_eco59109, w_eco59110, w_eco59111, w_eco59112, w_eco59113, w_eco59114, w_eco59115, w_eco59116, w_eco59117, w_eco59118, w_eco59119, w_eco59120, w_eco59121, w_eco59122, w_eco59123, w_eco59124, w_eco59125, w_eco59126, w_eco59127, w_eco59128, w_eco59129, w_eco59130, w_eco59131, w_eco59132, w_eco59133, w_eco59134, w_eco59135, w_eco59136, w_eco59137, w_eco59138, w_eco59139, w_eco59140, w_eco59141, w_eco59142, w_eco59143, w_eco59144, w_eco59145, w_eco59146, w_eco59147, w_eco59148, w_eco59149, w_eco59150, w_eco59151, w_eco59152, w_eco59153, w_eco59154, w_eco59155, w_eco59156, w_eco59157, w_eco59158, w_eco59159, w_eco59160, w_eco59161, w_eco59162, w_eco59163, w_eco59164, w_eco59165, w_eco59166, w_eco59167, w_eco59168, w_eco59169, w_eco59170, w_eco59171, w_eco59172, w_eco59173, w_eco59174, w_eco59175, w_eco59176, w_eco59177, w_eco59178, w_eco59179, w_eco59180, w_eco59181, w_eco59182, w_eco59183, w_eco59184, w_eco59185, w_eco59186, w_eco59187, w_eco59188, w_eco59189, w_eco59190, w_eco59191, w_eco59192, w_eco59193, w_eco59194, w_eco59195, w_eco59196, w_eco59197, w_eco59198, w_eco59199, w_eco59200, w_eco59201, w_eco59202, w_eco59203, w_eco59204, w_eco59205, w_eco59206, w_eco59207, w_eco59208, w_eco59209, w_eco59210, w_eco59211, w_eco59212, w_eco59213, w_eco59214, w_eco59215, w_eco59216, w_eco59217, w_eco59218, w_eco59219, w_eco59220, w_eco59221, w_eco59222, w_eco59223, w_eco59224, w_eco59225, w_eco59226, w_eco59227, w_eco59228, w_eco59229, w_eco59230, w_eco59231, w_eco59232, w_eco59233, w_eco59234, w_eco59235, w_eco59236, w_eco59237, w_eco59238, w_eco59239, w_eco59240, w_eco59241, w_eco59242, w_eco59243, w_eco59244, w_eco59245, w_eco59246, w_eco59247, w_eco59248, w_eco59249, w_eco59250, w_eco59251, w_eco59252, w_eco59253, w_eco59254, w_eco59255, w_eco59256, w_eco59257, w_eco59258, w_eco59259, w_eco59260, w_eco59261, w_eco59262, w_eco59263, w_eco59264, w_eco59265, w_eco59266, w_eco59267, w_eco59268, w_eco59269, w_eco59270, w_eco59271, w_eco59272, w_eco59273, w_eco59274, w_eco59275, w_eco59276, w_eco59277, w_eco59278, w_eco59279, w_eco59280, w_eco59281, w_eco59282, w_eco59283, w_eco59284, w_eco59285, w_eco59286, w_eco59287, w_eco59288, w_eco59289, w_eco59290, w_eco59291, w_eco59292, w_eco59293, w_eco59294, w_eco59295, w_eco59296, w_eco59297, w_eco59298, w_eco59299, w_eco59300, w_eco59301, w_eco59302, w_eco59303, w_eco59304, w_eco59305, w_eco59306, w_eco59307, w_eco59308, w_eco59309, w_eco59310, w_eco59311, w_eco59312, w_eco59313, w_eco59314, w_eco59315, w_eco59316, w_eco59317, w_eco59318, w_eco59319, w_eco59320, w_eco59321, w_eco59322, w_eco59323, w_eco59324, w_eco59325, w_eco59326, w_eco59327, w_eco59328, w_eco59329, w_eco59330, w_eco59331, w_eco59332, w_eco59333, w_eco59334, w_eco59335, w_eco59336, w_eco59337, w_eco59338, w_eco59339, w_eco59340, w_eco59341, w_eco59342, w_eco59343, w_eco59344, w_eco59345, w_eco59346, w_eco59347, w_eco59348, w_eco59349, w_eco59350, w_eco59351, w_eco59352, w_eco59353, w_eco59354, w_eco59355, w_eco59356, w_eco59357, w_eco59358, w_eco59359, w_eco59360, w_eco59361, w_eco59362, w_eco59363, w_eco59364, w_eco59365, w_eco59366, w_eco59367, w_eco59368, w_eco59369, w_eco59370, w_eco59371, w_eco59372, w_eco59373, w_eco59374, w_eco59375, w_eco59376, w_eco59377, w_eco59378, w_eco59379, w_eco59380, w_eco59381, w_eco59382, w_eco59383, w_eco59384, w_eco59385, w_eco59386, w_eco59387, w_eco59388, w_eco59389, w_eco59390, w_eco59391, w_eco59392, w_eco59393, w_eco59394, w_eco59395, w_eco59396, w_eco59397, w_eco59398, w_eco59399, w_eco59400, w_eco59401, w_eco59402, w_eco59403, w_eco59404, w_eco59405, w_eco59406, w_eco59407, w_eco59408, w_eco59409, w_eco59410, w_eco59411, w_eco59412, w_eco59413, w_eco59414, w_eco59415, w_eco59416, w_eco59417, w_eco59418, w_eco59419, w_eco59420, w_eco59421, w_eco59422, w_eco59423, w_eco59424, w_eco59425, w_eco59426, w_eco59427, w_eco59428, w_eco59429, w_eco59430, w_eco59431, w_eco59432, w_eco59433, w_eco59434, w_eco59435, w_eco59436, w_eco59437, w_eco59438, w_eco59439, w_eco59440, w_eco59441, w_eco59442, w_eco59443, w_eco59444, w_eco59445, w_eco59446, w_eco59447, w_eco59448, w_eco59449, w_eco59450, w_eco59451, w_eco59452, w_eco59453, w_eco59454, w_eco59455, w_eco59456, w_eco59457, w_eco59458, w_eco59459, w_eco59460, w_eco59461, w_eco59462, w_eco59463, w_eco59464, w_eco59465, w_eco59466, w_eco59467, w_eco59468, w_eco59469, w_eco59470, w_eco59471, w_eco59472, w_eco59473, w_eco59474, w_eco59475, w_eco59476, w_eco59477, w_eco59478, w_eco59479, w_eco59480, w_eco59481, w_eco59482, w_eco59483, w_eco59484, w_eco59485, w_eco59486, w_eco59487, w_eco59488, w_eco59489, w_eco59490, w_eco59491, w_eco59492, w_eco59493, w_eco59494, w_eco59495, w_eco59496, w_eco59497, w_eco59498, w_eco59499, w_eco59500, w_eco59501, w_eco59502, w_eco59503, w_eco59504, w_eco59505, w_eco59506, w_eco59507, w_eco59508, w_eco59509, w_eco59510, w_eco59511, w_eco59512, w_eco59513, w_eco59514, w_eco59515, w_eco59516, w_eco59517, w_eco59518, w_eco59519, w_eco59520, w_eco59521, w_eco59522, w_eco59523, w_eco59524, w_eco59525, w_eco59526, w_eco59527, w_eco59528, w_eco59529, w_eco59530, w_eco59531, w_eco59532, w_eco59533, w_eco59534, w_eco59535, w_eco59536, w_eco59537, w_eco59538, w_eco59539, w_eco59540, w_eco59541, w_eco59542, w_eco59543, w_eco59544, w_eco59545, w_eco59546, w_eco59547, w_eco59548, w_eco59549, w_eco59550, w_eco59551, w_eco59552, w_eco59553, w_eco59554, w_eco59555, w_eco59556, w_eco59557, w_eco59558, w_eco59559, w_eco59560, w_eco59561, w_eco59562, w_eco59563, w_eco59564, w_eco59565, w_eco59566, w_eco59567, w_eco59568, w_eco59569, w_eco59570, w_eco59571, w_eco59572, w_eco59573, w_eco59574, w_eco59575, w_eco59576, w_eco59577, w_eco59578, w_eco59579, w_eco59580, w_eco59581, w_eco59582, w_eco59583, w_eco59584, w_eco59585, w_eco59586, w_eco59587, w_eco59588, w_eco59589, w_eco59590, w_eco59591, w_eco59592, w_eco59593, w_eco59594, w_eco59595, w_eco59596, w_eco59597, w_eco59598, w_eco59599, w_eco59600, w_eco59601, w_eco59602, w_eco59603, w_eco59604, w_eco59605, w_eco59606, w_eco59607, w_eco59608, w_eco59609, w_eco59610, w_eco59611, w_eco59612, w_eco59613, w_eco59614, w_eco59615, w_eco59616, w_eco59617, w_eco59618, w_eco59619, w_eco59620, w_eco59621, w_eco59622, w_eco59623, w_eco59624, w_eco59625, w_eco59626, w_eco59627, w_eco59628, w_eco59629, w_eco59630, w_eco59631, w_eco59632, w_eco59633, w_eco59634, w_eco59635, w_eco59636, w_eco59637, w_eco59638, w_eco59639, w_eco59640, w_eco59641, w_eco59642, w_eco59643, w_eco59644, w_eco59645, w_eco59646, w_eco59647, w_eco59648, w_eco59649, w_eco59650, w_eco59651, w_eco59652, w_eco59653, w_eco59654, w_eco59655, w_eco59656, w_eco59657, w_eco59658, w_eco59659, w_eco59660, w_eco59661, w_eco59662, w_eco59663, w_eco59664, w_eco59665, w_eco59666, w_eco59667, w_eco59668, w_eco59669, w_eco59670, w_eco59671, w_eco59672, w_eco59673, w_eco59674, w_eco59675, w_eco59676, w_eco59677, w_eco59678, w_eco59679, w_eco59680, w_eco59681, w_eco59682, w_eco59683, w_eco59684, w_eco59685, w_eco59686, w_eco59687, w_eco59688, w_eco59689, w_eco59690, w_eco59691, w_eco59692, w_eco59693, w_eco59694, w_eco59695, w_eco59696, w_eco59697, w_eco59698, w_eco59699, w_eco59700, w_eco59701, w_eco59702, w_eco59703, w_eco59704, w_eco59705, w_eco59706, w_eco59707, w_eco59708, w_eco59709, w_eco59710, w_eco59711, w_eco59712, w_eco59713, w_eco59714, w_eco59715, w_eco59716, w_eco59717, w_eco59718, w_eco59719, w_eco59720, w_eco59721, w_eco59722, w_eco59723, w_eco59724, w_eco59725, w_eco59726, w_eco59727, w_eco59728, w_eco59729, w_eco59730, w_eco59731, w_eco59732, w_eco59733, w_eco59734, w_eco59735, w_eco59736, w_eco59737, w_eco59738, w_eco59739, w_eco59740, w_eco59741, w_eco59742, w_eco59743, w_eco59744, w_eco59745, w_eco59746, w_eco59747, w_eco59748, w_eco59749, w_eco59750, w_eco59751, w_eco59752, w_eco59753, w_eco59754, w_eco59755, w_eco59756, w_eco59757, w_eco59758, w_eco59759, w_eco59760, w_eco59761, w_eco59762, w_eco59763, w_eco59764, w_eco59765, w_eco59766, w_eco59767, w_eco59768, w_eco59769, w_eco59770, w_eco59771, w_eco59772, w_eco59773, w_eco59774, w_eco59775, w_eco59776, w_eco59777, w_eco59778, w_eco59779, w_eco59780, w_eco59781, w_eco59782, w_eco59783, w_eco59784, w_eco59785, w_eco59786, w_eco59787, w_eco59788, w_eco59789, w_eco59790, w_eco59791, w_eco59792, w_eco59793, w_eco59794, w_eco59795, w_eco59796, w_eco59797, w_eco59798, w_eco59799, w_eco59800, w_eco59801, w_eco59802, w_eco59803, w_eco59804, w_eco59805, w_eco59806, w_eco59807, w_eco59808, w_eco59809, w_eco59810, w_eco59811, w_eco59812, w_eco59813, w_eco59814, w_eco59815, w_eco59816, w_eco59817, w_eco59818, w_eco59819, w_eco59820, w_eco59821, w_eco59822, w_eco59823, w_eco59824, w_eco59825, w_eco59826, w_eco59827, w_eco59828, w_eco59829, w_eco59830, w_eco59831, w_eco59832, w_eco59833, w_eco59834, w_eco59835, w_eco59836, w_eco59837, w_eco59838, w_eco59839, w_eco59840, w_eco59841, w_eco59842, w_eco59843, w_eco59844, w_eco59845, w_eco59846, w_eco59847, w_eco59848, w_eco59849, w_eco59850, w_eco59851, w_eco59852, w_eco59853, w_eco59854, w_eco59855, w_eco59856, w_eco59857, w_eco59858, w_eco59859, w_eco59860, w_eco59861, w_eco59862, w_eco59863, w_eco59864, w_eco59865, w_eco59866, w_eco59867, w_eco59868, w_eco59869, w_eco59870, w_eco59871, w_eco59872, w_eco59873, w_eco59874, w_eco59875, w_eco59876, w_eco59877, w_eco59878, w_eco59879, w_eco59880, w_eco59881, w_eco59882, w_eco59883, w_eco59884, w_eco59885, w_eco59886, w_eco59887, w_eco59888, w_eco59889, w_eco59890, w_eco59891, w_eco59892, w_eco59893, w_eco59894, w_eco59895, w_eco59896, w_eco59897, w_eco59898, w_eco59899, w_eco59900, w_eco59901, w_eco59902, w_eco59903, w_eco59904, w_eco59905, w_eco59906, w_eco59907, w_eco59908, w_eco59909, w_eco59910, w_eco59911, w_eco59912, w_eco59913, w_eco59914, w_eco59915, w_eco59916, w_eco59917, w_eco59918, w_eco59919, w_eco59920, w_eco59921, w_eco59922, w_eco59923, w_eco59924, w_eco59925, w_eco59926, w_eco59927, w_eco59928, w_eco59929, w_eco59930, w_eco59931, w_eco59932, w_eco59933, w_eco59934, w_eco59935, w_eco59936, w_eco59937, w_eco59938, w_eco59939, w_eco59940, w_eco59941, w_eco59942, w_eco59943, w_eco59944, w_eco59945, w_eco59946, w_eco59947, w_eco59948, w_eco59949, w_eco59950, w_eco59951, w_eco59952, w_eco59953, w_eco59954, w_eco59955, w_eco59956, w_eco59957, w_eco59958, w_eco59959, w_eco59960, w_eco59961, w_eco59962, w_eco59963, w_eco59964, w_eco59965, w_eco59966, w_eco59967, w_eco59968, w_eco59969, w_eco59970, w_eco59971, w_eco59972, w_eco59973, w_eco59974, w_eco59975, w_eco59976, w_eco59977, w_eco59978, w_eco59979, w_eco59980, w_eco59981, w_eco59982, w_eco59983, w_eco59984, w_eco59985, w_eco59986, w_eco59987, w_eco59988, w_eco59989, w_eco59990, w_eco59991, w_eco59992, w_eco59993, w_eco59994, w_eco59995, w_eco59996, w_eco59997, w_eco59998, w_eco59999, w_eco60000, w_eco60001, w_eco60002, w_eco60003, w_eco60004, w_eco60005, w_eco60006, w_eco60007, w_eco60008, w_eco60009, w_eco60010, w_eco60011, w_eco60012, w_eco60013, w_eco60014, w_eco60015, w_eco60016, w_eco60017, w_eco60018, w_eco60019, w_eco60020, w_eco60021, w_eco60022, w_eco60023, w_eco60024, w_eco60025, w_eco60026, w_eco60027, w_eco60028, w_eco60029, w_eco60030, w_eco60031, w_eco60032, w_eco60033, w_eco60034, w_eco60035, w_eco60036, w_eco60037, w_eco60038, w_eco60039, w_eco60040, w_eco60041, w_eco60042, w_eco60043, w_eco60044, w_eco60045, w_eco60046, w_eco60047, w_eco60048, w_eco60049, w_eco60050, w_eco60051, w_eco60052, w_eco60053, w_eco60054, w_eco60055, w_eco60056, w_eco60057, w_eco60058, w_eco60059, w_eco60060, w_eco60061, w_eco60062, w_eco60063, w_eco60064, w_eco60065, w_eco60066, w_eco60067, w_eco60068, w_eco60069, w_eco60070, w_eco60071, w_eco60072, w_eco60073, w_eco60074, w_eco60075, w_eco60076, w_eco60077, w_eco60078, w_eco60079, w_eco60080, w_eco60081, w_eco60082, w_eco60083, w_eco60084, w_eco60085, w_eco60086, w_eco60087, w_eco60088, w_eco60089, w_eco60090, w_eco60091, w_eco60092, w_eco60093, w_eco60094, w_eco60095, w_eco60096, w_eco60097, w_eco60098, w_eco60099, w_eco60100, w_eco60101, w_eco60102, w_eco60103, w_eco60104, w_eco60105, w_eco60106, w_eco60107, w_eco60108, w_eco60109, w_eco60110, w_eco60111, w_eco60112, w_eco60113, w_eco60114, w_eco60115, w_eco60116, w_eco60117, w_eco60118, w_eco60119, w_eco60120, w_eco60121, w_eco60122, w_eco60123, w_eco60124, w_eco60125, w_eco60126, w_eco60127, w_eco60128, w_eco60129, w_eco60130, w_eco60131, w_eco60132, w_eco60133, w_eco60134, w_eco60135, w_eco60136, w_eco60137, w_eco60138, w_eco60139, w_eco60140, w_eco60141, w_eco60142, w_eco60143, w_eco60144, w_eco60145, w_eco60146, w_eco60147, w_eco60148, w_eco60149, w_eco60150, w_eco60151, w_eco60152, w_eco60153, w_eco60154, w_eco60155, w_eco60156, w_eco60157, w_eco60158, w_eco60159, w_eco60160, w_eco60161, w_eco60162, w_eco60163, w_eco60164, w_eco60165, w_eco60166, w_eco60167, w_eco60168, w_eco60169, w_eco60170, w_eco60171, w_eco60172, w_eco60173, w_eco60174, w_eco60175, w_eco60176, w_eco60177, w_eco60178, w_eco60179, w_eco60180, w_eco60181, w_eco60182, w_eco60183, w_eco60184, w_eco60185, w_eco60186, w_eco60187, w_eco60188, w_eco60189, w_eco60190, w_eco60191, w_eco60192, w_eco60193, w_eco60194, w_eco60195, w_eco60196, w_eco60197, w_eco60198, w_eco60199, w_eco60200, w_eco60201, w_eco60202, w_eco60203, w_eco60204, w_eco60205, w_eco60206, w_eco60207, w_eco60208, w_eco60209, w_eco60210, w_eco60211, w_eco60212, w_eco60213, w_eco60214, w_eco60215, w_eco60216, w_eco60217, w_eco60218, w_eco60219, w_eco60220, w_eco60221, w_eco60222, w_eco60223, w_eco60224, w_eco60225, w_eco60226, w_eco60227, w_eco60228, w_eco60229, w_eco60230, w_eco60231, w_eco60232, w_eco60233, w_eco60234, w_eco60235, w_eco60236, w_eco60237, w_eco60238, w_eco60239, w_eco60240, w_eco60241, w_eco60242, w_eco60243, w_eco60244, w_eco60245, w_eco60246, w_eco60247, w_eco60248, w_eco60249, w_eco60250, w_eco60251, w_eco60252, w_eco60253, w_eco60254, w_eco60255, w_eco60256, w_eco60257, w_eco60258, w_eco60259, w_eco60260, w_eco60261, w_eco60262, w_eco60263, w_eco60264, w_eco60265, w_eco60266, w_eco60267, w_eco60268, w_eco60269, w_eco60270, w_eco60271, w_eco60272, w_eco60273, w_eco60274, w_eco60275, w_eco60276, w_eco60277, w_eco60278, w_eco60279, w_eco60280, w_eco60281, w_eco60282, w_eco60283, w_eco60284, w_eco60285, w_eco60286, w_eco60287, w_eco60288, w_eco60289, w_eco60290, w_eco60291, w_eco60292, w_eco60293, w_eco60294, w_eco60295, w_eco60296, w_eco60297, w_eco60298, w_eco60299, w_eco60300, w_eco60301, w_eco60302, w_eco60303, w_eco60304, w_eco60305, w_eco60306, w_eco60307, w_eco60308, w_eco60309, w_eco60310, w_eco60311, w_eco60312, w_eco60313, w_eco60314, w_eco60315, w_eco60316, w_eco60317, w_eco60318, w_eco60319, w_eco60320, w_eco60321, w_eco60322, w_eco60323, w_eco60324, w_eco60325, w_eco60326, w_eco60327, w_eco60328, w_eco60329, w_eco60330, w_eco60331, w_eco60332, w_eco60333, w_eco60334, w_eco60335, w_eco60336, w_eco60337, w_eco60338, w_eco60339, w_eco60340, w_eco60341, w_eco60342, w_eco60343, w_eco60344, w_eco60345, w_eco60346, w_eco60347, w_eco60348, w_eco60349, w_eco60350, w_eco60351, w_eco60352, w_eco60353, w_eco60354, w_eco60355, w_eco60356, w_eco60357, w_eco60358, w_eco60359, w_eco60360, w_eco60361, w_eco60362, w_eco60363, w_eco60364, w_eco60365, w_eco60366, w_eco60367, w_eco60368, w_eco60369, w_eco60370, w_eco60371, w_eco60372, w_eco60373, w_eco60374, w_eco60375, w_eco60376, w_eco60377, w_eco60378, w_eco60379, w_eco60380, w_eco60381, w_eco60382, w_eco60383, w_eco60384, w_eco60385, w_eco60386, w_eco60387, w_eco60388, w_eco60389, w_eco60390, w_eco60391, w_eco60392, w_eco60393, w_eco60394, w_eco60395, w_eco60396, w_eco60397, w_eco60398, w_eco60399, w_eco60400, w_eco60401, w_eco60402, w_eco60403, w_eco60404, w_eco60405, w_eco60406, w_eco60407, w_eco60408, w_eco60409, w_eco60410, w_eco60411, w_eco60412, w_eco60413, w_eco60414, w_eco60415, w_eco60416, w_eco60417, w_eco60418, w_eco60419, w_eco60420, w_eco60421, w_eco60422, w_eco60423, w_eco60424, w_eco60425, w_eco60426, w_eco60427, w_eco60428, w_eco60429, w_eco60430, w_eco60431, w_eco60432, w_eco60433, w_eco60434, w_eco60435, w_eco60436, w_eco60437, w_eco60438, w_eco60439, w_eco60440, w_eco60441, w_eco60442, w_eco60443, w_eco60444, w_eco60445, w_eco60446, w_eco60447, w_eco60448, w_eco60449, w_eco60450, w_eco60451, w_eco60452, w_eco60453, w_eco60454, w_eco60455, w_eco60456, w_eco60457, w_eco60458, w_eco60459, w_eco60460, w_eco60461, w_eco60462, w_eco60463, w_eco60464, w_eco60465, w_eco60466, w_eco60467, w_eco60468, w_eco60469, w_eco60470, w_eco60471, w_eco60472, w_eco60473, w_eco60474, w_eco60475, w_eco60476, w_eco60477, w_eco60478, w_eco60479, w_eco60480, w_eco60481, w_eco60482, w_eco60483, w_eco60484, w_eco60485, w_eco60486, w_eco60487, w_eco60488, w_eco60489, w_eco60490, w_eco60491, w_eco60492, w_eco60493, w_eco60494, w_eco60495, w_eco60496, w_eco60497, w_eco60498, w_eco60499, w_eco60500, w_eco60501, w_eco60502, w_eco60503, w_eco60504, w_eco60505, w_eco60506, w_eco60507, w_eco60508, w_eco60509, w_eco60510, w_eco60511, w_eco60512, w_eco60513, w_eco60514, w_eco60515, w_eco60516, w_eco60517, w_eco60518, w_eco60519, w_eco60520, w_eco60521, w_eco60522, w_eco60523, w_eco60524, w_eco60525, w_eco60526, w_eco60527, w_eco60528, w_eco60529, w_eco60530, w_eco60531, w_eco60532, w_eco60533, w_eco60534, w_eco60535, w_eco60536, w_eco60537, w_eco60538, w_eco60539, w_eco60540, w_eco60541, w_eco60542, w_eco60543, w_eco60544, w_eco60545, w_eco60546, w_eco60547, w_eco60548, w_eco60549, w_eco60550, w_eco60551, w_eco60552, w_eco60553, w_eco60554, w_eco60555, w_eco60556, w_eco60557, w_eco60558, w_eco60559, w_eco60560, w_eco60561, w_eco60562, w_eco60563, w_eco60564, w_eco60565, w_eco60566, w_eco60567, w_eco60568, w_eco60569, w_eco60570, w_eco60571, w_eco60572, w_eco60573, w_eco60574, w_eco60575, w_eco60576, w_eco60577, w_eco60578, w_eco60579, w_eco60580, w_eco60581, w_eco60582, w_eco60583, w_eco60584, w_eco60585, w_eco60586, w_eco60587, w_eco60588, w_eco60589, w_eco60590, w_eco60591, w_eco60592, w_eco60593, w_eco60594, w_eco60595, w_eco60596, w_eco60597, w_eco60598, w_eco60599, w_eco60600, w_eco60601, w_eco60602, w_eco60603, w_eco60604, w_eco60605, w_eco60606, w_eco60607, w_eco60608, w_eco60609, w_eco60610, w_eco60611, w_eco60612, w_eco60613, w_eco60614, w_eco60615, w_eco60616, w_eco60617, w_eco60618, w_eco60619, w_eco60620, w_eco60621, w_eco60622, w_eco60623, w_eco60624, w_eco60625, w_eco60626, w_eco60627, w_eco60628, w_eco60629, w_eco60630, w_eco60631, w_eco60632, w_eco60633, w_eco60634, w_eco60635, w_eco60636, w_eco60637, w_eco60638, w_eco60639, w_eco60640, w_eco60641, w_eco60642, w_eco60643, w_eco60644, w_eco60645, w_eco60646, w_eco60647, w_eco60648, w_eco60649, w_eco60650, w_eco60651, w_eco60652, w_eco60653, w_eco60654, w_eco60655, w_eco60656, w_eco60657, w_eco60658, w_eco60659, w_eco60660, w_eco60661, w_eco60662, w_eco60663, w_eco60664, w_eco60665, w_eco60666, w_eco60667, w_eco60668, w_eco60669, w_eco60670, w_eco60671, w_eco60672, w_eco60673, w_eco60674, w_eco60675, w_eco60676, w_eco60677, w_eco60678, w_eco60679, w_eco60680, w_eco60681, w_eco60682, w_eco60683, w_eco60684, w_eco60685, w_eco60686, w_eco60687, w_eco60688, w_eco60689, w_eco60690, w_eco60691, w_eco60692, w_eco60693, w_eco60694, w_eco60695, w_eco60696, w_eco60697, w_eco60698, w_eco60699, w_eco60700, w_eco60701, w_eco60702, w_eco60703, w_eco60704, w_eco60705, w_eco60706, w_eco60707, w_eco60708, w_eco60709, w_eco60710, w_eco60711, w_eco60712, w_eco60713, w_eco60714, w_eco60715, w_eco60716, w_eco60717, w_eco60718, w_eco60719, w_eco60720, w_eco60721, w_eco60722, w_eco60723, w_eco60724, w_eco60725, w_eco60726, w_eco60727, w_eco60728, w_eco60729, w_eco60730, w_eco60731, w_eco60732, w_eco60733, w_eco60734, w_eco60735, w_eco60736, w_eco60737, w_eco60738, w_eco60739, w_eco60740, w_eco60741, w_eco60742, w_eco60743, w_eco60744, w_eco60745, w_eco60746, w_eco60747, w_eco60748, w_eco60749, w_eco60750, w_eco60751, w_eco60752, w_eco60753, w_eco60754, w_eco60755, w_eco60756, w_eco60757, w_eco60758, w_eco60759, w_eco60760, w_eco60761, w_eco60762, w_eco60763, w_eco60764, w_eco60765, w_eco60766, w_eco60767, w_eco60768, w_eco60769, w_eco60770, w_eco60771, w_eco60772, w_eco60773, w_eco60774, w_eco60775, w_eco60776, w_eco60777, w_eco60778, w_eco60779, w_eco60780, w_eco60781, w_eco60782, w_eco60783, w_eco60784, w_eco60785, w_eco60786, w_eco60787, w_eco60788, w_eco60789, w_eco60790, w_eco60791, w_eco60792, w_eco60793, w_eco60794, w_eco60795, w_eco60796, w_eco60797, w_eco60798, w_eco60799, w_eco60800, w_eco60801, w_eco60802, w_eco60803, w_eco60804, w_eco60805, w_eco60806, w_eco60807, w_eco60808, w_eco60809, w_eco60810, w_eco60811, w_eco60812, w_eco60813, w_eco60814, w_eco60815, w_eco60816, w_eco60817, w_eco60818, w_eco60819, w_eco60820, w_eco60821, w_eco60822, w_eco60823, w_eco60824, w_eco60825, w_eco60826, w_eco60827, w_eco60828, w_eco60829, w_eco60830, w_eco60831, w_eco60832, w_eco60833, w_eco60834, w_eco60835, w_eco60836, w_eco60837, w_eco60838, w_eco60839, w_eco60840, w_eco60841, w_eco60842, w_eco60843, w_eco60844, w_eco60845, w_eco60846, w_eco60847, w_eco60848, w_eco60849, w_eco60850, w_eco60851, w_eco60852, w_eco60853, w_eco60854, w_eco60855, w_eco60856, w_eco60857, w_eco60858, w_eco60859, w_eco60860, w_eco60861, w_eco60862, w_eco60863, w_eco60864, w_eco60865, w_eco60866, w_eco60867, w_eco60868, w_eco60869, w_eco60870, w_eco60871, w_eco60872, w_eco60873, w_eco60874, w_eco60875, w_eco60876, w_eco60877, w_eco60878, w_eco60879, w_eco60880, w_eco60881, w_eco60882, w_eco60883, w_eco60884, w_eco60885, w_eco60886, w_eco60887, w_eco60888, w_eco60889, w_eco60890, w_eco60891, w_eco60892, w_eco60893, w_eco60894, w_eco60895, w_eco60896, w_eco60897, w_eco60898, w_eco60899, w_eco60900, w_eco60901, w_eco60902, w_eco60903, w_eco60904, w_eco60905, w_eco60906, w_eco60907, w_eco60908, w_eco60909, w_eco60910, w_eco60911, w_eco60912, w_eco60913, w_eco60914, w_eco60915, w_eco60916, w_eco60917, w_eco60918, w_eco60919, w_eco60920, w_eco60921, w_eco60922, w_eco60923, w_eco60924, w_eco60925, w_eco60926, w_eco60927, w_eco60928, w_eco60929, w_eco60930, w_eco60931, w_eco60932, w_eco60933, w_eco60934, w_eco60935, w_eco60936, w_eco60937, w_eco60938, w_eco60939, w_eco60940, w_eco60941, w_eco60942, w_eco60943, w_eco60944, w_eco60945, w_eco60946, w_eco60947, w_eco60948, w_eco60949, w_eco60950, w_eco60951, w_eco60952, w_eco60953, w_eco60954, w_eco60955, w_eco60956, w_eco60957, w_eco60958, w_eco60959, w_eco60960, w_eco60961, w_eco60962, w_eco60963, w_eco60964, w_eco60965, w_eco60966, w_eco60967, w_eco60968, w_eco60969, w_eco60970, w_eco60971, w_eco60972, w_eco60973, w_eco60974, w_eco60975, w_eco60976, w_eco60977, w_eco60978, w_eco60979, w_eco60980, w_eco60981, w_eco60982, w_eco60983, w_eco60984, w_eco60985, w_eco60986, w_eco60987, w_eco60988, w_eco60989, w_eco60990, w_eco60991, w_eco60992, w_eco60993, w_eco60994, w_eco60995, w_eco60996, w_eco60997, w_eco60998, w_eco60999, w_eco61000, w_eco61001, w_eco61002, w_eco61003, w_eco61004, w_eco61005, w_eco61006, w_eco61007, w_eco61008, w_eco61009, w_eco61010, w_eco61011, w_eco61012, w_eco61013, w_eco61014, w_eco61015, w_eco61016, w_eco61017, w_eco61018, w_eco61019, w_eco61020, w_eco61021, w_eco61022, w_eco61023, w_eco61024, w_eco61025, w_eco61026, w_eco61027, w_eco61028, w_eco61029, w_eco61030, w_eco61031, w_eco61032, w_eco61033, w_eco61034, w_eco61035, w_eco61036, w_eco61037, w_eco61038, w_eco61039, w_eco61040, w_eco61041, w_eco61042, w_eco61043, w_eco61044, w_eco61045, w_eco61046, w_eco61047, w_eco61048, w_eco61049, w_eco61050, w_eco61051, w_eco61052, w_eco61053, w_eco61054, w_eco61055, w_eco61056, w_eco61057, w_eco61058, w_eco61059, w_eco61060, w_eco61061, w_eco61062, w_eco61063, w_eco61064, w_eco61065, w_eco61066, w_eco61067, w_eco61068, w_eco61069, w_eco61070, w_eco61071, w_eco61072, w_eco61073, w_eco61074, w_eco61075, w_eco61076, w_eco61077, w_eco61078, w_eco61079, w_eco61080, w_eco61081, w_eco61082, w_eco61083, w_eco61084, w_eco61085, w_eco61086, w_eco61087, w_eco61088, w_eco61089, w_eco61090, w_eco61091, w_eco61092, w_eco61093, w_eco61094, w_eco61095, w_eco61096, w_eco61097, w_eco61098, w_eco61099, w_eco61100, w_eco61101, w_eco61102, w_eco61103, w_eco61104, w_eco61105, w_eco61106, w_eco61107, w_eco61108, w_eco61109, w_eco61110, w_eco61111, w_eco61112, w_eco61113, w_eco61114, w_eco61115, w_eco61116, w_eco61117, w_eco61118, w_eco61119, w_eco61120, w_eco61121, w_eco61122, w_eco61123, w_eco61124, w_eco61125, w_eco61126, w_eco61127, w_eco61128, w_eco61129, w_eco61130, w_eco61131, w_eco61132, w_eco61133, w_eco61134, w_eco61135, w_eco61136, w_eco61137, w_eco61138, w_eco61139, w_eco61140, w_eco61141, w_eco61142, w_eco61143, w_eco61144, w_eco61145, w_eco61146, w_eco61147, w_eco61148, w_eco61149, w_eco61150, w_eco61151, w_eco61152, w_eco61153, w_eco61154, w_eco61155, w_eco61156, w_eco61157, w_eco61158, w_eco61159, w_eco61160, w_eco61161, w_eco61162, w_eco61163, w_eco61164, w_eco61165, w_eco61166, w_eco61167, w_eco61168, w_eco61169, w_eco61170, w_eco61171, w_eco61172, w_eco61173, w_eco61174, w_eco61175, w_eco61176, w_eco61177, w_eco61178, w_eco61179, w_eco61180, w_eco61181, w_eco61182, w_eco61183, w_eco61184, w_eco61185, w_eco61186, w_eco61187, w_eco61188, w_eco61189, w_eco61190, w_eco61191, w_eco61192, w_eco61193, w_eco61194, w_eco61195, w_eco61196, w_eco61197, w_eco61198, w_eco61199, w_eco61200, w_eco61201, w_eco61202, w_eco61203, w_eco61204, w_eco61205, w_eco61206, w_eco61207, w_eco61208, w_eco61209, w_eco61210, w_eco61211, w_eco61212, w_eco61213, w_eco61214, w_eco61215, w_eco61216, w_eco61217, w_eco61218, w_eco61219, w_eco61220, w_eco61221, w_eco61222, w_eco61223, w_eco61224, w_eco61225, w_eco61226, w_eco61227, w_eco61228, w_eco61229, w_eco61230, w_eco61231, w_eco61232, w_eco61233, w_eco61234, w_eco61235, w_eco61236, w_eco61237, w_eco61238, w_eco61239, w_eco61240, w_eco61241, w_eco61242, w_eco61243, w_eco61244, w_eco61245, w_eco61246, w_eco61247, w_eco61248, w_eco61249, w_eco61250, w_eco61251, w_eco61252, w_eco61253, w_eco61254, w_eco61255, w_eco61256, w_eco61257, w_eco61258, w_eco61259, w_eco61260, w_eco61261, w_eco61262, w_eco61263, w_eco61264, w_eco61265, w_eco61266, w_eco61267, w_eco61268, w_eco61269, w_eco61270, w_eco61271, w_eco61272, w_eco61273, w_eco61274, w_eco61275, w_eco61276, w_eco61277, w_eco61278, w_eco61279, w_eco61280, w_eco61281, w_eco61282, w_eco61283, w_eco61284, w_eco61285, w_eco61286, w_eco61287, w_eco61288, w_eco61289, w_eco61290, w_eco61291, w_eco61292, w_eco61293, w_eco61294, w_eco61295, w_eco61296, w_eco61297, w_eco61298, w_eco61299, w_eco61300, w_eco61301, w_eco61302, w_eco61303, w_eco61304, w_eco61305, w_eco61306, w_eco61307, w_eco61308, w_eco61309, w_eco61310, w_eco61311, w_eco61312, w_eco61313, w_eco61314, w_eco61315, w_eco61316, w_eco61317, w_eco61318, w_eco61319, w_eco61320, w_eco61321, w_eco61322, w_eco61323, w_eco61324, w_eco61325, w_eco61326, w_eco61327, w_eco61328, w_eco61329, w_eco61330, w_eco61331, w_eco61332, w_eco61333, w_eco61334, w_eco61335, w_eco61336, w_eco61337, w_eco61338, w_eco61339, w_eco61340, w_eco61341, w_eco61342, w_eco61343, w_eco61344, w_eco61345, w_eco61346, w_eco61347, w_eco61348, w_eco61349, w_eco61350, w_eco61351, w_eco61352, w_eco61353, w_eco61354, w_eco61355, w_eco61356, w_eco61357, w_eco61358, w_eco61359, w_eco61360, w_eco61361, w_eco61362, w_eco61363, w_eco61364, w_eco61365, w_eco61366, w_eco61367, w_eco61368, w_eco61369, w_eco61370, w_eco61371, w_eco61372, w_eco61373, w_eco61374, w_eco61375, w_eco61376, w_eco61377, w_eco61378, w_eco61379, w_eco61380, w_eco61381, w_eco61382, w_eco61383, w_eco61384, w_eco61385, w_eco61386, w_eco61387, w_eco61388, w_eco61389, w_eco61390, w_eco61391, w_eco61392, w_eco61393, w_eco61394, w_eco61395, w_eco61396, w_eco61397, w_eco61398, w_eco61399, w_eco61400, w_eco61401, w_eco61402, w_eco61403, w_eco61404, w_eco61405, w_eco61406, w_eco61407, w_eco61408, w_eco61409, w_eco61410, w_eco61411, w_eco61412, w_eco61413, w_eco61414, w_eco61415, w_eco61416, w_eco61417, w_eco61418, w_eco61419, w_eco61420, w_eco61421, w_eco61422, w_eco61423, w_eco61424, w_eco61425, w_eco61426, w_eco61427, w_eco61428, w_eco61429, w_eco61430, w_eco61431, w_eco61432, w_eco61433, w_eco61434, w_eco61435, w_eco61436, w_eco61437, w_eco61438, w_eco61439, w_eco61440, w_eco61441, w_eco61442, w_eco61443, w_eco61444, w_eco61445, w_eco61446, w_eco61447, w_eco61448, w_eco61449, w_eco61450, w_eco61451, w_eco61452, w_eco61453, w_eco61454, w_eco61455, w_eco61456, w_eco61457, w_eco61458, w_eco61459, w_eco61460, w_eco61461, w_eco61462, w_eco61463, w_eco61464, w_eco61465, w_eco61466, w_eco61467, w_eco61468, w_eco61469, w_eco61470, w_eco61471, w_eco61472, w_eco61473, w_eco61474, w_eco61475, w_eco61476, w_eco61477, w_eco61478, w_eco61479, w_eco61480, w_eco61481, w_eco61482, w_eco61483, w_eco61484, w_eco61485, w_eco61486, w_eco61487, w_eco61488, w_eco61489, w_eco61490, w_eco61491, w_eco61492, w_eco61493, w_eco61494, w_eco61495, w_eco61496, w_eco61497, w_eco61498, w_eco61499, w_eco61500, w_eco61501, w_eco61502, w_eco61503, w_eco61504, w_eco61505, w_eco61506, w_eco61507, w_eco61508, w_eco61509, w_eco61510, w_eco61511, w_eco61512, w_eco61513, w_eco61514, w_eco61515, w_eco61516, w_eco61517, w_eco61518, w_eco61519, w_eco61520, w_eco61521, w_eco61522, w_eco61523, w_eco61524, w_eco61525, w_eco61526, w_eco61527, w_eco61528, w_eco61529, w_eco61530, w_eco61531, w_eco61532, w_eco61533, w_eco61534, w_eco61535, w_eco61536, w_eco61537, w_eco61538, w_eco61539, w_eco61540, w_eco61541, w_eco61542, w_eco61543, w_eco61544, w_eco61545, w_eco61546, w_eco61547, w_eco61548, w_eco61549, w_eco61550, w_eco61551, w_eco61552, w_eco61553, w_eco61554, w_eco61555, w_eco61556, w_eco61557, w_eco61558, w_eco61559, w_eco61560, w_eco61561, w_eco61562, w_eco61563, w_eco61564, w_eco61565, w_eco61566, w_eco61567, w_eco61568, w_eco61569, w_eco61570, w_eco61571, w_eco61572, w_eco61573, w_eco61574, w_eco61575, w_eco61576, w_eco61577, w_eco61578, w_eco61579, w_eco61580, w_eco61581, w_eco61582, w_eco61583, w_eco61584, w_eco61585, w_eco61586, w_eco61587, w_eco61588, w_eco61589, w_eco61590, w_eco61591, w_eco61592, w_eco61593, w_eco61594, w_eco61595, w_eco61596, w_eco61597, w_eco61598, w_eco61599, w_eco61600, w_eco61601, w_eco61602, w_eco61603, w_eco61604, w_eco61605, w_eco61606, w_eco61607, w_eco61608, w_eco61609, w_eco61610, w_eco61611, w_eco61612, w_eco61613, w_eco61614, w_eco61615, w_eco61616, w_eco61617, w_eco61618, w_eco61619, w_eco61620, w_eco61621, w_eco61622, w_eco61623, w_eco61624, w_eco61625, w_eco61626, w_eco61627, w_eco61628, w_eco61629, w_eco61630, w_eco61631, w_eco61632, w_eco61633, w_eco61634, w_eco61635, w_eco61636, w_eco61637, w_eco61638, w_eco61639, w_eco61640, w_eco61641, w_eco61642, w_eco61643, w_eco61644, w_eco61645, w_eco61646, w_eco61647, w_eco61648, w_eco61649, w_eco61650, w_eco61651, w_eco61652, w_eco61653, w_eco61654, w_eco61655, w_eco61656, w_eco61657, w_eco61658, w_eco61659, w_eco61660, w_eco61661, w_eco61662, w_eco61663, w_eco61664, w_eco61665, w_eco61666, w_eco61667, w_eco61668, w_eco61669, w_eco61670, w_eco61671, w_eco61672, w_eco61673, w_eco61674, w_eco61675, w_eco61676, w_eco61677, w_eco61678, w_eco61679, w_eco61680, w_eco61681, w_eco61682, w_eco61683, w_eco61684, w_eco61685, w_eco61686, w_eco61687, w_eco61688, w_eco61689, w_eco61690, w_eco61691, w_eco61692, w_eco61693, w_eco61694, w_eco61695, w_eco61696, w_eco61697, w_eco61698, w_eco61699, w_eco61700, w_eco61701, w_eco61702, w_eco61703, w_eco61704, w_eco61705, w_eco61706, w_eco61707, w_eco61708, w_eco61709, w_eco61710, w_eco61711, w_eco61712, w_eco61713, w_eco61714, w_eco61715, w_eco61716, w_eco61717, w_eco61718, w_eco61719, w_eco61720, w_eco61721, w_eco61722, w_eco61723, w_eco61724, w_eco61725, w_eco61726, w_eco61727, w_eco61728, w_eco61729, w_eco61730, w_eco61731, w_eco61732, w_eco61733, w_eco61734, w_eco61735, w_eco61736, w_eco61737, w_eco61738, w_eco61739, w_eco61740, w_eco61741, w_eco61742, w_eco61743, w_eco61744, w_eco61745, w_eco61746, w_eco61747, w_eco61748, w_eco61749, w_eco61750, w_eco61751, w_eco61752, w_eco61753, w_eco61754, w_eco61755, w_eco61756, w_eco61757, w_eco61758, w_eco61759, w_eco61760, w_eco61761, w_eco61762, w_eco61763, w_eco61764, w_eco61765, w_eco61766, w_eco61767, w_eco61768, w_eco61769, w_eco61770, w_eco61771, w_eco61772, w_eco61773, w_eco61774, w_eco61775, w_eco61776, w_eco61777, w_eco61778, w_eco61779, w_eco61780, w_eco61781, w_eco61782, w_eco61783, w_eco61784, w_eco61785, w_eco61786, w_eco61787, w_eco61788, w_eco61789, w_eco61790, w_eco61791, w_eco61792, w_eco61793, w_eco61794, w_eco61795, w_eco61796, w_eco61797, w_eco61798, w_eco61799, w_eco61800, w_eco61801, w_eco61802, w_eco61803, w_eco61804, w_eco61805, w_eco61806, w_eco61807, w_eco61808, w_eco61809, w_eco61810, w_eco61811, w_eco61812, w_eco61813, w_eco61814, w_eco61815, w_eco61816, w_eco61817, w_eco61818, w_eco61819, w_eco61820, w_eco61821, w_eco61822, w_eco61823, w_eco61824, w_eco61825, w_eco61826, w_eco61827, w_eco61828, w_eco61829, w_eco61830, w_eco61831, w_eco61832, w_eco61833, w_eco61834, w_eco61835, w_eco61836, w_eco61837, w_eco61838, w_eco61839, w_eco61840, w_eco61841, w_eco61842, w_eco61843, w_eco61844, w_eco61845, w_eco61846, w_eco61847, w_eco61848, w_eco61849, w_eco61850, w_eco61851, w_eco61852, w_eco61853, w_eco61854, w_eco61855, w_eco61856, w_eco61857, w_eco61858, w_eco61859, w_eco61860, w_eco61861, w_eco61862, w_eco61863, w_eco61864, w_eco61865, w_eco61866, w_eco61867, w_eco61868, w_eco61869, w_eco61870, w_eco61871, w_eco61872, w_eco61873, w_eco61874, w_eco61875, w_eco61876, w_eco61877, w_eco61878, w_eco61879, w_eco61880, w_eco61881, w_eco61882, w_eco61883, w_eco61884, w_eco61885, w_eco61886, w_eco61887, w_eco61888, w_eco61889, w_eco61890, w_eco61891, w_eco61892, w_eco61893, w_eco61894, w_eco61895, w_eco61896, w_eco61897, w_eco61898, w_eco61899, w_eco61900, w_eco61901, w_eco61902, w_eco61903, w_eco61904, w_eco61905, w_eco61906, w_eco61907, w_eco61908, w_eco61909, w_eco61910, w_eco61911, w_eco61912, w_eco61913, w_eco61914, w_eco61915, w_eco61916, w_eco61917, w_eco61918, w_eco61919, w_eco61920, w_eco61921, w_eco61922, w_eco61923, w_eco61924, w_eco61925, w_eco61926, w_eco61927, w_eco61928, w_eco61929, w_eco61930, w_eco61931, w_eco61932, w_eco61933, w_eco61934, w_eco61935, w_eco61936, w_eco61937, w_eco61938, w_eco61939, w_eco61940, w_eco61941, w_eco61942, w_eco61943, w_eco61944, w_eco61945, w_eco61946, w_eco61947, w_eco61948, w_eco61949, w_eco61950, w_eco61951, w_eco61952, w_eco61953, w_eco61954, w_eco61955, w_eco61956, w_eco61957, w_eco61958, w_eco61959, w_eco61960, w_eco61961, w_eco61962, w_eco61963, w_eco61964, w_eco61965, w_eco61966, w_eco61967, w_eco61968, w_eco61969, w_eco61970, w_eco61971, w_eco61972, w_eco61973, w_eco61974, w_eco61975, w_eco61976, w_eco61977, w_eco61978, w_eco61979, w_eco61980, w_eco61981, w_eco61982, w_eco61983, w_eco61984, w_eco61985, w_eco61986, w_eco61987, w_eco61988, w_eco61989, w_eco61990, w_eco61991, w_eco61992, w_eco61993, w_eco61994, w_eco61995, w_eco61996, w_eco61997, w_eco61998, w_eco61999, w_eco62000, w_eco62001, w_eco62002, w_eco62003, w_eco62004, w_eco62005, w_eco62006, w_eco62007, w_eco62008, w_eco62009, w_eco62010, w_eco62011, w_eco62012, w_eco62013, w_eco62014, w_eco62015, w_eco62016, w_eco62017, w_eco62018, w_eco62019, w_eco62020, w_eco62021, w_eco62022, w_eco62023, w_eco62024, w_eco62025, w_eco62026, w_eco62027, w_eco62028, w_eco62029, w_eco62030, w_eco62031, w_eco62032, w_eco62033, w_eco62034, w_eco62035, w_eco62036, w_eco62037, w_eco62038, w_eco62039, w_eco62040, w_eco62041, w_eco62042, w_eco62043, w_eco62044, w_eco62045, w_eco62046, w_eco62047, w_eco62048, w_eco62049, w_eco62050, w_eco62051, w_eco62052, w_eco62053, w_eco62054, w_eco62055, w_eco62056, w_eco62057, w_eco62058, w_eco62059, w_eco62060, w_eco62061, w_eco62062, w_eco62063, w_eco62064, w_eco62065, w_eco62066, w_eco62067, w_eco62068, w_eco62069, w_eco62070, w_eco62071, w_eco62072, w_eco62073, w_eco62074, w_eco62075, w_eco62076, w_eco62077, w_eco62078, w_eco62079, w_eco62080, w_eco62081, w_eco62082, w_eco62083, w_eco62084, w_eco62085, w_eco62086, w_eco62087, w_eco62088, w_eco62089, w_eco62090, w_eco62091, w_eco62092, w_eco62093, w_eco62094, w_eco62095, w_eco62096, w_eco62097, w_eco62098, w_eco62099, w_eco62100, w_eco62101, w_eco62102, w_eco62103, w_eco62104, w_eco62105, w_eco62106, w_eco62107, w_eco62108, w_eco62109, w_eco62110, w_eco62111, w_eco62112, w_eco62113, w_eco62114, w_eco62115, w_eco62116, w_eco62117, w_eco62118, w_eco62119, w_eco62120, w_eco62121, w_eco62122, w_eco62123, w_eco62124, w_eco62125, w_eco62126, w_eco62127, w_eco62128, w_eco62129, w_eco62130, w_eco62131, w_eco62132, w_eco62133, w_eco62134, w_eco62135, w_eco62136, w_eco62137, w_eco62138, w_eco62139, w_eco62140, w_eco62141, w_eco62142, w_eco62143, w_eco62144, w_eco62145, w_eco62146, w_eco62147, w_eco62148, w_eco62149, w_eco62150, w_eco62151, w_eco62152, w_eco62153, w_eco62154, w_eco62155, w_eco62156, w_eco62157, w_eco62158, w_eco62159, w_eco62160, w_eco62161, w_eco62162, w_eco62163, w_eco62164, w_eco62165, w_eco62166, w_eco62167, w_eco62168, w_eco62169, w_eco62170, w_eco62171, w_eco62172, w_eco62173, w_eco62174, w_eco62175, w_eco62176, w_eco62177, w_eco62178, w_eco62179, w_eco62180, w_eco62181, w_eco62182, w_eco62183, w_eco62184, w_eco62185, w_eco62186, w_eco62187, w_eco62188, w_eco62189, w_eco62190, w_eco62191, w_eco62192, w_eco62193, w_eco62194, w_eco62195, w_eco62196, w_eco62197, w_eco62198, w_eco62199, w_eco62200, w_eco62201, w_eco62202, w_eco62203, w_eco62204, w_eco62205, w_eco62206, w_eco62207, w_eco62208, w_eco62209, w_eco62210, w_eco62211, w_eco62212, w_eco62213, w_eco62214, w_eco62215, w_eco62216, w_eco62217, w_eco62218, w_eco62219, w_eco62220, w_eco62221, w_eco62222, w_eco62223, w_eco62224, w_eco62225, w_eco62226, w_eco62227, w_eco62228, w_eco62229, w_eco62230, w_eco62231, w_eco62232, w_eco62233, w_eco62234, w_eco62235, w_eco62236, w_eco62237, w_eco62238, w_eco62239, w_eco62240, w_eco62241, w_eco62242, w_eco62243, w_eco62244, w_eco62245, w_eco62246, w_eco62247, w_eco62248, w_eco62249, w_eco62250, w_eco62251, w_eco62252, w_eco62253, w_eco62254, w_eco62255, w_eco62256, w_eco62257, w_eco62258, w_eco62259, w_eco62260, w_eco62261, w_eco62262, w_eco62263, w_eco62264, w_eco62265, w_eco62266, w_eco62267, w_eco62268, w_eco62269, w_eco62270, w_eco62271, w_eco62272, w_eco62273, w_eco62274, w_eco62275, w_eco62276, w_eco62277, w_eco62278, w_eco62279, w_eco62280, w_eco62281, w_eco62282, w_eco62283, w_eco62284, w_eco62285, w_eco62286, w_eco62287, w_eco62288, w_eco62289, w_eco62290, w_eco62291, w_eco62292, w_eco62293, w_eco62294, w_eco62295, w_eco62296, w_eco62297, w_eco62298, w_eco62299, w_eco62300, w_eco62301, w_eco62302, w_eco62303, w_eco62304, w_eco62305, w_eco62306, w_eco62307, w_eco62308, w_eco62309, w_eco62310, w_eco62311, w_eco62312, w_eco62313, w_eco62314, w_eco62315, w_eco62316, w_eco62317, w_eco62318, w_eco62319, w_eco62320, w_eco62321, w_eco62322, w_eco62323, w_eco62324, w_eco62325, w_eco62326, w_eco62327, w_eco62328, w_eco62329, w_eco62330, w_eco62331, w_eco62332, w_eco62333, w_eco62334, w_eco62335, w_eco62336, w_eco62337, w_eco62338, w_eco62339, w_eco62340, w_eco62341, w_eco62342, w_eco62343, w_eco62344, w_eco62345, w_eco62346, w_eco62347, w_eco62348, w_eco62349, w_eco62350, w_eco62351, w_eco62352, w_eco62353, w_eco62354, w_eco62355, w_eco62356, w_eco62357, w_eco62358, w_eco62359, w_eco62360, w_eco62361, w_eco62362, w_eco62363, w_eco62364, w_eco62365, w_eco62366, w_eco62367, w_eco62368, w_eco62369, w_eco62370, w_eco62371, w_eco62372, w_eco62373, w_eco62374, w_eco62375, w_eco62376, w_eco62377, w_eco62378, w_eco62379, w_eco62380, w_eco62381, w_eco62382, w_eco62383, w_eco62384, w_eco62385, w_eco62386, w_eco62387, w_eco62388, w_eco62389, w_eco62390, w_eco62391, w_eco62392, w_eco62393, w_eco62394, w_eco62395, w_eco62396, w_eco62397, w_eco62398, w_eco62399, w_eco62400, w_eco62401, w_eco62402, w_eco62403, w_eco62404, w_eco62405, w_eco62406, w_eco62407, w_eco62408, w_eco62409, w_eco62410, w_eco62411, w_eco62412, w_eco62413, w_eco62414, w_eco62415, w_eco62416, w_eco62417, w_eco62418, w_eco62419, w_eco62420, w_eco62421, w_eco62422, w_eco62423, w_eco62424, w_eco62425, w_eco62426, w_eco62427, w_eco62428, w_eco62429, w_eco62430, w_eco62431, w_eco62432, w_eco62433, w_eco62434, w_eco62435, w_eco62436, w_eco62437, w_eco62438, w_eco62439, w_eco62440, w_eco62441, w_eco62442, w_eco62443, w_eco62444, w_eco62445, w_eco62446, w_eco62447, w_eco62448, w_eco62449, w_eco62450, w_eco62451, w_eco62452, w_eco62453, w_eco62454, w_eco62455, w_eco62456, w_eco62457, w_eco62458, w_eco62459, w_eco62460, w_eco62461, w_eco62462, w_eco62463, w_eco62464, w_eco62465, w_eco62466, w_eco62467, w_eco62468, w_eco62469, w_eco62470, w_eco62471, w_eco62472, w_eco62473, w_eco62474, w_eco62475, w_eco62476, w_eco62477, w_eco62478, w_eco62479, w_eco62480, w_eco62481, w_eco62482, w_eco62483, w_eco62484, w_eco62485, w_eco62486, w_eco62487, w_eco62488, w_eco62489, w_eco62490, w_eco62491, w_eco62492, w_eco62493, w_eco62494, w_eco62495, w_eco62496, w_eco62497, w_eco62498, w_eco62499, w_eco62500, w_eco62501, w_eco62502, w_eco62503, w_eco62504, w_eco62505, w_eco62506, w_eco62507, w_eco62508, w_eco62509, w_eco62510, w_eco62511, w_eco62512, w_eco62513, w_eco62514, w_eco62515, w_eco62516, w_eco62517, w_eco62518, w_eco62519, w_eco62520, w_eco62521, w_eco62522, w_eco62523, w_eco62524, w_eco62525, w_eco62526, w_eco62527, w_eco62528, w_eco62529, w_eco62530, w_eco62531, w_eco62532, w_eco62533, w_eco62534, w_eco62535, w_eco62536, w_eco62537, w_eco62538, w_eco62539, w_eco62540, w_eco62541, w_eco62542, w_eco62543, w_eco62544, w_eco62545, w_eco62546, w_eco62547, w_eco62548, w_eco62549, w_eco62550, w_eco62551, w_eco62552, w_eco62553, w_eco62554, w_eco62555, w_eco62556, w_eco62557, w_eco62558, w_eco62559, w_eco62560, w_eco62561, w_eco62562, w_eco62563, w_eco62564, w_eco62565, w_eco62566, w_eco62567, w_eco62568, w_eco62569, w_eco62570, w_eco62571, w_eco62572, w_eco62573, w_eco62574, w_eco62575, w_eco62576, w_eco62577, w_eco62578, w_eco62579, w_eco62580, w_eco62581, w_eco62582, w_eco62583, w_eco62584, w_eco62585, w_eco62586, w_eco62587, w_eco62588, w_eco62589, w_eco62590, w_eco62591, w_eco62592, w_eco62593, w_eco62594, w_eco62595, w_eco62596, w_eco62597, w_eco62598, w_eco62599, w_eco62600, w_eco62601, w_eco62602, w_eco62603, w_eco62604, w_eco62605, w_eco62606, w_eco62607, w_eco62608, w_eco62609, w_eco62610, w_eco62611, w_eco62612, w_eco62613, w_eco62614, w_eco62615, w_eco62616, w_eco62617, w_eco62618, w_eco62619, w_eco62620, w_eco62621, w_eco62622, w_eco62623, w_eco62624, w_eco62625, w_eco62626, w_eco62627, w_eco62628, w_eco62629, w_eco62630, w_eco62631, w_eco62632, w_eco62633, w_eco62634, w_eco62635, w_eco62636, w_eco62637, w_eco62638, w_eco62639, w_eco62640, w_eco62641, w_eco62642, w_eco62643, w_eco62644, w_eco62645, w_eco62646, w_eco62647, w_eco62648, w_eco62649, w_eco62650, w_eco62651, w_eco62652, w_eco62653, w_eco62654, w_eco62655, w_eco62656, w_eco62657, w_eco62658, w_eco62659, w_eco62660, w_eco62661, w_eco62662, w_eco62663, w_eco62664, w_eco62665, w_eco62666, w_eco62667, w_eco62668, w_eco62669, w_eco62670, w_eco62671, w_eco62672, w_eco62673, w_eco62674, w_eco62675, w_eco62676, w_eco62677, w_eco62678, w_eco62679, w_eco62680, w_eco62681, w_eco62682, w_eco62683, w_eco62684, w_eco62685, w_eco62686, w_eco62687, w_eco62688, w_eco62689, w_eco62690, w_eco62691, w_eco62692, w_eco62693, w_eco62694, w_eco62695, w_eco62696, w_eco62697, w_eco62698, w_eco62699, w_eco62700, w_eco62701, w_eco62702, w_eco62703, w_eco62704, w_eco62705, w_eco62706, w_eco62707, w_eco62708, w_eco62709, w_eco62710, w_eco62711, w_eco62712, w_eco62713, w_eco62714, w_eco62715, w_eco62716, w_eco62717, w_eco62718, w_eco62719, w_eco62720, w_eco62721, w_eco62722, w_eco62723, w_eco62724, w_eco62725, w_eco62726, w_eco62727, w_eco62728, w_eco62729, w_eco62730, w_eco62731, w_eco62732, w_eco62733, w_eco62734, w_eco62735, w_eco62736, w_eco62737, w_eco62738, w_eco62739, w_eco62740, w_eco62741, w_eco62742, w_eco62743, w_eco62744, w_eco62745, w_eco62746, w_eco62747, w_eco62748, w_eco62749, w_eco62750, w_eco62751, w_eco62752, w_eco62753, w_eco62754, w_eco62755, w_eco62756, w_eco62757, w_eco62758, w_eco62759, w_eco62760, w_eco62761, w_eco62762, w_eco62763, w_eco62764, w_eco62765, w_eco62766, w_eco62767, w_eco62768, w_eco62769, w_eco62770, w_eco62771, w_eco62772, w_eco62773, w_eco62774, w_eco62775, w_eco62776, w_eco62777, w_eco62778, w_eco62779, w_eco62780, w_eco62781, w_eco62782, w_eco62783, w_eco62784, w_eco62785, w_eco62786, w_eco62787, w_eco62788, w_eco62789, w_eco62790, w_eco62791, w_eco62792, w_eco62793, w_eco62794, w_eco62795, w_eco62796, w_eco62797, w_eco62798, w_eco62799, w_eco62800, w_eco62801, w_eco62802, w_eco62803, w_eco62804, w_eco62805, w_eco62806, w_eco62807, w_eco62808, w_eco62809, w_eco62810, w_eco62811, w_eco62812, w_eco62813, w_eco62814, w_eco62815, w_eco62816, w_eco62817, w_eco62818, w_eco62819, w_eco62820, w_eco62821, w_eco62822, w_eco62823, w_eco62824, w_eco62825, w_eco62826, w_eco62827, w_eco62828, w_eco62829, w_eco62830, w_eco62831, w_eco62832, w_eco62833, w_eco62834, w_eco62835, w_eco62836, w_eco62837, w_eco62838, w_eco62839, w_eco62840, w_eco62841, w_eco62842, w_eco62843, w_eco62844, w_eco62845, w_eco62846, w_eco62847, w_eco62848, w_eco62849, w_eco62850, w_eco62851, w_eco62852, w_eco62853, w_eco62854, w_eco62855, w_eco62856, w_eco62857, w_eco62858, w_eco62859, w_eco62860, w_eco62861, w_eco62862, w_eco62863, w_eco62864, w_eco62865, w_eco62866, w_eco62867, w_eco62868, w_eco62869, w_eco62870, w_eco62871, w_eco62872, w_eco62873, w_eco62874, w_eco62875, w_eco62876, w_eco62877, w_eco62878, w_eco62879, w_eco62880, w_eco62881, w_eco62882, w_eco62883, w_eco62884, w_eco62885, w_eco62886, w_eco62887, w_eco62888, w_eco62889, w_eco62890, w_eco62891, w_eco62892, w_eco62893, w_eco62894, w_eco62895, w_eco62896, w_eco62897, w_eco62898, w_eco62899, w_eco62900, w_eco62901, w_eco62902, w_eco62903, w_eco62904, w_eco62905, w_eco62906, w_eco62907, w_eco62908, w_eco62909, w_eco62910, w_eco62911, w_eco62912, w_eco62913, w_eco62914, w_eco62915, w_eco62916, w_eco62917, w_eco62918, w_eco62919, w_eco62920, w_eco62921, w_eco62922, w_eco62923, w_eco62924, w_eco62925, w_eco62926, w_eco62927, w_eco62928, w_eco62929, w_eco62930, w_eco62931, w_eco62932, w_eco62933, w_eco62934, w_eco62935, w_eco62936, w_eco62937, w_eco62938, w_eco62939, w_eco62940, w_eco62941, w_eco62942, w_eco62943, w_eco62944, w_eco62945, w_eco62946, w_eco62947, w_eco62948, w_eco62949, w_eco62950, w_eco62951, w_eco62952, w_eco62953, w_eco62954, w_eco62955, w_eco62956, w_eco62957, w_eco62958, w_eco62959, w_eco62960, w_eco62961, w_eco62962, w_eco62963, w_eco62964, w_eco62965, w_eco62966, w_eco62967, w_eco62968, w_eco62969, w_eco62970, w_eco62971, w_eco62972, w_eco62973, w_eco62974, w_eco62975, w_eco62976, w_eco62977, w_eco62978, w_eco62979, w_eco62980, w_eco62981, w_eco62982, w_eco62983, w_eco62984, w_eco62985, w_eco62986, w_eco62987, w_eco62988, w_eco62989, w_eco62990, w_eco62991, w_eco62992, w_eco62993, w_eco62994, w_eco62995, w_eco62996, w_eco62997, w_eco62998, w_eco62999, w_eco63000, w_eco63001, w_eco63002, w_eco63003, w_eco63004, w_eco63005, w_eco63006, w_eco63007, w_eco63008, w_eco63009, w_eco63010, w_eco63011, w_eco63012, w_eco63013, w_eco63014, w_eco63015, w_eco63016, w_eco63017, w_eco63018, w_eco63019, w_eco63020, w_eco63021, w_eco63022, w_eco63023, w_eco63024, w_eco63025, w_eco63026, w_eco63027, w_eco63028, w_eco63029, w_eco63030, w_eco63031, w_eco63032, w_eco63033, w_eco63034, w_eco63035, w_eco63036, w_eco63037, w_eco63038, w_eco63039, w_eco63040, w_eco63041, w_eco63042, w_eco63043, w_eco63044, w_eco63045, w_eco63046, w_eco63047, w_eco63048, w_eco63049, w_eco63050, w_eco63051, w_eco63052, w_eco63053, w_eco63054, w_eco63055, w_eco63056, w_eco63057, w_eco63058, w_eco63059, w_eco63060, w_eco63061, w_eco63062, w_eco63063, w_eco63064, w_eco63065, w_eco63066, w_eco63067, w_eco63068, w_eco63069, w_eco63070, w_eco63071, w_eco63072, w_eco63073, w_eco63074, w_eco63075, w_eco63076, w_eco63077, w_eco63078, w_eco63079, w_eco63080, w_eco63081, w_eco63082, w_eco63083, w_eco63084, w_eco63085, w_eco63086, w_eco63087, w_eco63088, w_eco63089, w_eco63090, w_eco63091, w_eco63092, w_eco63093, w_eco63094, w_eco63095, w_eco63096, w_eco63097, w_eco63098, w_eco63099, w_eco63100, w_eco63101, w_eco63102, w_eco63103, w_eco63104, w_eco63105, w_eco63106, w_eco63107, w_eco63108, w_eco63109, w_eco63110, w_eco63111, w_eco63112, w_eco63113, w_eco63114, w_eco63115, w_eco63116, w_eco63117, w_eco63118, w_eco63119, w_eco63120, w_eco63121, w_eco63122, w_eco63123, w_eco63124, w_eco63125, w_eco63126, w_eco63127, w_eco63128, w_eco63129, w_eco63130, w_eco63131, w_eco63132, w_eco63133, w_eco63134, w_eco63135, w_eco63136, w_eco63137, w_eco63138, w_eco63139, w_eco63140, w_eco63141, w_eco63142, w_eco63143, w_eco63144, w_eco63145, w_eco63146, w_eco63147, w_eco63148, w_eco63149, w_eco63150, w_eco63151, w_eco63152, w_eco63153, w_eco63154, w_eco63155, w_eco63156, w_eco63157, w_eco63158, w_eco63159, w_eco63160, w_eco63161, w_eco63162, w_eco63163, w_eco63164, w_eco63165, w_eco63166, w_eco63167, w_eco63168, w_eco63169, w_eco63170, w_eco63171, w_eco63172, w_eco63173, w_eco63174, w_eco63175, w_eco63176, w_eco63177, w_eco63178, w_eco63179, w_eco63180, w_eco63181, w_eco63182, w_eco63183, w_eco63184, w_eco63185, w_eco63186, w_eco63187, w_eco63188, w_eco63189, w_eco63190, w_eco63191, w_eco63192, w_eco63193, w_eco63194, w_eco63195, w_eco63196, w_eco63197, w_eco63198, w_eco63199, w_eco63200, w_eco63201, w_eco63202, w_eco63203, w_eco63204, w_eco63205, w_eco63206, w_eco63207, w_eco63208, w_eco63209, w_eco63210, w_eco63211, w_eco63212, w_eco63213, w_eco63214, w_eco63215, w_eco63216, w_eco63217, w_eco63218, w_eco63219, w_eco63220, w_eco63221, w_eco63222, w_eco63223, w_eco63224, w_eco63225, w_eco63226, w_eco63227, w_eco63228, w_eco63229, w_eco63230, w_eco63231, w_eco63232, w_eco63233, w_eco63234, w_eco63235, w_eco63236, w_eco63237, w_eco63238, w_eco63239, w_eco63240, w_eco63241, w_eco63242, w_eco63243, w_eco63244, w_eco63245, w_eco63246, w_eco63247, w_eco63248, w_eco63249, w_eco63250, w_eco63251, w_eco63252, w_eco63253, w_eco63254, w_eco63255, w_eco63256, w_eco63257, w_eco63258, w_eco63259, w_eco63260, w_eco63261, w_eco63262, w_eco63263, w_eco63264, w_eco63265, w_eco63266, w_eco63267, w_eco63268, w_eco63269, w_eco63270, w_eco63271, w_eco63272, w_eco63273, w_eco63274, w_eco63275, w_eco63276, w_eco63277, w_eco63278, w_eco63279, w_eco63280, w_eco63281, w_eco63282, w_eco63283, w_eco63284, w_eco63285, w_eco63286, w_eco63287, w_eco63288, w_eco63289, w_eco63290, w_eco63291, w_eco63292, w_eco63293, w_eco63294, w_eco63295, w_eco63296, w_eco63297, w_eco63298, w_eco63299, w_eco63300, w_eco63301, w_eco63302, w_eco63303, w_eco63304, w_eco63305, w_eco63306, w_eco63307, w_eco63308, w_eco63309, w_eco63310, w_eco63311, w_eco63312, w_eco63313, w_eco63314, w_eco63315, w_eco63316, w_eco63317, w_eco63318, w_eco63319, w_eco63320, w_eco63321, w_eco63322, w_eco63323, w_eco63324, w_eco63325, w_eco63326, w_eco63327, w_eco63328, w_eco63329, w_eco63330, w_eco63331, w_eco63332, w_eco63333, w_eco63334, w_eco63335, w_eco63336, w_eco63337, w_eco63338, w_eco63339, w_eco63340, w_eco63341, w_eco63342, w_eco63343, w_eco63344, w_eco63345, w_eco63346, w_eco63347, w_eco63348, w_eco63349, w_eco63350, w_eco63351, w_eco63352, w_eco63353, w_eco63354, w_eco63355, w_eco63356, w_eco63357, w_eco63358, w_eco63359, w_eco63360, w_eco63361, w_eco63362, w_eco63363, w_eco63364, w_eco63365, w_eco63366, w_eco63367, w_eco63368, w_eco63369, w_eco63370, w_eco63371, w_eco63372, w_eco63373, w_eco63374, w_eco63375, w_eco63376, w_eco63377, w_eco63378, w_eco63379, w_eco63380, w_eco63381, w_eco63382, w_eco63383, w_eco63384, w_eco63385, w_eco63386, w_eco63387, w_eco63388, w_eco63389, w_eco63390, w_eco63391, w_eco63392, w_eco63393, w_eco63394, w_eco63395, w_eco63396, w_eco63397, w_eco63398, w_eco63399, w_eco63400, w_eco63401, w_eco63402, w_eco63403, w_eco63404, w_eco63405, w_eco63406, w_eco63407, w_eco63408, w_eco63409, w_eco63410, w_eco63411, w_eco63412, w_eco63413, w_eco63414, w_eco63415, w_eco63416, w_eco63417, w_eco63418, w_eco63419, w_eco63420, w_eco63421, w_eco63422, w_eco63423, w_eco63424, w_eco63425, w_eco63426, w_eco63427, w_eco63428, w_eco63429, w_eco63430, w_eco63431, w_eco63432, w_eco63433, w_eco63434, w_eco63435, w_eco63436, w_eco63437, w_eco63438, w_eco63439, w_eco63440, w_eco63441, w_eco63442, w_eco63443, w_eco63444, w_eco63445, w_eco63446, w_eco63447, w_eco63448, w_eco63449, w_eco63450, w_eco63451, w_eco63452, w_eco63453, w_eco63454, w_eco63455, w_eco63456, w_eco63457, w_eco63458, w_eco63459, w_eco63460, w_eco63461, w_eco63462, w_eco63463, w_eco63464, w_eco63465, w_eco63466, w_eco63467, w_eco63468, w_eco63469, w_eco63470, w_eco63471, w_eco63472, w_eco63473, w_eco63474, w_eco63475, w_eco63476, w_eco63477, w_eco63478, w_eco63479, w_eco63480, w_eco63481, w_eco63482, w_eco63483, w_eco63484, w_eco63485, w_eco63486, w_eco63487, w_eco63488, w_eco63489, w_eco63490, w_eco63491, w_eco63492, w_eco63493, w_eco63494, w_eco63495, w_eco63496, w_eco63497, w_eco63498, w_eco63499, w_eco63500, w_eco63501, w_eco63502, w_eco63503, w_eco63504, w_eco63505, w_eco63506, w_eco63507, w_eco63508, w_eco63509, w_eco63510, w_eco63511, w_eco63512, w_eco63513, w_eco63514, w_eco63515, w_eco63516, w_eco63517, w_eco63518, w_eco63519, w_eco63520, w_eco63521, w_eco63522, w_eco63523, w_eco63524, w_eco63525, w_eco63526, w_eco63527, w_eco63528, w_eco63529, w_eco63530, w_eco63531, w_eco63532, w_eco63533, w_eco63534, w_eco63535, w_eco63536, w_eco63537, w_eco63538, w_eco63539, w_eco63540, w_eco63541, w_eco63542, w_eco63543, w_eco63544, w_eco63545, w_eco63546, w_eco63547, w_eco63548, w_eco63549, w_eco63550, w_eco63551, w_eco63552, w_eco63553, w_eco63554, w_eco63555, w_eco63556, w_eco63557, w_eco63558, w_eco63559, w_eco63560, w_eco63561, w_eco63562, w_eco63563, w_eco63564, w_eco63565, w_eco63566, w_eco63567, w_eco63568, w_eco63569, w_eco63570, w_eco63571, w_eco63572, w_eco63573, w_eco63574, w_eco63575, w_eco63576, w_eco63577, w_eco63578, w_eco63579, w_eco63580, w_eco63581, w_eco63582, w_eco63583, w_eco63584, w_eco63585, w_eco63586, w_eco63587, w_eco63588, w_eco63589, w_eco63590, w_eco63591, w_eco63592, w_eco63593, w_eco63594, w_eco63595, w_eco63596, w_eco63597, w_eco63598, w_eco63599, w_eco63600, w_eco63601, w_eco63602, w_eco63603, w_eco63604, w_eco63605, w_eco63606, w_eco63607, w_eco63608, w_eco63609, w_eco63610, w_eco63611, w_eco63612, w_eco63613, w_eco63614, w_eco63615, w_eco63616, w_eco63617, w_eco63618, w_eco63619, w_eco63620, w_eco63621, w_eco63622, w_eco63623, w_eco63624, w_eco63625, w_eco63626, w_eco63627, w_eco63628, w_eco63629, w_eco63630, w_eco63631, w_eco63632, w_eco63633, w_eco63634, w_eco63635, w_eco63636, w_eco63637, w_eco63638, w_eco63639, w_eco63640, w_eco63641, w_eco63642, w_eco63643, w_eco63644, w_eco63645, w_eco63646, w_eco63647, w_eco63648, w_eco63649, w_eco63650, w_eco63651, w_eco63652, w_eco63653, w_eco63654, w_eco63655, w_eco63656, w_eco63657, w_eco63658, w_eco63659, w_eco63660, w_eco63661, w_eco63662, w_eco63663, w_eco63664, w_eco63665, w_eco63666, w_eco63667, w_eco63668, w_eco63669, w_eco63670, w_eco63671, w_eco63672, w_eco63673, w_eco63674, w_eco63675, w_eco63676, w_eco63677, w_eco63678, w_eco63679, w_eco63680, w_eco63681, w_eco63682, w_eco63683, w_eco63684, w_eco63685, w_eco63686, w_eco63687, w_eco63688, w_eco63689, w_eco63690, w_eco63691, w_eco63692, w_eco63693, w_eco63694, w_eco63695, w_eco63696, w_eco63697, w_eco63698, w_eco63699, w_eco63700, w_eco63701, w_eco63702, w_eco63703, w_eco63704, w_eco63705, w_eco63706, w_eco63707, w_eco63708, w_eco63709, w_eco63710, w_eco63711, w_eco63712, w_eco63713, w_eco63714, w_eco63715, w_eco63716, w_eco63717, w_eco63718, w_eco63719, w_eco63720, w_eco63721, w_eco63722, w_eco63723, w_eco63724, w_eco63725, w_eco63726, w_eco63727, w_eco63728, w_eco63729, w_eco63730, w_eco63731, w_eco63732, w_eco63733, w_eco63734, w_eco63735, w_eco63736, w_eco63737, w_eco63738, w_eco63739, w_eco63740, w_eco63741, w_eco63742, w_eco63743, w_eco63744, w_eco63745, w_eco63746, w_eco63747, w_eco63748, w_eco63749, w_eco63750, w_eco63751, w_eco63752, w_eco63753, w_eco63754, w_eco63755, w_eco63756, w_eco63757, w_eco63758, w_eco63759, w_eco63760, w_eco63761, w_eco63762, w_eco63763, w_eco63764, w_eco63765, w_eco63766, w_eco63767, w_eco63768, w_eco63769, w_eco63770, w_eco63771, w_eco63772, w_eco63773, w_eco63774, w_eco63775, w_eco63776, w_eco63777, w_eco63778, w_eco63779, w_eco63780, w_eco63781, w_eco63782, w_eco63783, w_eco63784, w_eco63785, w_eco63786, w_eco63787, w_eco63788, w_eco63789, w_eco63790, w_eco63791, w_eco63792, w_eco63793, w_eco63794, w_eco63795, w_eco63796, w_eco63797, w_eco63798, w_eco63799, w_eco63800, w_eco63801, w_eco63802, w_eco63803, w_eco63804, w_eco63805, w_eco63806, w_eco63807, w_eco63808, w_eco63809, w_eco63810, w_eco63811, w_eco63812, w_eco63813, w_eco63814, w_eco63815, w_eco63816, w_eco63817, w_eco63818, w_eco63819, w_eco63820, w_eco63821, w_eco63822, w_eco63823, w_eco63824, w_eco63825, w_eco63826, w_eco63827, w_eco63828, w_eco63829, w_eco63830, w_eco63831, w_eco63832, w_eco63833, w_eco63834, w_eco63835, w_eco63836, w_eco63837, w_eco63838, w_eco63839, w_eco63840, w_eco63841, w_eco63842, w_eco63843, w_eco63844, w_eco63845, w_eco63846, w_eco63847, w_eco63848, w_eco63849, w_eco63850, w_eco63851, w_eco63852, w_eco63853, w_eco63854, w_eco63855, w_eco63856, w_eco63857, w_eco63858, w_eco63859, w_eco63860, w_eco63861, w_eco63862, w_eco63863, w_eco63864, w_eco63865, w_eco63866, w_eco63867, w_eco63868, w_eco63869, w_eco63870, w_eco63871, w_eco63872, w_eco63873, w_eco63874, w_eco63875, w_eco63876, w_eco63877, w_eco63878, w_eco63879, w_eco63880, w_eco63881, w_eco63882, w_eco63883, w_eco63884, w_eco63885, w_eco63886, w_eco63887, w_eco63888, w_eco63889, w_eco63890, w_eco63891, w_eco63892, w_eco63893, w_eco63894, w_eco63895, w_eco63896, w_eco63897, w_eco63898, w_eco63899, w_eco63900, w_eco63901, w_eco63902, w_eco63903, w_eco63904, w_eco63905, w_eco63906, w_eco63907, w_eco63908, w_eco63909, w_eco63910, w_eco63911, w_eco63912, w_eco63913, w_eco63914, w_eco63915, w_eco63916, w_eco63917, w_eco63918, w_eco63919, w_eco63920, w_eco63921, w_eco63922, w_eco63923, w_eco63924, w_eco63925, w_eco63926, w_eco63927, w_eco63928, w_eco63929, w_eco63930, w_eco63931, w_eco63932, w_eco63933, w_eco63934, w_eco63935, w_eco63936, w_eco63937, w_eco63938, w_eco63939, w_eco63940, w_eco63941, w_eco63942, w_eco63943, w_eco63944, w_eco63945, w_eco63946, w_eco63947, w_eco63948, w_eco63949, w_eco63950, w_eco63951, w_eco63952, w_eco63953, w_eco63954, w_eco63955, w_eco63956, w_eco63957, w_eco63958, w_eco63959, w_eco63960, w_eco63961, w_eco63962, w_eco63963, w_eco63964, w_eco63965, w_eco63966, w_eco63967, w_eco63968, w_eco63969, w_eco63970, w_eco63971, w_eco63972, w_eco63973, w_eco63974, w_eco63975, w_eco63976, w_eco63977, w_eco63978, w_eco63979, w_eco63980, w_eco63981, w_eco63982, w_eco63983, w_eco63984, w_eco63985, w_eco63986, w_eco63987, w_eco63988, w_eco63989, w_eco63990, w_eco63991, w_eco63992, w_eco63993, w_eco63994, w_eco63995, w_eco63996, w_eco63997, w_eco63998, w_eco63999, w_eco64000, w_eco64001, w_eco64002, w_eco64003, w_eco64004, w_eco64005, w_eco64006, w_eco64007, w_eco64008, w_eco64009, w_eco64010, w_eco64011, w_eco64012, w_eco64013, w_eco64014, w_eco64015, w_eco64016, w_eco64017, w_eco64018, w_eco64019, w_eco64020, w_eco64021, w_eco64022, w_eco64023, w_eco64024, w_eco64025, w_eco64026, w_eco64027, w_eco64028, w_eco64029, w_eco64030, w_eco64031, w_eco64032, w_eco64033, w_eco64034, w_eco64035, w_eco64036, w_eco64037, w_eco64038, w_eco64039, w_eco64040, w_eco64041, w_eco64042, w_eco64043, w_eco64044, w_eco64045, w_eco64046, w_eco64047, w_eco64048, w_eco64049, w_eco64050, w_eco64051, w_eco64052, w_eco64053, w_eco64054, w_eco64055, w_eco64056, w_eco64057, w_eco64058, w_eco64059, w_eco64060, w_eco64061, w_eco64062, w_eco64063, w_eco64064, w_eco64065, w_eco64066, w_eco64067, w_eco64068, w_eco64069, w_eco64070, w_eco64071, w_eco64072, w_eco64073, w_eco64074, w_eco64075, w_eco64076, w_eco64077, w_eco64078, w_eco64079, w_eco64080, w_eco64081, w_eco64082, w_eco64083, w_eco64084, w_eco64085, w_eco64086, w_eco64087, w_eco64088, w_eco64089, w_eco64090, w_eco64091, w_eco64092, w_eco64093, w_eco64094, w_eco64095, w_eco64096, w_eco64097, w_eco64098, w_eco64099, w_eco64100, w_eco64101, w_eco64102, w_eco64103, w_eco64104, w_eco64105, w_eco64106, w_eco64107, w_eco64108, w_eco64109, w_eco64110, w_eco64111, w_eco64112, w_eco64113, w_eco64114, w_eco64115, w_eco64116, w_eco64117, w_eco64118, w_eco64119, w_eco64120, w_eco64121, w_eco64122, w_eco64123, w_eco64124, w_eco64125, w_eco64126, w_eco64127, w_eco64128, w_eco64129, w_eco64130, w_eco64131, w_eco64132, w_eco64133, w_eco64134, w_eco64135, w_eco64136, w_eco64137, w_eco64138, w_eco64139, w_eco64140, w_eco64141, w_eco64142, w_eco64143, w_eco64144, w_eco64145, w_eco64146, w_eco64147, w_eco64148, w_eco64149, w_eco64150, w_eco64151, w_eco64152, w_eco64153, w_eco64154, w_eco64155, w_eco64156, w_eco64157, w_eco64158, w_eco64159, w_eco64160, w_eco64161, w_eco64162, w_eco64163, w_eco64164, w_eco64165, w_eco64166, w_eco64167, w_eco64168, w_eco64169, w_eco64170, w_eco64171, w_eco64172, w_eco64173, w_eco64174, w_eco64175, w_eco64176, w_eco64177, w_eco64178, w_eco64179, w_eco64180, w_eco64181, w_eco64182, w_eco64183, w_eco64184, w_eco64185, w_eco64186, w_eco64187, w_eco64188, w_eco64189, w_eco64190, w_eco64191, w_eco64192, w_eco64193, w_eco64194, w_eco64195, w_eco64196, w_eco64197, w_eco64198, w_eco64199, w_eco64200, w_eco64201, w_eco64202, w_eco64203, w_eco64204, w_eco64205, w_eco64206, w_eco64207, w_eco64208, w_eco64209, w_eco64210, w_eco64211, w_eco64212, w_eco64213, w_eco64214, w_eco64215, w_eco64216, w_eco64217, w_eco64218, w_eco64219, w_eco64220, w_eco64221, w_eco64222, w_eco64223, w_eco64224, w_eco64225, w_eco64226, w_eco64227, w_eco64228, w_eco64229, w_eco64230, w_eco64231, w_eco64232, w_eco64233, w_eco64234, w_eco64235, w_eco64236, w_eco64237, w_eco64238, w_eco64239, w_eco64240, w_eco64241, w_eco64242, w_eco64243, w_eco64244, w_eco64245, w_eco64246, w_eco64247, w_eco64248, w_eco64249, w_eco64250, w_eco64251, w_eco64252, w_eco64253, w_eco64254, w_eco64255, w_eco64256, w_eco64257, w_eco64258, w_eco64259, w_eco64260, w_eco64261, w_eco64262, w_eco64263, w_eco64264, w_eco64265, w_eco64266, w_eco64267, w_eco64268, w_eco64269, w_eco64270, w_eco64271, w_eco64272, w_eco64273, w_eco64274, w_eco64275, w_eco64276, w_eco64277, w_eco64278, w_eco64279, w_eco64280, w_eco64281, w_eco64282, w_eco64283, w_eco64284, w_eco64285, w_eco64286, w_eco64287, w_eco64288, w_eco64289, w_eco64290, w_eco64291, w_eco64292, w_eco64293, w_eco64294, w_eco64295, w_eco64296, w_eco64297, w_eco64298, w_eco64299, w_eco64300, w_eco64301, w_eco64302, w_eco64303, w_eco64304, w_eco64305, w_eco64306, w_eco64307, w_eco64308, w_eco64309, w_eco64310, w_eco64311, w_eco64312, w_eco64313, w_eco64314, w_eco64315, w_eco64316, w_eco64317, w_eco64318, w_eco64319, w_eco64320, w_eco64321, w_eco64322, w_eco64323, w_eco64324, w_eco64325, w_eco64326, w_eco64327, w_eco64328, w_eco64329, w_eco64330, w_eco64331, w_eco64332, w_eco64333, w_eco64334, w_eco64335, w_eco64336, w_eco64337, w_eco64338, w_eco64339, w_eco64340, w_eco64341, w_eco64342, w_eco64343, w_eco64344, w_eco64345, w_eco64346, w_eco64347, w_eco64348, w_eco64349, w_eco64350, w_eco64351, w_eco64352, w_eco64353, w_eco64354, w_eco64355, w_eco64356, w_eco64357, w_eco64358, w_eco64359, w_eco64360, w_eco64361, w_eco64362, w_eco64363, w_eco64364, w_eco64365, w_eco64366, w_eco64367, w_eco64368, w_eco64369, w_eco64370, w_eco64371, w_eco64372, w_eco64373, w_eco64374, w_eco64375, w_eco64376, w_eco64377, w_eco64378, w_eco64379, w_eco64380, w_eco64381, w_eco64382, w_eco64383, w_eco64384, w_eco64385, w_eco64386, w_eco64387, w_eco64388, w_eco64389, w_eco64390, w_eco64391, w_eco64392, w_eco64393, w_eco64394, w_eco64395, w_eco64396, w_eco64397, w_eco64398, w_eco64399, w_eco64400, w_eco64401, w_eco64402, w_eco64403, w_eco64404, w_eco64405, w_eco64406, w_eco64407, w_eco64408, w_eco64409, w_eco64410, w_eco64411, w_eco64412, w_eco64413, w_eco64414, w_eco64415, w_eco64416, w_eco64417, w_eco64418, w_eco64419, w_eco64420, w_eco64421, w_eco64422, w_eco64423, w_eco64424, w_eco64425, w_eco64426, w_eco64427, w_eco64428, w_eco64429, w_eco64430, w_eco64431, w_eco64432, w_eco64433, w_eco64434, w_eco64435, w_eco64436, w_eco64437, w_eco64438, w_eco64439, w_eco64440, w_eco64441, w_eco64442, w_eco64443, w_eco64444, w_eco64445, w_eco64446, w_eco64447, w_eco64448, w_eco64449, w_eco64450, w_eco64451, w_eco64452, w_eco64453, w_eco64454, w_eco64455, w_eco64456, w_eco64457, w_eco64458, w_eco64459, w_eco64460, w_eco64461, w_eco64462, w_eco64463, w_eco64464, w_eco64465, w_eco64466, w_eco64467, w_eco64468, w_eco64469, w_eco64470, w_eco64471, w_eco64472, w_eco64473, w_eco64474, w_eco64475, w_eco64476, w_eco64477, w_eco64478, w_eco64479, w_eco64480, w_eco64481, w_eco64482, w_eco64483, w_eco64484, w_eco64485, w_eco64486, w_eco64487, w_eco64488, w_eco64489, w_eco64490, w_eco64491, w_eco64492, w_eco64493, w_eco64494, w_eco64495, w_eco64496, w_eco64497, w_eco64498, w_eco64499, w_eco64500, w_eco64501, w_eco64502, w_eco64503, w_eco64504, w_eco64505, w_eco64506, w_eco64507, w_eco64508, w_eco64509, w_eco64510, w_eco64511, w_eco64512, w_eco64513, w_eco64514, w_eco64515, w_eco64516, w_eco64517, w_eco64518, w_eco64519, w_eco64520, w_eco64521, w_eco64522, w_eco64523, w_eco64524, w_eco64525, w_eco64526, w_eco64527, w_eco64528, w_eco64529, w_eco64530, w_eco64531, w_eco64532, w_eco64533, w_eco64534, w_eco64535, w_eco64536, w_eco64537, w_eco64538, w_eco64539, w_eco64540, w_eco64541, w_eco64542, w_eco64543, w_eco64544, w_eco64545, w_eco64546, w_eco64547, w_eco64548, w_eco64549, w_eco64550, w_eco64551, w_eco64552, w_eco64553, w_eco64554, w_eco64555, w_eco64556, w_eco64557, w_eco64558, w_eco64559, w_eco64560, w_eco64561, w_eco64562, w_eco64563, w_eco64564, w_eco64565, w_eco64566, w_eco64567, w_eco64568, w_eco64569, w_eco64570, w_eco64571, w_eco64572, w_eco64573, w_eco64574, w_eco64575, w_eco64576, w_eco64577, w_eco64578, w_eco64579, w_eco64580, w_eco64581, w_eco64582, w_eco64583, w_eco64584, w_eco64585, w_eco64586, w_eco64587, w_eco64588, w_eco64589, w_eco64590, w_eco64591, w_eco64592, w_eco64593, w_eco64594, w_eco64595, w_eco64596, w_eco64597, w_eco64598, w_eco64599, w_eco64600, w_eco64601, w_eco64602, w_eco64603, w_eco64604, w_eco64605, w_eco64606, w_eco64607, w_eco64608, w_eco64609, w_eco64610, w_eco64611, w_eco64612, w_eco64613, w_eco64614, w_eco64615, w_eco64616, w_eco64617, w_eco64618, w_eco64619, w_eco64620, w_eco64621, w_eco64622, w_eco64623, w_eco64624, w_eco64625, w_eco64626, w_eco64627, w_eco64628, w_eco64629, w_eco64630, w_eco64631, w_eco64632, w_eco64633, w_eco64634, w_eco64635, w_eco64636, w_eco64637, w_eco64638, w_eco64639, w_eco64640, w_eco64641, w_eco64642, w_eco64643, w_eco64644, w_eco64645, w_eco64646, w_eco64647, w_eco64648, w_eco64649, w_eco64650, w_eco64651, w_eco64652, w_eco64653, w_eco64654, w_eco64655, w_eco64656, w_eco64657, w_eco64658, w_eco64659, w_eco64660, w_eco64661, w_eco64662, w_eco64663, w_eco64664, w_eco64665, w_eco64666, w_eco64667, w_eco64668, w_eco64669, w_eco64670, w_eco64671, w_eco64672, w_eco64673, w_eco64674, w_eco64675, w_eco64676, w_eco64677, w_eco64678, w_eco64679, w_eco64680, w_eco64681, w_eco64682, w_eco64683, w_eco64684, w_eco64685, w_eco64686, w_eco64687, w_eco64688, w_eco64689, w_eco64690, w_eco64691, w_eco64692, w_eco64693, w_eco64694, w_eco64695, w_eco64696, w_eco64697, w_eco64698, w_eco64699, w_eco64700, w_eco64701, w_eco64702, w_eco64703, w_eco64704, w_eco64705, w_eco64706, w_eco64707, w_eco64708, w_eco64709, w_eco64710, w_eco64711, w_eco64712, w_eco64713, w_eco64714, w_eco64715, w_eco64716, w_eco64717, w_eco64718, w_eco64719, w_eco64720, w_eco64721, w_eco64722, w_eco64723, w_eco64724, w_eco64725, w_eco64726, w_eco64727, w_eco64728, w_eco64729, w_eco64730, w_eco64731, w_eco64732, w_eco64733, w_eco64734, w_eco64735, w_eco64736, w_eco64737, w_eco64738, w_eco64739, w_eco64740, w_eco64741, w_eco64742, w_eco64743, w_eco64744, w_eco64745, w_eco64746, w_eco64747, w_eco64748, w_eco64749, w_eco64750, w_eco64751, w_eco64752, w_eco64753, w_eco64754, w_eco64755, w_eco64756, w_eco64757, w_eco64758, w_eco64759, w_eco64760, w_eco64761, w_eco64762, w_eco64763, w_eco64764, w_eco64765, w_eco64766, w_eco64767, w_eco64768, w_eco64769, w_eco64770, w_eco64771, w_eco64772, w_eco64773, w_eco64774, w_eco64775, w_eco64776, w_eco64777, w_eco64778, w_eco64779, w_eco64780, w_eco64781, w_eco64782, w_eco64783, w_eco64784, w_eco64785, w_eco64786, w_eco64787, w_eco64788, w_eco64789, w_eco64790, w_eco64791, w_eco64792, w_eco64793, w_eco64794, w_eco64795, w_eco64796, w_eco64797, w_eco64798, w_eco64799, w_eco64800, w_eco64801, w_eco64802, w_eco64803, w_eco64804, w_eco64805, w_eco64806, w_eco64807, w_eco64808, w_eco64809, w_eco64810, w_eco64811, w_eco64812, w_eco64813, w_eco64814, w_eco64815, w_eco64816, w_eco64817, w_eco64818, w_eco64819, w_eco64820, w_eco64821, w_eco64822, w_eco64823, w_eco64824, w_eco64825, w_eco64826, w_eco64827, w_eco64828, w_eco64829, w_eco64830, w_eco64831, w_eco64832, w_eco64833, w_eco64834, w_eco64835, w_eco64836, w_eco64837, w_eco64838, w_eco64839, w_eco64840, w_eco64841, w_eco64842, w_eco64843, w_eco64844, w_eco64845, w_eco64846, w_eco64847, w_eco64848, w_eco64849, w_eco64850, w_eco64851, w_eco64852, w_eco64853, w_eco64854, w_eco64855, w_eco64856, w_eco64857, w_eco64858, w_eco64859, w_eco64860, w_eco64861, w_eco64862, w_eco64863, w_eco64864, w_eco64865, w_eco64866, w_eco64867, w_eco64868, w_eco64869, w_eco64870, w_eco64871, w_eco64872, w_eco64873, w_eco64874, w_eco64875, w_eco64876, w_eco64877, w_eco64878, w_eco64879, w_eco64880, w_eco64881, w_eco64882, w_eco64883, w_eco64884, w_eco64885, w_eco64886, w_eco64887, w_eco64888, w_eco64889, w_eco64890, w_eco64891, w_eco64892, w_eco64893, w_eco64894, w_eco64895, w_eco64896, w_eco64897, w_eco64898, w_eco64899, w_eco64900, w_eco64901, w_eco64902, w_eco64903, w_eco64904, w_eco64905, w_eco64906, w_eco64907, w_eco64908, w_eco64909, w_eco64910, w_eco64911, w_eco64912, w_eco64913, w_eco64914, w_eco64915, w_eco64916, w_eco64917, w_eco64918, w_eco64919, w_eco64920, w_eco64921, w_eco64922, w_eco64923, w_eco64924, w_eco64925, w_eco64926, w_eco64927, w_eco64928, w_eco64929, w_eco64930, w_eco64931, w_eco64932, w_eco64933, w_eco64934, w_eco64935, w_eco64936, w_eco64937, w_eco64938, w_eco64939, w_eco64940, w_eco64941, w_eco64942, w_eco64943, w_eco64944, w_eco64945, w_eco64946, w_eco64947, w_eco64948, w_eco64949, w_eco64950, w_eco64951, w_eco64952, w_eco64953, w_eco64954, w_eco64955, w_eco64956, w_eco64957, w_eco64958, w_eco64959, w_eco64960, w_eco64961, w_eco64962, w_eco64963, w_eco64964, w_eco64965, w_eco64966, w_eco64967, w_eco64968, w_eco64969, w_eco64970, w_eco64971, w_eco64972, w_eco64973, w_eco64974, w_eco64975, w_eco64976, w_eco64977, w_eco64978, w_eco64979, w_eco64980, w_eco64981, w_eco64982, w_eco64983, w_eco64984, w_eco64985, w_eco64986, w_eco64987, w_eco64988, w_eco64989, w_eco64990, w_eco64991, w_eco64992, w_eco64993, w_eco64994, w_eco64995, w_eco64996, w_eco64997, w_eco64998, w_eco64999, w_eco65000, w_eco65001, w_eco65002, w_eco65003, w_eco65004, w_eco65005, w_eco65006, w_eco65007, w_eco65008, w_eco65009, w_eco65010, w_eco65011, w_eco65012, w_eco65013, w_eco65014, w_eco65015, w_eco65016, w_eco65017, w_eco65018, w_eco65019, w_eco65020, w_eco65021, w_eco65022, w_eco65023, w_eco65024, w_eco65025, w_eco65026, w_eco65027, w_eco65028, w_eco65029, w_eco65030, w_eco65031, w_eco65032, w_eco65033, w_eco65034, w_eco65035, w_eco65036, w_eco65037, w_eco65038, w_eco65039, w_eco65040, w_eco65041, w_eco65042, w_eco65043, w_eco65044, w_eco65045, w_eco65046, w_eco65047, w_eco65048, w_eco65049, w_eco65050, w_eco65051, w_eco65052, w_eco65053, w_eco65054, w_eco65055, w_eco65056, w_eco65057, w_eco65058, w_eco65059, w_eco65060, w_eco65061, w_eco65062, w_eco65063, w_eco65064, w_eco65065, w_eco65066, w_eco65067, w_eco65068, w_eco65069, w_eco65070, w_eco65071, w_eco65072, w_eco65073, w_eco65074, w_eco65075, w_eco65076, w_eco65077, w_eco65078, w_eco65079, w_eco65080, w_eco65081, w_eco65082, w_eco65083, w_eco65084, w_eco65085, w_eco65086, w_eco65087, w_eco65088, w_eco65089, w_eco65090, w_eco65091, w_eco65092, w_eco65093, w_eco65094, w_eco65095, w_eco65096, w_eco65097, w_eco65098, w_eco65099, w_eco65100, w_eco65101, w_eco65102, w_eco65103, w_eco65104, w_eco65105, w_eco65106, w_eco65107, w_eco65108, w_eco65109, w_eco65110, w_eco65111, w_eco65112, w_eco65113, w_eco65114, w_eco65115, w_eco65116, w_eco65117, w_eco65118, w_eco65119, w_eco65120, w_eco65121, w_eco65122, w_eco65123, w_eco65124, w_eco65125, w_eco65126, w_eco65127, w_eco65128, w_eco65129, w_eco65130, w_eco65131, w_eco65132, w_eco65133, w_eco65134, w_eco65135, w_eco65136, w_eco65137, w_eco65138, w_eco65139, w_eco65140, w_eco65141, w_eco65142, w_eco65143, w_eco65144, w_eco65145, w_eco65146, w_eco65147, w_eco65148, w_eco65149, w_eco65150, w_eco65151, w_eco65152, w_eco65153, w_eco65154, w_eco65155, w_eco65156, w_eco65157, w_eco65158, w_eco65159, w_eco65160, w_eco65161, w_eco65162, w_eco65163, w_eco65164, w_eco65165, w_eco65166, w_eco65167, w_eco65168, w_eco65169, w_eco65170, w_eco65171, w_eco65172, w_eco65173, w_eco65174, w_eco65175, w_eco65176, w_eco65177, w_eco65178, w_eco65179, w_eco65180, w_eco65181, w_eco65182, w_eco65183, w_eco65184, w_eco65185, w_eco65186, w_eco65187, w_eco65188, w_eco65189, w_eco65190, w_eco65191, w_eco65192, w_eco65193, w_eco65194, w_eco65195, w_eco65196, w_eco65197, w_eco65198, w_eco65199, w_eco65200, w_eco65201, w_eco65202, w_eco65203, w_eco65204, w_eco65205, w_eco65206, w_eco65207, w_eco65208, w_eco65209, w_eco65210, w_eco65211, w_eco65212, w_eco65213, w_eco65214, w_eco65215, w_eco65216, w_eco65217, w_eco65218, w_eco65219, w_eco65220, w_eco65221, w_eco65222, w_eco65223, w_eco65224, w_eco65225, w_eco65226, w_eco65227, w_eco65228, w_eco65229, w_eco65230, w_eco65231, w_eco65232, w_eco65233, w_eco65234, w_eco65235, w_eco65236, w_eco65237, w_eco65238, w_eco65239, w_eco65240, w_eco65241, w_eco65242, w_eco65243, w_eco65244, w_eco65245, w_eco65246, w_eco65247, w_eco65248, w_eco65249, w_eco65250, w_eco65251, w_eco65252, w_eco65253, w_eco65254, w_eco65255, w_eco65256, w_eco65257, w_eco65258, w_eco65259, w_eco65260, w_eco65261, w_eco65262, w_eco65263, w_eco65264, w_eco65265, w_eco65266, w_eco65267, w_eco65268, w_eco65269, w_eco65270, w_eco65271, w_eco65272, w_eco65273, w_eco65274, w_eco65275, w_eco65276, w_eco65277, w_eco65278, w_eco65279, w_eco65280, w_eco65281, w_eco65282, w_eco65283, w_eco65284, w_eco65285, w_eco65286, w_eco65287, w_eco65288, w_eco65289, w_eco65290, w_eco65291, w_eco65292, w_eco65293, w_eco65294, w_eco65295, w_eco65296, w_eco65297, w_eco65298, w_eco65299, w_eco65300, w_eco65301, w_eco65302, w_eco65303, w_eco65304, w_eco65305, w_eco65306, w_eco65307, w_eco65308, w_eco65309, w_eco65310, w_eco65311, w_eco65312, w_eco65313, w_eco65314, w_eco65315, w_eco65316, w_eco65317, w_eco65318, w_eco65319, w_eco65320, w_eco65321, w_eco65322, w_eco65323, w_eco65324, w_eco65325, w_eco65326, w_eco65327, w_eco65328, w_eco65329, w_eco65330, w_eco65331, w_eco65332, w_eco65333, w_eco65334, w_eco65335, w_eco65336, w_eco65337, w_eco65338, w_eco65339, w_eco65340, w_eco65341, w_eco65342, w_eco65343, w_eco65344, w_eco65345, w_eco65346, w_eco65347, w_eco65348, w_eco65349, w_eco65350, w_eco65351, w_eco65352, w_eco65353, w_eco65354, w_eco65355, w_eco65356, w_eco65357, w_eco65358, w_eco65359, w_eco65360, w_eco65361, w_eco65362, w_eco65363, w_eco65364, w_eco65365, w_eco65366, w_eco65367, w_eco65368, w_eco65369, w_eco65370, w_eco65371, w_eco65372, w_eco65373, w_eco65374, w_eco65375, w_eco65376, w_eco65377, w_eco65378, w_eco65379, w_eco65380, w_eco65381, w_eco65382, w_eco65383, w_eco65384, w_eco65385, w_eco65386, w_eco65387, w_eco65388, w_eco65389, w_eco65390, w_eco65391, w_eco65392, w_eco65393, w_eco65394, w_eco65395, w_eco65396, w_eco65397, w_eco65398, w_eco65399, w_eco65400, w_eco65401, w_eco65402, w_eco65403, w_eco65404, w_eco65405, w_eco65406, w_eco65407, w_eco65408, w_eco65409, w_eco65410, w_eco65411, w_eco65412, w_eco65413, w_eco65414, w_eco65415, w_eco65416, w_eco65417, w_eco65418, w_eco65419, w_eco65420, w_eco65421, w_eco65422, w_eco65423, w_eco65424, w_eco65425, w_eco65426, w_eco65427, w_eco65428, w_eco65429, w_eco65430, w_eco65431, w_eco65432, w_eco65433, w_eco65434, w_eco65435, w_eco65436, w_eco65437, w_eco65438, w_eco65439, w_eco65440, w_eco65441, w_eco65442, w_eco65443, w_eco65444, w_eco65445, w_eco65446, w_eco65447, w_eco65448, w_eco65449, w_eco65450, w_eco65451, w_eco65452, w_eco65453, w_eco65454, w_eco65455, w_eco65456, w_eco65457, w_eco65458, w_eco65459, w_eco65460, w_eco65461, w_eco65462, w_eco65463, w_eco65464, w_eco65465, w_eco65466, w_eco65467, w_eco65468, w_eco65469, w_eco65470, w_eco65471, w_eco65472, w_eco65473, w_eco65474, w_eco65475, w_eco65476, w_eco65477, w_eco65478, w_eco65479, w_eco65480, w_eco65481, w_eco65482, w_eco65483, w_eco65484, w_eco65485, w_eco65486, w_eco65487, w_eco65488, w_eco65489, w_eco65490, w_eco65491, w_eco65492, w_eco65493, w_eco65494, w_eco65495, w_eco65496, w_eco65497, w_eco65498, w_eco65499, w_eco65500, w_eco65501, w_eco65502, w_eco65503, w_eco65504, w_eco65505, w_eco65506, w_eco65507, w_eco65508, w_eco65509, w_eco65510, w_eco65511, w_eco65512, w_eco65513, w_eco65514, w_eco65515, w_eco65516, w_eco65517, w_eco65518, w_eco65519, w_eco65520, w_eco65521, w_eco65522, w_eco65523, w_eco65524, w_eco65525, w_eco65526, w_eco65527, w_eco65528, w_eco65529, w_eco65530, w_eco65531, w_eco65532, w_eco65533, w_eco65534, w_eco65535, w_eco65536, w_eco65537, w_eco65538, w_eco65539, w_eco65540, w_eco65541, w_eco65542, w_eco65543, w_eco65544, w_eco65545, w_eco65546, w_eco65547, w_eco65548, w_eco65549, w_eco65550, w_eco65551, w_eco65552, w_eco65553, w_eco65554, w_eco65555, w_eco65556, w_eco65557, w_eco65558, w_eco65559, w_eco65560, w_eco65561, w_eco65562, w_eco65563, w_eco65564, w_eco65565, w_eco65566, w_eco65567, w_eco65568, w_eco65569, w_eco65570, w_eco65571, w_eco65572, w_eco65573, w_eco65574, w_eco65575, w_eco65576, w_eco65577, w_eco65578, w_eco65579, w_eco65580, w_eco65581, w_eco65582, w_eco65583, w_eco65584, w_eco65585, w_eco65586, w_eco65587, w_eco65588, w_eco65589, w_eco65590, w_eco65591, w_eco65592, w_eco65593, w_eco65594, w_eco65595, w_eco65596, w_eco65597, w_eco65598, w_eco65599, w_eco65600, w_eco65601, w_eco65602, w_eco65603, w_eco65604, w_eco65605, w_eco65606, w_eco65607, w_eco65608, w_eco65609, w_eco65610, w_eco65611, w_eco65612, w_eco65613, w_eco65614, w_eco65615, w_eco65616, w_eco65617, w_eco65618, w_eco65619, w_eco65620, w_eco65621, w_eco65622, w_eco65623, w_eco65624, w_eco65625, w_eco65626, w_eco65627, w_eco65628, w_eco65629, w_eco65630, w_eco65631, w_eco65632, w_eco65633, w_eco65634, w_eco65635, w_eco65636, w_eco65637, w_eco65638, w_eco65639, w_eco65640, w_eco65641, w_eco65642, w_eco65643, w_eco65644, w_eco65645, w_eco65646, w_eco65647, w_eco65648, w_eco65649, w_eco65650, w_eco65651, w_eco65652, w_eco65653, w_eco65654, w_eco65655, w_eco65656, w_eco65657, w_eco65658, w_eco65659, w_eco65660, w_eco65661, w_eco65662, w_eco65663, w_eco65664, w_eco65665, w_eco65666, w_eco65667, w_eco65668, w_eco65669, w_eco65670, w_eco65671, w_eco65672, w_eco65673, w_eco65674, w_eco65675, w_eco65676, w_eco65677, w_eco65678, w_eco65679, w_eco65680, w_eco65681, w_eco65682, w_eco65683, w_eco65684, w_eco65685, w_eco65686, w_eco65687, w_eco65688, w_eco65689, w_eco65690, w_eco65691, w_eco65692, w_eco65693, w_eco65694, w_eco65695, w_eco65696, w_eco65697, w_eco65698, w_eco65699, w_eco65700, w_eco65701, w_eco65702, w_eco65703, w_eco65704, w_eco65705, w_eco65706, w_eco65707, w_eco65708, w_eco65709, w_eco65710, w_eco65711, w_eco65712, w_eco65713, w_eco65714, w_eco65715, w_eco65716, w_eco65717, w_eco65718, w_eco65719, w_eco65720, w_eco65721, w_eco65722, w_eco65723, w_eco65724, w_eco65725, w_eco65726, w_eco65727, w_eco65728, w_eco65729, w_eco65730, w_eco65731, w_eco65732, w_eco65733, w_eco65734, w_eco65735, w_eco65736, w_eco65737, w_eco65738, w_eco65739, w_eco65740, w_eco65741, w_eco65742, w_eco65743, w_eco65744, w_eco65745, w_eco65746, w_eco65747, w_eco65748, w_eco65749, w_eco65750, w_eco65751, w_eco65752, w_eco65753, w_eco65754, w_eco65755, w_eco65756, w_eco65757, w_eco65758, w_eco65759, w_eco65760, w_eco65761, w_eco65762, w_eco65763, w_eco65764, w_eco65765, w_eco65766, w_eco65767, w_eco65768, w_eco65769, w_eco65770, w_eco65771, w_eco65772, w_eco65773, w_eco65774, w_eco65775, w_eco65776, w_eco65777, w_eco65778, w_eco65779, w_eco65780, w_eco65781, w_eco65782, w_eco65783, w_eco65784, w_eco65785, w_eco65786, w_eco65787, w_eco65788, w_eco65789, w_eco65790, w_eco65791, w_eco65792, w_eco65793, w_eco65794, w_eco65795, w_eco65796, w_eco65797, w_eco65798, w_eco65799, w_eco65800, w_eco65801, w_eco65802, w_eco65803, w_eco65804, w_eco65805, w_eco65806, w_eco65807, w_eco65808, w_eco65809, w_eco65810, w_eco65811, w_eco65812, w_eco65813, w_eco65814, w_eco65815, w_eco65816, w_eco65817, w_eco65818, w_eco65819, w_eco65820, w_eco65821, w_eco65822, w_eco65823, w_eco65824, w_eco65825, w_eco65826, w_eco65827, w_eco65828, w_eco65829, w_eco65830, w_eco65831, w_eco65832, w_eco65833, w_eco65834, w_eco65835, w_eco65836, w_eco65837, w_eco65838, w_eco65839, w_eco65840, w_eco65841, w_eco65842, w_eco65843, w_eco65844, w_eco65845, w_eco65846, w_eco65847, w_eco65848, w_eco65849, w_eco65850, w_eco65851, w_eco65852, w_eco65853, w_eco65854, w_eco65855, w_eco65856, w_eco65857, w_eco65858, w_eco65859, w_eco65860, w_eco65861, w_eco65862, w_eco65863, w_eco65864, w_eco65865, w_eco65866, w_eco65867, w_eco65868, w_eco65869, w_eco65870, w_eco65871, w_eco65872, w_eco65873, w_eco65874, w_eco65875, w_eco65876, w_eco65877, w_eco65878, w_eco65879, w_eco65880, w_eco65881, w_eco65882, w_eco65883, w_eco65884, w_eco65885, w_eco65886, w_eco65887, w_eco65888, w_eco65889, w_eco65890, w_eco65891, w_eco65892, w_eco65893, w_eco65894, w_eco65895, w_eco65896, w_eco65897, w_eco65898, w_eco65899, w_eco65900, w_eco65901, w_eco65902, w_eco65903, w_eco65904, w_eco65905, w_eco65906, w_eco65907, w_eco65908, w_eco65909, w_eco65910, w_eco65911, w_eco65912, w_eco65913, w_eco65914, w_eco65915, w_eco65916, w_eco65917, w_eco65918, w_eco65919, w_eco65920, w_eco65921, w_eco65922, w_eco65923, w_eco65924, w_eco65925, w_eco65926, w_eco65927, w_eco65928, w_eco65929, w_eco65930, w_eco65931, w_eco65932, w_eco65933, w_eco65934, w_eco65935, w_eco65936, w_eco65937, w_eco65938, w_eco65939, w_eco65940, w_eco65941, w_eco65942, w_eco65943, w_eco65944, w_eco65945, w_eco65946, w_eco65947, w_eco65948, w_eco65949, w_eco65950, w_eco65951, w_eco65952, w_eco65953, w_eco65954, w_eco65955, w_eco65956, w_eco65957, w_eco65958, w_eco65959, w_eco65960, w_eco65961, w_eco65962, w_eco65963, w_eco65964, w_eco65965, w_eco65966, w_eco65967, w_eco65968, w_eco65969, w_eco65970, w_eco65971, w_eco65972, w_eco65973, w_eco65974, w_eco65975, w_eco65976, w_eco65977, w_eco65978, w_eco65979, w_eco65980, w_eco65981, w_eco65982, w_eco65983, w_eco65984, w_eco65985, w_eco65986, w_eco65987, w_eco65988, w_eco65989, w_eco65990, w_eco65991, w_eco65992, w_eco65993, w_eco65994, w_eco65995, w_eco65996, w_eco65997, w_eco65998, w_eco65999, w_eco66000, w_eco66001, w_eco66002, w_eco66003, w_eco66004, w_eco66005, w_eco66006, w_eco66007, w_eco66008, w_eco66009, w_eco66010, w_eco66011, w_eco66012, w_eco66013, w_eco66014, w_eco66015, w_eco66016, w_eco66017, w_eco66018, w_eco66019, w_eco66020, w_eco66021, w_eco66022, w_eco66023, w_eco66024, w_eco66025, w_eco66026, w_eco66027, w_eco66028, w_eco66029, w_eco66030, w_eco66031, w_eco66032, w_eco66033, w_eco66034, w_eco66035, w_eco66036, w_eco66037, w_eco66038, w_eco66039, w_eco66040, w_eco66041, w_eco66042, w_eco66043, w_eco66044, w_eco66045, w_eco66046, w_eco66047, w_eco66048, w_eco66049, w_eco66050, w_eco66051, w_eco66052, w_eco66053, w_eco66054, w_eco66055, w_eco66056, w_eco66057, w_eco66058, w_eco66059, w_eco66060, w_eco66061, w_eco66062, w_eco66063, w_eco66064, w_eco66065, w_eco66066, w_eco66067, w_eco66068, w_eco66069, w_eco66070, w_eco66071, w_eco66072, w_eco66073, w_eco66074, w_eco66075, w_eco66076, w_eco66077, w_eco66078, w_eco66079, w_eco66080, w_eco66081, w_eco66082, w_eco66083, w_eco66084, w_eco66085, w_eco66086, w_eco66087, w_eco66088, w_eco66089, w_eco66090, w_eco66091, w_eco66092, w_eco66093, w_eco66094, w_eco66095, w_eco66096, w_eco66097, w_eco66098, w_eco66099, w_eco66100, w_eco66101, w_eco66102, w_eco66103, w_eco66104, w_eco66105, w_eco66106, w_eco66107, w_eco66108, w_eco66109, w_eco66110, w_eco66111, w_eco66112, w_eco66113, w_eco66114, w_eco66115, w_eco66116, w_eco66117, w_eco66118, w_eco66119, w_eco66120, w_eco66121, w_eco66122, w_eco66123, w_eco66124, w_eco66125, w_eco66126, w_eco66127, w_eco66128, w_eco66129, w_eco66130, w_eco66131, w_eco66132, w_eco66133, w_eco66134, w_eco66135, w_eco66136, w_eco66137, w_eco66138, w_eco66139, w_eco66140, w_eco66141, w_eco66142, w_eco66143, w_eco66144, w_eco66145, w_eco66146, w_eco66147, w_eco66148, w_eco66149, w_eco66150, w_eco66151, w_eco66152, w_eco66153, w_eco66154, w_eco66155, w_eco66156, w_eco66157, w_eco66158, w_eco66159, w_eco66160, w_eco66161, w_eco66162, w_eco66163, w_eco66164, w_eco66165, w_eco66166, w_eco66167, w_eco66168, w_eco66169, w_eco66170, w_eco66171, w_eco66172, w_eco66173, w_eco66174, w_eco66175, w_eco66176, w_eco66177, w_eco66178, w_eco66179, w_eco66180, w_eco66181, w_eco66182, w_eco66183, w_eco66184, w_eco66185, w_eco66186, w_eco66187, w_eco66188, w_eco66189, w_eco66190, w_eco66191, w_eco66192, w_eco66193, w_eco66194, w_eco66195, w_eco66196, w_eco66197, w_eco66198, w_eco66199, w_eco66200, w_eco66201, w_eco66202, w_eco66203, w_eco66204, w_eco66205, w_eco66206, w_eco66207, w_eco66208, w_eco66209, w_eco66210, w_eco66211, w_eco66212, w_eco66213, w_eco66214, w_eco66215, w_eco66216, w_eco66217, w_eco66218, w_eco66219, w_eco66220, w_eco66221, w_eco66222, w_eco66223, w_eco66224, w_eco66225, w_eco66226, w_eco66227, w_eco66228, w_eco66229, w_eco66230, w_eco66231, w_eco66232, w_eco66233, w_eco66234, w_eco66235, w_eco66236, w_eco66237, w_eco66238, w_eco66239, w_eco66240, w_eco66241, w_eco66242, w_eco66243, w_eco66244, w_eco66245, w_eco66246, w_eco66247, w_eco66248, w_eco66249, w_eco66250, w_eco66251, w_eco66252, w_eco66253, w_eco66254, w_eco66255, w_eco66256, w_eco66257, w_eco66258, w_eco66259, w_eco66260, w_eco66261, w_eco66262, w_eco66263, w_eco66264, w_eco66265, w_eco66266, w_eco66267, w_eco66268, w_eco66269, w_eco66270, w_eco66271, w_eco66272, w_eco66273, w_eco66274, w_eco66275, w_eco66276, w_eco66277, w_eco66278, w_eco66279, w_eco66280, w_eco66281, w_eco66282, w_eco66283, w_eco66284, w_eco66285, w_eco66286, w_eco66287, w_eco66288, w_eco66289, w_eco66290, w_eco66291, w_eco66292, w_eco66293, w_eco66294, w_eco66295, w_eco66296, w_eco66297, w_eco66298, w_eco66299, w_eco66300, w_eco66301, w_eco66302, w_eco66303, w_eco66304, w_eco66305, w_eco66306, w_eco66307, w_eco66308, w_eco66309, w_eco66310, w_eco66311, w_eco66312, w_eco66313, w_eco66314, w_eco66315, w_eco66316, w_eco66317, w_eco66318, w_eco66319, w_eco66320, w_eco66321, w_eco66322, w_eco66323, w_eco66324, w_eco66325, w_eco66326, w_eco66327, w_eco66328, w_eco66329, w_eco66330, w_eco66331, w_eco66332, w_eco66333, w_eco66334, w_eco66335, w_eco66336, w_eco66337, w_eco66338, w_eco66339, w_eco66340, w_eco66341, w_eco66342, w_eco66343, w_eco66344, w_eco66345, w_eco66346, w_eco66347, w_eco66348, w_eco66349, w_eco66350, w_eco66351, w_eco66352, w_eco66353, w_eco66354, w_eco66355, w_eco66356, w_eco66357, w_eco66358, w_eco66359, w_eco66360, w_eco66361, w_eco66362, w_eco66363, w_eco66364, w_eco66365, w_eco66366, w_eco66367, w_eco66368, w_eco66369, w_eco66370, w_eco66371, w_eco66372, w_eco66373, w_eco66374, w_eco66375, w_eco66376, w_eco66377, w_eco66378, w_eco66379, w_eco66380, w_eco66381, w_eco66382, w_eco66383, w_eco66384, w_eco66385, w_eco66386, w_eco66387, w_eco66388, w_eco66389, w_eco66390, w_eco66391, w_eco66392, w_eco66393, w_eco66394, w_eco66395, w_eco66396, w_eco66397, w_eco66398, w_eco66399, w_eco66400, w_eco66401, w_eco66402, w_eco66403, w_eco66404, w_eco66405, w_eco66406, w_eco66407, w_eco66408, w_eco66409, w_eco66410, w_eco66411, w_eco66412, w_eco66413, w_eco66414, w_eco66415, w_eco66416, w_eco66417, w_eco66418, w_eco66419, w_eco66420, w_eco66421, w_eco66422, w_eco66423, w_eco66424, w_eco66425, w_eco66426, w_eco66427, w_eco66428, w_eco66429, w_eco66430, w_eco66431, w_eco66432, w_eco66433, w_eco66434, w_eco66435, w_eco66436, w_eco66437, w_eco66438, w_eco66439, w_eco66440, w_eco66441, w_eco66442, w_eco66443, w_eco66444, w_eco66445, w_eco66446, w_eco66447, w_eco66448, w_eco66449, w_eco66450, w_eco66451, w_eco66452, w_eco66453, w_eco66454, w_eco66455, w_eco66456, w_eco66457, w_eco66458, w_eco66459, w_eco66460, w_eco66461, w_eco66462, w_eco66463, w_eco66464, w_eco66465, w_eco66466, w_eco66467, w_eco66468, w_eco66469, w_eco66470, w_eco66471, w_eco66472, w_eco66473, w_eco66474, w_eco66475, w_eco66476, w_eco66477, w_eco66478, w_eco66479, w_eco66480, w_eco66481, w_eco66482, w_eco66483, w_eco66484, w_eco66485, w_eco66486, w_eco66487, w_eco66488, w_eco66489, w_eco66490, w_eco66491, w_eco66492, w_eco66493, w_eco66494, w_eco66495, w_eco66496, w_eco66497, w_eco66498, w_eco66499, w_eco66500, w_eco66501, w_eco66502, w_eco66503, w_eco66504, w_eco66505, w_eco66506, w_eco66507, w_eco66508, w_eco66509, w_eco66510, w_eco66511, w_eco66512, w_eco66513, w_eco66514, w_eco66515, w_eco66516, w_eco66517, w_eco66518, w_eco66519, w_eco66520, w_eco66521, w_eco66522, w_eco66523, w_eco66524, w_eco66525, w_eco66526, w_eco66527, w_eco66528, w_eco66529, w_eco66530, w_eco66531, w_eco66532, w_eco66533, w_eco66534, w_eco66535, w_eco66536, w_eco66537, w_eco66538, w_eco66539, w_eco66540, w_eco66541, w_eco66542, w_eco66543, w_eco66544, w_eco66545, w_eco66546, w_eco66547, w_eco66548, w_eco66549, w_eco66550, w_eco66551, w_eco66552, w_eco66553, w_eco66554, w_eco66555, w_eco66556, w_eco66557, w_eco66558, w_eco66559, w_eco66560, w_eco66561, w_eco66562, w_eco66563, w_eco66564, w_eco66565, w_eco66566, w_eco66567, w_eco66568, w_eco66569, w_eco66570, w_eco66571, w_eco66572, w_eco66573, w_eco66574, w_eco66575, w_eco66576, w_eco66577, w_eco66578, w_eco66579, w_eco66580, w_eco66581, w_eco66582, w_eco66583, w_eco66584, w_eco66585, w_eco66586, w_eco66587, w_eco66588, w_eco66589, w_eco66590, w_eco66591, w_eco66592, w_eco66593, w_eco66594, w_eco66595, w_eco66596, w_eco66597, w_eco66598, w_eco66599, w_eco66600, w_eco66601, w_eco66602, w_eco66603, w_eco66604, w_eco66605, w_eco66606, w_eco66607, w_eco66608, w_eco66609, w_eco66610, w_eco66611, w_eco66612, w_eco66613, w_eco66614, w_eco66615, w_eco66616, w_eco66617, w_eco66618, w_eco66619, w_eco66620, w_eco66621, w_eco66622, w_eco66623, w_eco66624, w_eco66625, w_eco66626, w_eco66627, w_eco66628, w_eco66629, w_eco66630, w_eco66631, w_eco66632, w_eco66633, w_eco66634, w_eco66635, w_eco66636, w_eco66637, w_eco66638, w_eco66639, w_eco66640, w_eco66641, w_eco66642, w_eco66643, w_eco66644, w_eco66645, w_eco66646, w_eco66647, w_eco66648, w_eco66649, w_eco66650, w_eco66651, w_eco66652, w_eco66653, w_eco66654, w_eco66655, w_eco66656, w_eco66657, w_eco66658, w_eco66659, w_eco66660, w_eco66661, w_eco66662, w_eco66663, w_eco66664, w_eco66665, w_eco66666, w_eco66667, w_eco66668, w_eco66669, w_eco66670, w_eco66671, w_eco66672, w_eco66673, w_eco66674, w_eco66675, w_eco66676, w_eco66677, w_eco66678, w_eco66679, w_eco66680, w_eco66681, w_eco66682, w_eco66683, w_eco66684, w_eco66685, w_eco66686, w_eco66687, w_eco66688, w_eco66689, w_eco66690, w_eco66691, w_eco66692, w_eco66693, w_eco66694, w_eco66695, w_eco66696, w_eco66697, w_eco66698, w_eco66699, w_eco66700, w_eco66701, w_eco66702, w_eco66703, w_eco66704, w_eco66705, w_eco66706, w_eco66707, w_eco66708, w_eco66709, w_eco66710, w_eco66711, w_eco66712, w_eco66713, w_eco66714, w_eco66715, w_eco66716, w_eco66717, w_eco66718, w_eco66719, w_eco66720, w_eco66721, w_eco66722, w_eco66723, w_eco66724, w_eco66725, w_eco66726, w_eco66727, w_eco66728, w_eco66729, w_eco66730, w_eco66731, w_eco66732, w_eco66733, w_eco66734, w_eco66735, w_eco66736, w_eco66737, w_eco66738, w_eco66739, w_eco66740, w_eco66741, w_eco66742, w_eco66743, w_eco66744, w_eco66745, w_eco66746, w_eco66747, w_eco66748, w_eco66749, w_eco66750, w_eco66751, w_eco66752, w_eco66753, w_eco66754, w_eco66755, w_eco66756, w_eco66757, w_eco66758, w_eco66759, w_eco66760, w_eco66761, w_eco66762, w_eco66763, w_eco66764, w_eco66765, w_eco66766, w_eco66767, w_eco66768, w_eco66769, w_eco66770, w_eco66771, w_eco66772, w_eco66773, w_eco66774, w_eco66775, w_eco66776, w_eco66777, w_eco66778, w_eco66779, w_eco66780, w_eco66781, w_eco66782, w_eco66783, w_eco66784, w_eco66785, w_eco66786, w_eco66787, w_eco66788, w_eco66789, w_eco66790, w_eco66791, w_eco66792, w_eco66793, w_eco66794, w_eco66795, w_eco66796, w_eco66797, w_eco66798, w_eco66799, w_eco66800, w_eco66801, w_eco66802, w_eco66803, w_eco66804, w_eco66805, w_eco66806, w_eco66807, w_eco66808, w_eco66809, w_eco66810, w_eco66811, w_eco66812, w_eco66813, w_eco66814, w_eco66815, w_eco66816, w_eco66817, w_eco66818, w_eco66819, w_eco66820, w_eco66821, w_eco66822, w_eco66823, w_eco66824, w_eco66825, w_eco66826, w_eco66827, w_eco66828, w_eco66829, w_eco66830, w_eco66831, w_eco66832, w_eco66833, w_eco66834, w_eco66835, w_eco66836, w_eco66837, w_eco66838, w_eco66839, w_eco66840, w_eco66841, w_eco66842, w_eco66843, w_eco66844, w_eco66845, w_eco66846, w_eco66847, w_eco66848, w_eco66849, w_eco66850, w_eco66851, w_eco66852, w_eco66853, w_eco66854, w_eco66855, w_eco66856, w_eco66857, w_eco66858, w_eco66859, w_eco66860, w_eco66861, w_eco66862, w_eco66863, w_eco66864, w_eco66865, w_eco66866, w_eco66867, w_eco66868, w_eco66869, w_eco66870, w_eco66871, w_eco66872, w_eco66873, w_eco66874, w_eco66875, w_eco66876, w_eco66877, w_eco66878, w_eco66879, w_eco66880, w_eco66881, w_eco66882, w_eco66883, w_eco66884, w_eco66885, w_eco66886, w_eco66887, w_eco66888, w_eco66889, w_eco66890, w_eco66891, w_eco66892, w_eco66893, w_eco66894, w_eco66895, w_eco66896, w_eco66897, w_eco66898, w_eco66899, w_eco66900, w_eco66901, w_eco66902, w_eco66903, w_eco66904, w_eco66905, w_eco66906, w_eco66907, w_eco66908, w_eco66909, w_eco66910, w_eco66911, w_eco66912, w_eco66913, w_eco66914, w_eco66915, w_eco66916, w_eco66917, w_eco66918, w_eco66919, w_eco66920, w_eco66921, w_eco66922, w_eco66923, w_eco66924, w_eco66925, w_eco66926, w_eco66927, w_eco66928, w_eco66929, w_eco66930, w_eco66931, w_eco66932, w_eco66933, w_eco66934, w_eco66935, w_eco66936, w_eco66937, w_eco66938, w_eco66939, w_eco66940, w_eco66941, w_eco66942, w_eco66943, w_eco66944, w_eco66945, w_eco66946, w_eco66947, w_eco66948, w_eco66949, w_eco66950, w_eco66951, w_eco66952, w_eco66953, w_eco66954, w_eco66955, w_eco66956, w_eco66957, w_eco66958, w_eco66959, w_eco66960, w_eco66961, w_eco66962, w_eco66963, w_eco66964, w_eco66965, w_eco66966, w_eco66967, w_eco66968, w_eco66969, w_eco66970, w_eco66971, w_eco66972, w_eco66973, w_eco66974, w_eco66975, w_eco66976, w_eco66977, w_eco66978, w_eco66979, w_eco66980, w_eco66981, w_eco66982, w_eco66983, w_eco66984, w_eco66985, w_eco66986, w_eco66987, w_eco66988, w_eco66989, w_eco66990, w_eco66991, w_eco66992, w_eco66993, w_eco66994, w_eco66995, w_eco66996, w_eco66997, w_eco66998, w_eco66999, w_eco67000, w_eco67001, w_eco67002, w_eco67003, w_eco67004, w_eco67005, w_eco67006, w_eco67007, w_eco67008, w_eco67009, w_eco67010, w_eco67011, w_eco67012, w_eco67013, w_eco67014, w_eco67015, w_eco67016, w_eco67017, w_eco67018, w_eco67019, w_eco67020, w_eco67021, w_eco67022, w_eco67023, w_eco67024, w_eco67025, w_eco67026, w_eco67027, w_eco67028, w_eco67029, w_eco67030, w_eco67031, w_eco67032, w_eco67033, w_eco67034, w_eco67035, w_eco67036, w_eco67037, w_eco67038, w_eco67039, w_eco67040, w_eco67041, w_eco67042, w_eco67043, w_eco67044, w_eco67045, w_eco67046, w_eco67047, w_eco67048, w_eco67049, w_eco67050, w_eco67051, w_eco67052, w_eco67053, w_eco67054, w_eco67055, w_eco67056, w_eco67057, w_eco67058, w_eco67059, w_eco67060, w_eco67061, w_eco67062, w_eco67063, w_eco67064, w_eco67065, w_eco67066, w_eco67067, w_eco67068, w_eco67069, w_eco67070, w_eco67071, w_eco67072, w_eco67073, w_eco67074, w_eco67075, w_eco67076, w_eco67077, w_eco67078, w_eco67079, w_eco67080, w_eco67081, w_eco67082, w_eco67083, w_eco67084, w_eco67085, w_eco67086, w_eco67087, w_eco67088, w_eco67089, w_eco67090, w_eco67091, w_eco67092, w_eco67093, w_eco67094, w_eco67095, w_eco67096, w_eco67097, w_eco67098, w_eco67099, w_eco67100, w_eco67101, w_eco67102, w_eco67103, w_eco67104, w_eco67105, w_eco67106, w_eco67107, w_eco67108, w_eco67109, w_eco67110, w_eco67111, w_eco67112, w_eco67113, w_eco67114, w_eco67115, w_eco67116, w_eco67117, w_eco67118, w_eco67119, w_eco67120, w_eco67121, w_eco67122, w_eco67123, w_eco67124, w_eco67125, w_eco67126, w_eco67127, w_eco67128, w_eco67129, w_eco67130, w_eco67131, w_eco67132, w_eco67133, w_eco67134, w_eco67135, w_eco67136, w_eco67137, w_eco67138, w_eco67139, w_eco67140, w_eco67141, w_eco67142, w_eco67143, w_eco67144, w_eco67145, w_eco67146, w_eco67147, w_eco67148, w_eco67149, w_eco67150, w_eco67151, w_eco67152, w_eco67153, w_eco67154, w_eco67155, w_eco67156, w_eco67157, w_eco67158, w_eco67159, w_eco67160, w_eco67161, w_eco67162, w_eco67163, w_eco67164, w_eco67165, w_eco67166, w_eco67167, w_eco67168, w_eco67169, w_eco67170, w_eco67171, w_eco67172, w_eco67173, w_eco67174, w_eco67175, w_eco67176, w_eco67177, w_eco67178, w_eco67179, w_eco67180, w_eco67181, w_eco67182, w_eco67183, w_eco67184, w_eco67185, w_eco67186, w_eco67187, w_eco67188, w_eco67189, w_eco67190, w_eco67191, w_eco67192, w_eco67193, w_eco67194, w_eco67195, w_eco67196, w_eco67197, w_eco67198, w_eco67199, w_eco67200, w_eco67201, w_eco67202, w_eco67203, w_eco67204, w_eco67205, w_eco67206, w_eco67207, w_eco67208, w_eco67209, w_eco67210, w_eco67211, w_eco67212, w_eco67213, w_eco67214, w_eco67215, w_eco67216, w_eco67217, w_eco67218, w_eco67219, w_eco67220, w_eco67221, w_eco67222, w_eco67223, w_eco67224, w_eco67225, w_eco67226, w_eco67227, w_eco67228, w_eco67229, w_eco67230, w_eco67231, w_eco67232, w_eco67233, w_eco67234, w_eco67235, w_eco67236, w_eco67237, w_eco67238, w_eco67239, w_eco67240, w_eco67241, w_eco67242, w_eco67243, w_eco67244, w_eco67245, w_eco67246, w_eco67247, w_eco67248, w_eco67249, w_eco67250, w_eco67251, w_eco67252, w_eco67253, w_eco67254, w_eco67255, w_eco67256, w_eco67257, w_eco67258, w_eco67259, w_eco67260, w_eco67261, w_eco67262, w_eco67263, w_eco67264, w_eco67265, w_eco67266, w_eco67267, w_eco67268, w_eco67269, w_eco67270, w_eco67271, w_eco67272, w_eco67273, w_eco67274, w_eco67275, w_eco67276, w_eco67277, w_eco67278, w_eco67279, w_eco67280, w_eco67281, w_eco67282, w_eco67283, w_eco67284, w_eco67285, w_eco67286, w_eco67287, w_eco67288, w_eco67289, w_eco67290, w_eco67291, w_eco67292, w_eco67293, w_eco67294, w_eco67295, w_eco67296, w_eco67297, w_eco67298, w_eco67299, w_eco67300, w_eco67301, w_eco67302, w_eco67303, w_eco67304, w_eco67305, w_eco67306, w_eco67307, w_eco67308, w_eco67309, w_eco67310, w_eco67311, w_eco67312, w_eco67313, w_eco67314, w_eco67315, w_eco67316, w_eco67317, w_eco67318, w_eco67319, w_eco67320, w_eco67321, w_eco67322, w_eco67323, w_eco67324, w_eco67325, w_eco67326, w_eco67327, w_eco67328, w_eco67329, w_eco67330, w_eco67331, w_eco67332, w_eco67333, w_eco67334, w_eco67335, w_eco67336, w_eco67337, w_eco67338, w_eco67339, w_eco67340, w_eco67341, w_eco67342, w_eco67343, w_eco67344, w_eco67345, w_eco67346, w_eco67347, w_eco67348, w_eco67349, w_eco67350, w_eco67351, w_eco67352, w_eco67353, w_eco67354, w_eco67355, w_eco67356, w_eco67357, w_eco67358, w_eco67359, w_eco67360, w_eco67361, w_eco67362, w_eco67363, w_eco67364, w_eco67365, w_eco67366, w_eco67367, w_eco67368, w_eco67369, w_eco67370, w_eco67371, w_eco67372, w_eco67373, w_eco67374, w_eco67375, w_eco67376, w_eco67377, w_eco67378, w_eco67379, w_eco67380, w_eco67381, w_eco67382, w_eco67383, w_eco67384, w_eco67385, w_eco67386, w_eco67387, w_eco67388, w_eco67389, w_eco67390, w_eco67391, w_eco67392, w_eco67393, w_eco67394, w_eco67395, w_eco67396, w_eco67397, w_eco67398, w_eco67399, w_eco67400, w_eco67401, w_eco67402, w_eco67403, w_eco67404, w_eco67405, w_eco67406, w_eco67407, w_eco67408, w_eco67409, w_eco67410, w_eco67411, w_eco67412, w_eco67413, w_eco67414, w_eco67415, w_eco67416, w_eco67417, w_eco67418, w_eco67419, w_eco67420, w_eco67421, w_eco67422, w_eco67423, w_eco67424, w_eco67425, w_eco67426, w_eco67427, w_eco67428, w_eco67429, w_eco67430, w_eco67431, w_eco67432, w_eco67433, w_eco67434, w_eco67435, w_eco67436, w_eco67437, w_eco67438, w_eco67439, w_eco67440, w_eco67441, w_eco67442, w_eco67443, w_eco67444, w_eco67445, w_eco67446, w_eco67447, w_eco67448, w_eco67449, w_eco67450, w_eco67451, w_eco67452, w_eco67453, w_eco67454, w_eco67455, w_eco67456, w_eco67457, w_eco67458, w_eco67459, w_eco67460, w_eco67461, w_eco67462, w_eco67463, w_eco67464, w_eco67465, w_eco67466, w_eco67467, w_eco67468, w_eco67469, w_eco67470, w_eco67471, w_eco67472, w_eco67473, w_eco67474, w_eco67475, w_eco67476, w_eco67477, w_eco67478, w_eco67479, w_eco67480, w_eco67481, w_eco67482, w_eco67483, w_eco67484, w_eco67485, w_eco67486, w_eco67487, w_eco67488, w_eco67489, w_eco67490, w_eco67491, w_eco67492, w_eco67493, w_eco67494, w_eco67495, w_eco67496, w_eco67497, w_eco67498, w_eco67499, w_eco67500, w_eco67501, w_eco67502, w_eco67503, w_eco67504, w_eco67505, w_eco67506, w_eco67507, w_eco67508, w_eco67509, w_eco67510, w_eco67511, w_eco67512, w_eco67513, w_eco67514, w_eco67515, w_eco67516, w_eco67517, w_eco67518, w_eco67519, w_eco67520, w_eco67521, w_eco67522, w_eco67523, w_eco67524, w_eco67525, w_eco67526, w_eco67527, w_eco67528, w_eco67529, w_eco67530, w_eco67531, w_eco67532, w_eco67533, w_eco67534, w_eco67535, w_eco67536, w_eco67537, w_eco67538, w_eco67539, w_eco67540, w_eco67541, w_eco67542, w_eco67543, w_eco67544, w_eco67545, w_eco67546, w_eco67547, w_eco67548, w_eco67549, w_eco67550, w_eco67551, w_eco67552, w_eco67553, w_eco67554, w_eco67555, w_eco67556, w_eco67557, w_eco67558, w_eco67559, w_eco67560, w_eco67561, w_eco67562, w_eco67563, w_eco67564, w_eco67565, w_eco67566, w_eco67567, w_eco67568, w_eco67569, w_eco67570, w_eco67571, w_eco67572, w_eco67573, w_eco67574, w_eco67575, w_eco67576, w_eco67577, w_eco67578, w_eco67579, w_eco67580, w_eco67581, w_eco67582, w_eco67583, w_eco67584, w_eco67585, w_eco67586, w_eco67587, w_eco67588, w_eco67589, w_eco67590, w_eco67591, w_eco67592, w_eco67593, w_eco67594, w_eco67595, w_eco67596, w_eco67597, w_eco67598, w_eco67599, w_eco67600, w_eco67601, w_eco67602, w_eco67603, w_eco67604, w_eco67605, w_eco67606, w_eco67607, w_eco67608, w_eco67609, w_eco67610, w_eco67611, w_eco67612, w_eco67613, w_eco67614, w_eco67615, w_eco67616, w_eco67617, w_eco67618, w_eco67619, w_eco67620, w_eco67621, w_eco67622, w_eco67623, w_eco67624, w_eco67625, w_eco67626, w_eco67627, w_eco67628, w_eco67629, w_eco67630, w_eco67631, w_eco67632, w_eco67633, w_eco67634, w_eco67635, w_eco67636, w_eco67637, w_eco67638, w_eco67639, w_eco67640, w_eco67641, w_eco67642, w_eco67643, w_eco67644, w_eco67645, w_eco67646, w_eco67647, w_eco67648, w_eco67649, w_eco67650, w_eco67651, w_eco67652, w_eco67653, w_eco67654, w_eco67655, w_eco67656, w_eco67657, w_eco67658, w_eco67659, w_eco67660, w_eco67661, w_eco67662, w_eco67663, w_eco67664, w_eco67665, w_eco67666, w_eco67667, w_eco67668, w_eco67669, w_eco67670, w_eco67671, w_eco67672, w_eco67673, w_eco67674, w_eco67675, w_eco67676, w_eco67677, w_eco67678, w_eco67679, w_eco67680, w_eco67681, w_eco67682, w_eco67683, w_eco67684, w_eco67685, w_eco67686, w_eco67687, w_eco67688, w_eco67689, w_eco67690, w_eco67691, w_eco67692, w_eco67693, w_eco67694, w_eco67695, w_eco67696, w_eco67697, w_eco67698, w_eco67699, w_eco67700, w_eco67701, w_eco67702, w_eco67703, w_eco67704, w_eco67705, w_eco67706, w_eco67707, w_eco67708, w_eco67709, w_eco67710, w_eco67711, w_eco67712, w_eco67713, w_eco67714, w_eco67715, w_eco67716, w_eco67717, w_eco67718, w_eco67719, w_eco67720, w_eco67721, w_eco67722, w_eco67723, w_eco67724, w_eco67725, w_eco67726, w_eco67727, w_eco67728, w_eco67729, w_eco67730, w_eco67731, w_eco67732, w_eco67733, w_eco67734, w_eco67735, w_eco67736, w_eco67737, w_eco67738, w_eco67739, w_eco67740, w_eco67741, w_eco67742, w_eco67743, w_eco67744, w_eco67745, w_eco67746, w_eco67747, w_eco67748, w_eco67749, w_eco67750, w_eco67751, w_eco67752, w_eco67753, w_eco67754, w_eco67755, w_eco67756, w_eco67757, w_eco67758, w_eco67759, w_eco67760, w_eco67761, w_eco67762, w_eco67763, w_eco67764, w_eco67765, w_eco67766, w_eco67767, w_eco67768, w_eco67769, w_eco67770, w_eco67771, w_eco67772, w_eco67773, w_eco67774, w_eco67775, w_eco67776, w_eco67777, w_eco67778, w_eco67779, w_eco67780, w_eco67781, w_eco67782, w_eco67783, w_eco67784, w_eco67785, w_eco67786, w_eco67787, w_eco67788, w_eco67789, w_eco67790, w_eco67791, w_eco67792, w_eco67793, w_eco67794, w_eco67795, w_eco67796, w_eco67797, w_eco67798, w_eco67799, w_eco67800, w_eco67801, w_eco67802, w_eco67803, w_eco67804, w_eco67805, w_eco67806, w_eco67807, w_eco67808, w_eco67809, w_eco67810, w_eco67811, w_eco67812, w_eco67813, w_eco67814, w_eco67815, w_eco67816, w_eco67817, w_eco67818, w_eco67819, w_eco67820, w_eco67821, w_eco67822, w_eco67823, w_eco67824, w_eco67825, w_eco67826, w_eco67827, w_eco67828, w_eco67829, w_eco67830, w_eco67831, w_eco67832, w_eco67833, w_eco67834, w_eco67835, w_eco67836, w_eco67837, w_eco67838, w_eco67839, w_eco67840, w_eco67841, w_eco67842, w_eco67843, w_eco67844, w_eco67845, w_eco67846, w_eco67847, w_eco67848, w_eco67849, w_eco67850, w_eco67851, w_eco67852, w_eco67853, w_eco67854, w_eco67855, w_eco67856, w_eco67857, w_eco67858, w_eco67859, w_eco67860, w_eco67861, w_eco67862, w_eco67863, w_eco67864, w_eco67865, w_eco67866, w_eco67867, w_eco67868, w_eco67869, w_eco67870, w_eco67871, w_eco67872, w_eco67873, w_eco67874, w_eco67875, w_eco67876, w_eco67877, w_eco67878, w_eco67879, w_eco67880, w_eco67881, w_eco67882, w_eco67883, w_eco67884, w_eco67885, w_eco67886, w_eco67887, w_eco67888, w_eco67889, w_eco67890, w_eco67891, w_eco67892, w_eco67893, w_eco67894, w_eco67895, w_eco67896, w_eco67897, w_eco67898, w_eco67899, w_eco67900, w_eco67901, w_eco67902, w_eco67903, w_eco67904, w_eco67905, w_eco67906, w_eco67907, w_eco67908, w_eco67909, w_eco67910, w_eco67911, w_eco67912, w_eco67913, w_eco67914, w_eco67915, w_eco67916, w_eco67917, w_eco67918, w_eco67919, w_eco67920, w_eco67921, w_eco67922, w_eco67923, w_eco67924, w_eco67925, w_eco67926, w_eco67927, w_eco67928, w_eco67929, w_eco67930, w_eco67931, w_eco67932, w_eco67933, w_eco67934, w_eco67935, w_eco67936, w_eco67937, w_eco67938, w_eco67939, w_eco67940, w_eco67941, w_eco67942, w_eco67943, w_eco67944, w_eco67945, w_eco67946, w_eco67947, w_eco67948, w_eco67949, w_eco67950, w_eco67951, w_eco67952, w_eco67953, w_eco67954, w_eco67955, w_eco67956, w_eco67957, w_eco67958, w_eco67959, w_eco67960, w_eco67961, w_eco67962, w_eco67963, w_eco67964, w_eco67965, w_eco67966, w_eco67967, w_eco67968, w_eco67969, w_eco67970, w_eco67971, w_eco67972, w_eco67973, w_eco67974, w_eco67975, w_eco67976, w_eco67977, w_eco67978, w_eco67979, w_eco67980, w_eco67981, w_eco67982, w_eco67983, w_eco67984, w_eco67985, w_eco67986, w_eco67987, w_eco67988, w_eco67989, w_eco67990, w_eco67991, w_eco67992, w_eco67993, w_eco67994, w_eco67995, w_eco67996, w_eco67997, w_eco67998, w_eco67999, w_eco68000, w_eco68001, w_eco68002, w_eco68003, w_eco68004, w_eco68005, w_eco68006, w_eco68007, w_eco68008, w_eco68009, w_eco68010, w_eco68011, w_eco68012, w_eco68013, w_eco68014, w_eco68015, w_eco68016, w_eco68017, w_eco68018, w_eco68019, w_eco68020, w_eco68021, w_eco68022, w_eco68023, w_eco68024, w_eco68025, w_eco68026, w_eco68027, w_eco68028, w_eco68029, w_eco68030, w_eco68031, w_eco68032, w_eco68033, w_eco68034, w_eco68035, w_eco68036, w_eco68037, w_eco68038, w_eco68039, w_eco68040, w_eco68041, w_eco68042, w_eco68043, w_eco68044, w_eco68045, w_eco68046, w_eco68047, w_eco68048, w_eco68049, w_eco68050, w_eco68051, w_eco68052, w_eco68053, w_eco68054, w_eco68055, w_eco68056, w_eco68057, w_eco68058, w_eco68059, w_eco68060, w_eco68061, w_eco68062, w_eco68063, w_eco68064, w_eco68065, w_eco68066, w_eco68067, w_eco68068, w_eco68069, w_eco68070, w_eco68071, w_eco68072, w_eco68073, w_eco68074, w_eco68075, w_eco68076, w_eco68077, w_eco68078, w_eco68079, w_eco68080, w_eco68081, w_eco68082, w_eco68083, w_eco68084, w_eco68085, w_eco68086, w_eco68087, w_eco68088, w_eco68089, w_eco68090, w_eco68091, w_eco68092, w_eco68093, w_eco68094, w_eco68095, w_eco68096, w_eco68097, w_eco68098, w_eco68099, w_eco68100, w_eco68101, w_eco68102, w_eco68103, w_eco68104, w_eco68105, w_eco68106, w_eco68107, w_eco68108, w_eco68109, w_eco68110, w_eco68111, w_eco68112, w_eco68113, w_eco68114, w_eco68115, w_eco68116, w_eco68117, w_eco68118, w_eco68119, w_eco68120, w_eco68121, w_eco68122, w_eco68123, w_eco68124, w_eco68125, w_eco68126, w_eco68127, w_eco68128, w_eco68129, w_eco68130, w_eco68131, w_eco68132, w_eco68133, w_eco68134, w_eco68135, w_eco68136, w_eco68137, w_eco68138, w_eco68139, w_eco68140, w_eco68141, w_eco68142, w_eco68143, w_eco68144, w_eco68145, w_eco68146, w_eco68147, w_eco68148, w_eco68149, w_eco68150, w_eco68151, w_eco68152, w_eco68153, w_eco68154, w_eco68155, w_eco68156, w_eco68157, w_eco68158, w_eco68159, w_eco68160, w_eco68161, w_eco68162, w_eco68163, w_eco68164, w_eco68165, w_eco68166, w_eco68167, w_eco68168, w_eco68169, w_eco68170, w_eco68171, w_eco68172, w_eco68173, w_eco68174, w_eco68175, w_eco68176, w_eco68177, w_eco68178, w_eco68179, w_eco68180, w_eco68181, w_eco68182, w_eco68183, w_eco68184, w_eco68185, w_eco68186, w_eco68187, w_eco68188, w_eco68189, w_eco68190, w_eco68191, w_eco68192, w_eco68193, w_eco68194, w_eco68195, w_eco68196, w_eco68197, w_eco68198, w_eco68199, w_eco68200, w_eco68201, w_eco68202, w_eco68203, w_eco68204, w_eco68205, w_eco68206, w_eco68207, w_eco68208, w_eco68209, w_eco68210, w_eco68211, w_eco68212, w_eco68213, w_eco68214, w_eco68215, w_eco68216, w_eco68217, w_eco68218, w_eco68219, w_eco68220, w_eco68221, w_eco68222, w_eco68223, w_eco68224, w_eco68225, w_eco68226, w_eco68227, w_eco68228, w_eco68229, w_eco68230, w_eco68231, w_eco68232, w_eco68233, w_eco68234, w_eco68235, w_eco68236, w_eco68237, w_eco68238, w_eco68239, w_eco68240, w_eco68241, w_eco68242, w_eco68243, w_eco68244, w_eco68245, w_eco68246, w_eco68247, w_eco68248, w_eco68249, w_eco68250, w_eco68251, w_eco68252, w_eco68253, w_eco68254, w_eco68255, w_eco68256, w_eco68257, w_eco68258, w_eco68259, w_eco68260, w_eco68261, w_eco68262, w_eco68263, w_eco68264, w_eco68265, w_eco68266, w_eco68267, w_eco68268, w_eco68269, w_eco68270, w_eco68271, w_eco68272, w_eco68273, w_eco68274, w_eco68275, w_eco68276, w_eco68277, w_eco68278, w_eco68279, w_eco68280, w_eco68281, w_eco68282, w_eco68283, w_eco68284, w_eco68285, w_eco68286, w_eco68287, w_eco68288, w_eco68289, w_eco68290, w_eco68291, w_eco68292, w_eco68293, w_eco68294, w_eco68295, w_eco68296, w_eco68297, w_eco68298, w_eco68299, w_eco68300, w_eco68301, w_eco68302, w_eco68303, w_eco68304, w_eco68305, w_eco68306, w_eco68307, w_eco68308, w_eco68309, w_eco68310, w_eco68311, w_eco68312, w_eco68313, w_eco68314, w_eco68315, w_eco68316, w_eco68317, w_eco68318, w_eco68319, w_eco68320, w_eco68321, w_eco68322, w_eco68323, w_eco68324, w_eco68325, w_eco68326, w_eco68327, w_eco68328, w_eco68329, w_eco68330, w_eco68331, w_eco68332, w_eco68333, w_eco68334, w_eco68335, w_eco68336, w_eco68337, w_eco68338, w_eco68339, w_eco68340, w_eco68341, w_eco68342, w_eco68343, w_eco68344, w_eco68345, w_eco68346, w_eco68347, w_eco68348, w_eco68349, w_eco68350, w_eco68351, w_eco68352, w_eco68353, w_eco68354, w_eco68355, w_eco68356, w_eco68357, w_eco68358, w_eco68359, w_eco68360, w_eco68361, w_eco68362, w_eco68363, w_eco68364, w_eco68365, w_eco68366, w_eco68367, w_eco68368, w_eco68369, w_eco68370, w_eco68371, w_eco68372, w_eco68373, w_eco68374, w_eco68375, w_eco68376, w_eco68377, w_eco68378, w_eco68379, w_eco68380, w_eco68381, w_eco68382, w_eco68383, w_eco68384, w_eco68385, w_eco68386, w_eco68387, w_eco68388, w_eco68389, w_eco68390, w_eco68391, w_eco68392, w_eco68393, w_eco68394, w_eco68395, w_eco68396, w_eco68397, w_eco68398, w_eco68399, w_eco68400, w_eco68401, w_eco68402, w_eco68403, w_eco68404, w_eco68405, w_eco68406, w_eco68407, w_eco68408, w_eco68409, w_eco68410, w_eco68411, w_eco68412, w_eco68413, w_eco68414, w_eco68415, w_eco68416, w_eco68417, w_eco68418, w_eco68419, w_eco68420, w_eco68421, w_eco68422, w_eco68423, w_eco68424, w_eco68425, w_eco68426, w_eco68427, w_eco68428, w_eco68429, w_eco68430, w_eco68431, w_eco68432, w_eco68433, w_eco68434, w_eco68435, w_eco68436, w_eco68437, w_eco68438, w_eco68439, w_eco68440, w_eco68441, w_eco68442, w_eco68443, w_eco68444, w_eco68445, w_eco68446, w_eco68447, w_eco68448, w_eco68449, w_eco68450, w_eco68451, w_eco68452, w_eco68453, w_eco68454, w_eco68455, w_eco68456, w_eco68457, w_eco68458, w_eco68459, w_eco68460, w_eco68461, w_eco68462, w_eco68463, w_eco68464, w_eco68465, w_eco68466, w_eco68467, w_eco68468, w_eco68469, w_eco68470, w_eco68471, w_eco68472, w_eco68473, w_eco68474, w_eco68475, w_eco68476, w_eco68477, w_eco68478, w_eco68479, w_eco68480, w_eco68481, w_eco68482, w_eco68483, w_eco68484, w_eco68485, w_eco68486, w_eco68487, w_eco68488, w_eco68489, w_eco68490, w_eco68491, w_eco68492, w_eco68493, w_eco68494, w_eco68495, w_eco68496, w_eco68497, w_eco68498, w_eco68499, w_eco68500, w_eco68501, w_eco68502, w_eco68503, w_eco68504, w_eco68505, w_eco68506, w_eco68507, w_eco68508, w_eco68509, w_eco68510, w_eco68511, w_eco68512, w_eco68513, w_eco68514, w_eco68515, w_eco68516, w_eco68517, w_eco68518, w_eco68519, w_eco68520, w_eco68521, w_eco68522, w_eco68523, w_eco68524, w_eco68525, w_eco68526, w_eco68527, w_eco68528, w_eco68529, w_eco68530, w_eco68531, w_eco68532, w_eco68533, w_eco68534, w_eco68535, w_eco68536, w_eco68537, w_eco68538, w_eco68539, w_eco68540, w_eco68541, w_eco68542, w_eco68543, w_eco68544, w_eco68545, w_eco68546, w_eco68547, w_eco68548, w_eco68549, w_eco68550, w_eco68551, w_eco68552, w_eco68553, w_eco68554, w_eco68555, w_eco68556, w_eco68557, w_eco68558, w_eco68559, w_eco68560, w_eco68561, w_eco68562, w_eco68563, w_eco68564, w_eco68565, w_eco68566, w_eco68567, w_eco68568, w_eco68569, w_eco68570, w_eco68571, w_eco68572, w_eco68573, w_eco68574, w_eco68575, w_eco68576, w_eco68577, w_eco68578, w_eco68579, w_eco68580, w_eco68581, w_eco68582, w_eco68583, w_eco68584, w_eco68585, w_eco68586, w_eco68587, w_eco68588, w_eco68589, w_eco68590, w_eco68591, w_eco68592, w_eco68593, w_eco68594, w_eco68595, w_eco68596, w_eco68597, w_eco68598, w_eco68599, w_eco68600, w_eco68601, w_eco68602, w_eco68603, w_eco68604, w_eco68605, w_eco68606, w_eco68607, w_eco68608, w_eco68609, w_eco68610, w_eco68611, w_eco68612, w_eco68613, w_eco68614, w_eco68615, w_eco68616, w_eco68617, w_eco68618, w_eco68619, w_eco68620, w_eco68621, w_eco68622, w_eco68623, w_eco68624, w_eco68625, w_eco68626, w_eco68627, w_eco68628, w_eco68629, w_eco68630, w_eco68631, w_eco68632, w_eco68633, w_eco68634, w_eco68635, w_eco68636, w_eco68637, w_eco68638, w_eco68639, w_eco68640, w_eco68641, w_eco68642, w_eco68643, w_eco68644, w_eco68645, w_eco68646, w_eco68647, w_eco68648, w_eco68649, w_eco68650, w_eco68651, w_eco68652, w_eco68653, w_eco68654, w_eco68655, w_eco68656, w_eco68657, w_eco68658, w_eco68659, w_eco68660, w_eco68661, w_eco68662, w_eco68663, w_eco68664, w_eco68665, w_eco68666, w_eco68667, w_eco68668, w_eco68669, w_eco68670, w_eco68671, w_eco68672, w_eco68673, w_eco68674, w_eco68675, w_eco68676, w_eco68677, w_eco68678, w_eco68679, w_eco68680, w_eco68681, w_eco68682, w_eco68683, w_eco68684, w_eco68685, w_eco68686, w_eco68687, w_eco68688, w_eco68689, w_eco68690, w_eco68691, w_eco68692, w_eco68693, w_eco68694, w_eco68695, w_eco68696, w_eco68697, w_eco68698, w_eco68699, w_eco68700, w_eco68701, w_eco68702, w_eco68703, w_eco68704, w_eco68705, w_eco68706, w_eco68707, w_eco68708, w_eco68709, w_eco68710, w_eco68711, w_eco68712, w_eco68713, w_eco68714, w_eco68715, w_eco68716, w_eco68717, w_eco68718, w_eco68719, w_eco68720, w_eco68721, w_eco68722, w_eco68723, w_eco68724, w_eco68725, w_eco68726, w_eco68727, w_eco68728, w_eco68729, w_eco68730, w_eco68731, w_eco68732, w_eco68733, w_eco68734, w_eco68735, w_eco68736, w_eco68737, w_eco68738, w_eco68739, w_eco68740, w_eco68741, w_eco68742, w_eco68743, w_eco68744, w_eco68745, w_eco68746, w_eco68747, w_eco68748, w_eco68749, w_eco68750, w_eco68751, w_eco68752, w_eco68753, w_eco68754, w_eco68755, w_eco68756, w_eco68757, w_eco68758, w_eco68759, w_eco68760, w_eco68761, w_eco68762, w_eco68763, w_eco68764, w_eco68765, w_eco68766, w_eco68767, w_eco68768, w_eco68769, w_eco68770, w_eco68771, w_eco68772, w_eco68773, w_eco68774, w_eco68775, w_eco68776, w_eco68777, w_eco68778, w_eco68779, w_eco68780, w_eco68781, w_eco68782, w_eco68783, w_eco68784, w_eco68785, w_eco68786, w_eco68787, w_eco68788, w_eco68789, w_eco68790, w_eco68791, w_eco68792, w_eco68793, w_eco68794, w_eco68795, w_eco68796, w_eco68797, w_eco68798, w_eco68799, w_eco68800, w_eco68801, w_eco68802, w_eco68803, w_eco68804, w_eco68805, w_eco68806, w_eco68807, w_eco68808, w_eco68809, w_eco68810, w_eco68811, w_eco68812, w_eco68813, w_eco68814, w_eco68815, w_eco68816, w_eco68817, w_eco68818, w_eco68819, w_eco68820, w_eco68821, w_eco68822, w_eco68823, w_eco68824, w_eco68825, w_eco68826, w_eco68827, w_eco68828, w_eco68829, w_eco68830, w_eco68831, w_eco68832, w_eco68833, w_eco68834, w_eco68835, w_eco68836, w_eco68837, w_eco68838, w_eco68839, w_eco68840, w_eco68841, w_eco68842, w_eco68843, w_eco68844, w_eco68845, w_eco68846, w_eco68847, w_eco68848, w_eco68849, w_eco68850, w_eco68851, w_eco68852, w_eco68853, w_eco68854, w_eco68855, w_eco68856, w_eco68857, w_eco68858, w_eco68859, w_eco68860, w_eco68861, w_eco68862, w_eco68863, w_eco68864, w_eco68865, w_eco68866, w_eco68867, w_eco68868, w_eco68869, w_eco68870, w_eco68871, w_eco68872, w_eco68873, w_eco68874, w_eco68875, w_eco68876, w_eco68877, w_eco68878, w_eco68879, w_eco68880, w_eco68881, w_eco68882, w_eco68883, w_eco68884, w_eco68885, w_eco68886, w_eco68887, w_eco68888, w_eco68889, w_eco68890, w_eco68891, w_eco68892, w_eco68893, w_eco68894, w_eco68895, w_eco68896, w_eco68897, w_eco68898, w_eco68899, w_eco68900, w_eco68901, w_eco68902, w_eco68903, w_eco68904, w_eco68905, w_eco68906, w_eco68907, w_eco68908, w_eco68909, w_eco68910, w_eco68911, w_eco68912, w_eco68913, w_eco68914, w_eco68915, w_eco68916, w_eco68917, w_eco68918, w_eco68919, w_eco68920, w_eco68921, w_eco68922, w_eco68923, w_eco68924, w_eco68925, w_eco68926, w_eco68927, w_eco68928, w_eco68929, w_eco68930, w_eco68931, w_eco68932, w_eco68933, w_eco68934, w_eco68935, w_eco68936, w_eco68937, w_eco68938, w_eco68939, w_eco68940, w_eco68941, w_eco68942, w_eco68943, w_eco68944, w_eco68945, w_eco68946, w_eco68947, w_eco68948, w_eco68949, w_eco68950, w_eco68951, w_eco68952, w_eco68953, w_eco68954, w_eco68955, w_eco68956, w_eco68957, w_eco68958, w_eco68959, w_eco68960, w_eco68961, w_eco68962, w_eco68963, w_eco68964, w_eco68965, w_eco68966, w_eco68967, w_eco68968, w_eco68969, w_eco68970, w_eco68971, w_eco68972, w_eco68973, w_eco68974, w_eco68975, w_eco68976, w_eco68977, w_eco68978, w_eco68979, w_eco68980, w_eco68981, w_eco68982, w_eco68983, w_eco68984, w_eco68985, w_eco68986, w_eco68987, w_eco68988, w_eco68989, w_eco68990, w_eco68991, w_eco68992, w_eco68993, w_eco68994, w_eco68995, w_eco68996, w_eco68997, w_eco68998, w_eco68999, w_eco69000, w_eco69001, w_eco69002, w_eco69003, w_eco69004, w_eco69005, w_eco69006, w_eco69007, w_eco69008, w_eco69009, w_eco69010, w_eco69011, w_eco69012, w_eco69013, w_eco69014, w_eco69015, w_eco69016, w_eco69017, w_eco69018, w_eco69019, w_eco69020, w_eco69021, w_eco69022, w_eco69023, w_eco69024, w_eco69025, w_eco69026, w_eco69027, w_eco69028, w_eco69029, w_eco69030, w_eco69031, w_eco69032, w_eco69033, w_eco69034, w_eco69035, w_eco69036, w_eco69037, w_eco69038, w_eco69039, w_eco69040, w_eco69041, w_eco69042, w_eco69043, w_eco69044, w_eco69045, w_eco69046, w_eco69047, w_eco69048, w_eco69049, w_eco69050, w_eco69051, w_eco69052, w_eco69053, w_eco69054, w_eco69055, w_eco69056, w_eco69057, w_eco69058, w_eco69059, w_eco69060, w_eco69061, w_eco69062, w_eco69063, w_eco69064, w_eco69065, w_eco69066, w_eco69067, w_eco69068, w_eco69069, w_eco69070, w_eco69071, w_eco69072, w_eco69073, w_eco69074, w_eco69075, w_eco69076, w_eco69077, w_eco69078, w_eco69079, w_eco69080, w_eco69081, w_eco69082, w_eco69083, w_eco69084, w_eco69085, w_eco69086, w_eco69087, w_eco69088, w_eco69089, w_eco69090, w_eco69091, w_eco69092, w_eco69093, w_eco69094, w_eco69095, w_eco69096, w_eco69097, w_eco69098, w_eco69099, w_eco69100, w_eco69101, w_eco69102, w_eco69103, w_eco69104, w_eco69105, w_eco69106, w_eco69107, w_eco69108, w_eco69109, w_eco69110, w_eco69111, w_eco69112, w_eco69113, w_eco69114, w_eco69115, w_eco69116, w_eco69117, w_eco69118, w_eco69119, w_eco69120, w_eco69121, w_eco69122, w_eco69123, w_eco69124, w_eco69125, w_eco69126, w_eco69127, w_eco69128, w_eco69129, w_eco69130, w_eco69131, w_eco69132, w_eco69133, w_eco69134, w_eco69135, w_eco69136, w_eco69137, w_eco69138, w_eco69139, w_eco69140, w_eco69141, w_eco69142, w_eco69143, w_eco69144, w_eco69145, w_eco69146, w_eco69147, w_eco69148, w_eco69149, w_eco69150, w_eco69151, w_eco69152, w_eco69153, w_eco69154, w_eco69155, w_eco69156, w_eco69157, w_eco69158, w_eco69159, w_eco69160, w_eco69161, w_eco69162, w_eco69163, w_eco69164, w_eco69165, w_eco69166, w_eco69167, w_eco69168, w_eco69169, w_eco69170, w_eco69171, w_eco69172, w_eco69173, w_eco69174, w_eco69175, w_eco69176, w_eco69177, w_eco69178, w_eco69179, w_eco69180, w_eco69181, w_eco69182, w_eco69183, w_eco69184, w_eco69185, w_eco69186, w_eco69187, w_eco69188, w_eco69189, w_eco69190, w_eco69191, w_eco69192, w_eco69193, w_eco69194, w_eco69195, w_eco69196, w_eco69197, w_eco69198, w_eco69199, w_eco69200, w_eco69201, w_eco69202, w_eco69203, w_eco69204, w_eco69205, w_eco69206, w_eco69207, w_eco69208, w_eco69209, w_eco69210, w_eco69211, w_eco69212, w_eco69213, w_eco69214, w_eco69215, w_eco69216, w_eco69217, w_eco69218, w_eco69219, w_eco69220, w_eco69221, w_eco69222, w_eco69223, w_eco69224, w_eco69225, w_eco69226, w_eco69227, w_eco69228, w_eco69229, w_eco69230, w_eco69231, w_eco69232, w_eco69233, w_eco69234, w_eco69235, w_eco69236, w_eco69237, w_eco69238, w_eco69239, w_eco69240, w_eco69241, w_eco69242, w_eco69243, w_eco69244, w_eco69245, w_eco69246, w_eco69247, w_eco69248, w_eco69249, w_eco69250, w_eco69251, w_eco69252, w_eco69253, w_eco69254, w_eco69255, w_eco69256, w_eco69257, w_eco69258, w_eco69259, w_eco69260, w_eco69261, w_eco69262, w_eco69263, w_eco69264, w_eco69265, w_eco69266, w_eco69267, w_eco69268, w_eco69269, w_eco69270, w_eco69271, w_eco69272, w_eco69273, w_eco69274, w_eco69275, w_eco69276, w_eco69277, w_eco69278, w_eco69279, w_eco69280, w_eco69281, w_eco69282, w_eco69283, w_eco69284, w_eco69285, w_eco69286, w_eco69287, w_eco69288, w_eco69289, w_eco69290, w_eco69291, w_eco69292, w_eco69293, w_eco69294, w_eco69295, w_eco69296, w_eco69297, w_eco69298, w_eco69299, w_eco69300, w_eco69301, w_eco69302, w_eco69303, w_eco69304, w_eco69305, w_eco69306, w_eco69307, w_eco69308, w_eco69309, w_eco69310, w_eco69311, w_eco69312, w_eco69313, w_eco69314, w_eco69315, w_eco69316, w_eco69317, w_eco69318, w_eco69319, w_eco69320, w_eco69321, w_eco69322, w_eco69323, w_eco69324, w_eco69325, w_eco69326, w_eco69327, w_eco69328, w_eco69329, w_eco69330, w_eco69331, w_eco69332, w_eco69333, w_eco69334, w_eco69335, w_eco69336, w_eco69337, w_eco69338, w_eco69339, w_eco69340, w_eco69341, w_eco69342, w_eco69343, w_eco69344, w_eco69345, w_eco69346, w_eco69347, w_eco69348, w_eco69349, w_eco69350, w_eco69351, w_eco69352, w_eco69353, w_eco69354, w_eco69355, w_eco69356, w_eco69357, w_eco69358, w_eco69359, w_eco69360, w_eco69361, w_eco69362, w_eco69363, w_eco69364, w_eco69365, w_eco69366, w_eco69367, w_eco69368, w_eco69369, w_eco69370, w_eco69371, w_eco69372, w_eco69373, w_eco69374, w_eco69375, w_eco69376, w_eco69377, w_eco69378, w_eco69379, w_eco69380, w_eco69381, w_eco69382, w_eco69383, w_eco69384, w_eco69385, w_eco69386, w_eco69387, w_eco69388, w_eco69389, w_eco69390, w_eco69391, w_eco69392, w_eco69393, w_eco69394, w_eco69395, w_eco69396, w_eco69397, w_eco69398, w_eco69399, w_eco69400, w_eco69401, w_eco69402, w_eco69403, w_eco69404, w_eco69405, w_eco69406, w_eco69407, w_eco69408, w_eco69409, w_eco69410, w_eco69411, w_eco69412, w_eco69413, w_eco69414, w_eco69415, w_eco69416, w_eco69417, w_eco69418, w_eco69419, w_eco69420, w_eco69421, w_eco69422, w_eco69423, w_eco69424, w_eco69425, w_eco69426, w_eco69427, w_eco69428, w_eco69429, w_eco69430, w_eco69431, w_eco69432, w_eco69433, w_eco69434, w_eco69435, w_eco69436, w_eco69437, w_eco69438, w_eco69439, w_eco69440, w_eco69441, w_eco69442, w_eco69443, w_eco69444, w_eco69445, w_eco69446, w_eco69447, w_eco69448, w_eco69449, w_eco69450, w_eco69451, w_eco69452, w_eco69453, w_eco69454, w_eco69455, w_eco69456, w_eco69457, w_eco69458, w_eco69459, w_eco69460, w_eco69461, w_eco69462, w_eco69463, w_eco69464, w_eco69465, w_eco69466, w_eco69467, w_eco69468, w_eco69469, w_eco69470, w_eco69471, w_eco69472, w_eco69473, w_eco69474, w_eco69475, w_eco69476, w_eco69477, w_eco69478, w_eco69479, w_eco69480, w_eco69481, w_eco69482, w_eco69483, w_eco69484, w_eco69485, w_eco69486, w_eco69487, w_eco69488, w_eco69489, w_eco69490, w_eco69491, w_eco69492, w_eco69493, w_eco69494, w_eco69495, w_eco69496, w_eco69497, w_eco69498, w_eco69499, w_eco69500, w_eco69501, w_eco69502, w_eco69503, w_eco69504, w_eco69505, w_eco69506, w_eco69507, w_eco69508, w_eco69509, w_eco69510, w_eco69511, w_eco69512, w_eco69513, w_eco69514, w_eco69515, w_eco69516, w_eco69517, w_eco69518, w_eco69519, w_eco69520, w_eco69521, w_eco69522, w_eco69523, w_eco69524, w_eco69525, w_eco69526, w_eco69527, w_eco69528, w_eco69529, w_eco69530, w_eco69531, w_eco69532, w_eco69533, w_eco69534, w_eco69535, w_eco69536, w_eco69537, w_eco69538, w_eco69539, w_eco69540, w_eco69541, w_eco69542, w_eco69543, w_eco69544, w_eco69545, w_eco69546, w_eco69547, w_eco69548, w_eco69549, w_eco69550, w_eco69551, w_eco69552, w_eco69553, w_eco69554, w_eco69555, w_eco69556, w_eco69557, w_eco69558, w_eco69559, w_eco69560, w_eco69561, w_eco69562, w_eco69563, w_eco69564, w_eco69565, w_eco69566, w_eco69567, w_eco69568, w_eco69569, w_eco69570, w_eco69571, w_eco69572, w_eco69573, w_eco69574, w_eco69575, w_eco69576, w_eco69577, w_eco69578, w_eco69579, w_eco69580, w_eco69581, w_eco69582, w_eco69583, w_eco69584, w_eco69585, w_eco69586, w_eco69587, w_eco69588, w_eco69589, w_eco69590, w_eco69591, w_eco69592, w_eco69593, w_eco69594, w_eco69595, w_eco69596, w_eco69597, w_eco69598, w_eco69599, w_eco69600, w_eco69601, w_eco69602, w_eco69603, w_eco69604, w_eco69605, w_eco69606, w_eco69607, w_eco69608, w_eco69609, w_eco69610, w_eco69611, w_eco69612, w_eco69613, w_eco69614, w_eco69615, w_eco69616, w_eco69617, w_eco69618, w_eco69619, w_eco69620, w_eco69621, w_eco69622, w_eco69623, w_eco69624, w_eco69625, w_eco69626, w_eco69627, w_eco69628, w_eco69629, w_eco69630, w_eco69631, w_eco69632, w_eco69633, w_eco69634, w_eco69635, w_eco69636, w_eco69637, w_eco69638, w_eco69639, w_eco69640, w_eco69641, w_eco69642, w_eco69643, w_eco69644, w_eco69645, w_eco69646, w_eco69647, w_eco69648, w_eco69649, w_eco69650, w_eco69651, w_eco69652, w_eco69653, w_eco69654, w_eco69655, w_eco69656, w_eco69657, w_eco69658, w_eco69659, w_eco69660, w_eco69661, w_eco69662, w_eco69663, w_eco69664, w_eco69665, w_eco69666, w_eco69667, w_eco69668, w_eco69669, w_eco69670, w_eco69671, w_eco69672, w_eco69673, w_eco69674, w_eco69675, w_eco69676, w_eco69677, w_eco69678, w_eco69679, w_eco69680, w_eco69681, w_eco69682, w_eco69683, w_eco69684, w_eco69685, w_eco69686, w_eco69687, w_eco69688, w_eco69689, w_eco69690, w_eco69691, w_eco69692, w_eco69693, w_eco69694, w_eco69695, w_eco69696, w_eco69697, w_eco69698, w_eco69699, w_eco69700, w_eco69701, w_eco69702, w_eco69703, w_eco69704, w_eco69705, w_eco69706, w_eco69707, w_eco69708, w_eco69709, w_eco69710, w_eco69711, w_eco69712, w_eco69713, w_eco69714, w_eco69715, w_eco69716, w_eco69717, w_eco69718, w_eco69719, w_eco69720, w_eco69721, w_eco69722, w_eco69723, w_eco69724, w_eco69725, w_eco69726, w_eco69727, w_eco69728, w_eco69729, w_eco69730, w_eco69731, w_eco69732, w_eco69733, w_eco69734, w_eco69735, w_eco69736, w_eco69737, w_eco69738, w_eco69739, w_eco69740, w_eco69741, w_eco69742, w_eco69743, w_eco69744, w_eco69745, w_eco69746, w_eco69747, w_eco69748, w_eco69749, w_eco69750, w_eco69751, w_eco69752, w_eco69753, w_eco69754, w_eco69755, w_eco69756, w_eco69757, w_eco69758, w_eco69759, w_eco69760, w_eco69761, w_eco69762, w_eco69763, w_eco69764, w_eco69765, w_eco69766, w_eco69767, w_eco69768, w_eco69769, w_eco69770, w_eco69771, w_eco69772, w_eco69773, w_eco69774, w_eco69775, w_eco69776, w_eco69777, w_eco69778, w_eco69779, w_eco69780, w_eco69781, w_eco69782, w_eco69783, w_eco69784, w_eco69785, w_eco69786, w_eco69787, w_eco69788, w_eco69789, w_eco69790, w_eco69791, w_eco69792, w_eco69793, w_eco69794, w_eco69795, w_eco69796, w_eco69797, w_eco69798, w_eco69799, w_eco69800, w_eco69801, w_eco69802, w_eco69803, w_eco69804, w_eco69805, w_eco69806, w_eco69807, w_eco69808, w_eco69809, w_eco69810, w_eco69811, w_eco69812, w_eco69813, w_eco69814, w_eco69815, w_eco69816, w_eco69817, w_eco69818, w_eco69819, w_eco69820, w_eco69821, w_eco69822, w_eco69823, w_eco69824, w_eco69825, w_eco69826, w_eco69827, w_eco69828, w_eco69829, w_eco69830, w_eco69831, w_eco69832, w_eco69833, w_eco69834, w_eco69835, w_eco69836, w_eco69837, w_eco69838, w_eco69839, w_eco69840, w_eco69841, w_eco69842, w_eco69843, w_eco69844, w_eco69845, w_eco69846, w_eco69847, w_eco69848, w_eco69849, w_eco69850, w_eco69851, w_eco69852, w_eco69853, w_eco69854, w_eco69855, w_eco69856, w_eco69857, w_eco69858, w_eco69859, w_eco69860, w_eco69861, w_eco69862, w_eco69863, w_eco69864, w_eco69865, w_eco69866, w_eco69867, w_eco69868, w_eco69869, w_eco69870, w_eco69871, w_eco69872, w_eco69873, w_eco69874, w_eco69875, w_eco69876, w_eco69877, w_eco69878, w_eco69879, w_eco69880, w_eco69881, w_eco69882, w_eco69883, w_eco69884, w_eco69885, w_eco69886, w_eco69887, w_eco69888, w_eco69889, w_eco69890, w_eco69891, w_eco69892, w_eco69893, w_eco69894, w_eco69895, w_eco69896, w_eco69897, w_eco69898, w_eco69899, w_eco69900, w_eco69901, w_eco69902, w_eco69903, w_eco69904, w_eco69905, w_eco69906, w_eco69907, w_eco69908, w_eco69909, w_eco69910, w_eco69911, w_eco69912, w_eco69913, w_eco69914, w_eco69915, w_eco69916, w_eco69917, w_eco69918, w_eco69919, w_eco69920, w_eco69921, w_eco69922, w_eco69923, w_eco69924, w_eco69925, w_eco69926, w_eco69927, w_eco69928, w_eco69929, w_eco69930, w_eco69931, w_eco69932, w_eco69933, w_eco69934, w_eco69935, w_eco69936, w_eco69937, w_eco69938, w_eco69939, w_eco69940, w_eco69941, w_eco69942, w_eco69943, w_eco69944, w_eco69945, w_eco69946, w_eco69947, w_eco69948, w_eco69949, w_eco69950, w_eco69951, w_eco69952, w_eco69953, w_eco69954, w_eco69955, w_eco69956, w_eco69957, w_eco69958, w_eco69959, w_eco69960, w_eco69961, w_eco69962, w_eco69963, w_eco69964, w_eco69965, w_eco69966, w_eco69967, w_eco69968, w_eco69969, w_eco69970, w_eco69971, w_eco69972, w_eco69973, w_eco69974, w_eco69975, w_eco69976, w_eco69977, w_eco69978, w_eco69979, w_eco69980, w_eco69981, w_eco69982, w_eco69983, w_eco69984, w_eco69985, w_eco69986, w_eco69987, w_eco69988, w_eco69989, w_eco69990, w_eco69991, w_eco69992, w_eco69993, w_eco69994, w_eco69995, w_eco69996, w_eco69997, w_eco69998, w_eco69999, w_eco70000, w_eco70001, w_eco70002, w_eco70003, w_eco70004, w_eco70005, w_eco70006, w_eco70007, w_eco70008, w_eco70009, w_eco70010, w_eco70011, w_eco70012, w_eco70013, w_eco70014, w_eco70015, w_eco70016, w_eco70017, w_eco70018, w_eco70019, w_eco70020, w_eco70021, w_eco70022, w_eco70023, w_eco70024, w_eco70025, w_eco70026, w_eco70027, w_eco70028, w_eco70029, w_eco70030, w_eco70031, w_eco70032, w_eco70033, w_eco70034, w_eco70035, w_eco70036, w_eco70037, w_eco70038, w_eco70039, w_eco70040, w_eco70041, w_eco70042, w_eco70043, w_eco70044, w_eco70045, w_eco70046, w_eco70047, w_eco70048, w_eco70049, w_eco70050, w_eco70051, w_eco70052, w_eco70053, w_eco70054, w_eco70055, w_eco70056, w_eco70057, w_eco70058, w_eco70059, w_eco70060, w_eco70061, w_eco70062, w_eco70063, w_eco70064, w_eco70065, w_eco70066, w_eco70067, w_eco70068, w_eco70069, w_eco70070, w_eco70071, w_eco70072, w_eco70073, w_eco70074, w_eco70075, w_eco70076, w_eco70077, w_eco70078, w_eco70079, w_eco70080, w_eco70081, w_eco70082, w_eco70083, w_eco70084, w_eco70085, w_eco70086, w_eco70087, w_eco70088, w_eco70089, w_eco70090, w_eco70091, w_eco70092, w_eco70093, w_eco70094, w_eco70095, w_eco70096, w_eco70097, w_eco70098, w_eco70099, w_eco70100, w_eco70101, w_eco70102, w_eco70103, w_eco70104, w_eco70105, w_eco70106, w_eco70107, w_eco70108, w_eco70109, w_eco70110, w_eco70111, w_eco70112, w_eco70113, w_eco70114, w_eco70115, w_eco70116, w_eco70117, w_eco70118, w_eco70119, w_eco70120, w_eco70121, w_eco70122, w_eco70123, w_eco70124, w_eco70125, w_eco70126, w_eco70127, w_eco70128, w_eco70129, w_eco70130, w_eco70131, w_eco70132, w_eco70133, w_eco70134, w_eco70135, w_eco70136, w_eco70137, w_eco70138, w_eco70139, w_eco70140, w_eco70141, w_eco70142, w_eco70143, w_eco70144, w_eco70145, w_eco70146, w_eco70147, w_eco70148, w_eco70149, w_eco70150, w_eco70151, w_eco70152, w_eco70153, w_eco70154, w_eco70155, w_eco70156, w_eco70157, w_eco70158, w_eco70159, w_eco70160, w_eco70161, w_eco70162, w_eco70163, w_eco70164, w_eco70165, w_eco70166, w_eco70167, w_eco70168, w_eco70169, w_eco70170, w_eco70171, w_eco70172, w_eco70173, w_eco70174, w_eco70175, w_eco70176, w_eco70177, w_eco70178, w_eco70179, w_eco70180, w_eco70181, w_eco70182, w_eco70183, w_eco70184, w_eco70185, w_eco70186, w_eco70187, w_eco70188, w_eco70189, w_eco70190, w_eco70191, w_eco70192, w_eco70193, w_eco70194, w_eco70195, w_eco70196, w_eco70197, w_eco70198, w_eco70199, w_eco70200, w_eco70201, w_eco70202, w_eco70203, w_eco70204, w_eco70205, w_eco70206, w_eco70207, w_eco70208, w_eco70209, w_eco70210, w_eco70211, w_eco70212, w_eco70213, w_eco70214, w_eco70215, w_eco70216, w_eco70217, w_eco70218, w_eco70219, w_eco70220, w_eco70221, w_eco70222, w_eco70223, w_eco70224, w_eco70225, w_eco70226, w_eco70227, w_eco70228, w_eco70229, w_eco70230, w_eco70231, w_eco70232, w_eco70233, w_eco70234, w_eco70235, w_eco70236, w_eco70237, w_eco70238, w_eco70239, w_eco70240, w_eco70241, w_eco70242, w_eco70243, w_eco70244, w_eco70245, w_eco70246, w_eco70247, w_eco70248, w_eco70249, w_eco70250, w_eco70251, w_eco70252, w_eco70253, w_eco70254, w_eco70255, w_eco70256, w_eco70257, w_eco70258, w_eco70259, w_eco70260, w_eco70261, w_eco70262, w_eco70263, w_eco70264, w_eco70265, w_eco70266, w_eco70267, w_eco70268, w_eco70269, w_eco70270, w_eco70271, w_eco70272, w_eco70273, w_eco70274, w_eco70275, w_eco70276, w_eco70277, w_eco70278, w_eco70279, w_eco70280, w_eco70281, w_eco70282, w_eco70283, w_eco70284, w_eco70285, w_eco70286, w_eco70287, w_eco70288, w_eco70289, w_eco70290, w_eco70291, w_eco70292, w_eco70293, w_eco70294, w_eco70295, w_eco70296, w_eco70297, w_eco70298, w_eco70299, w_eco70300, w_eco70301, w_eco70302, w_eco70303, w_eco70304, w_eco70305, w_eco70306, w_eco70307, w_eco70308, w_eco70309, w_eco70310, w_eco70311, w_eco70312, w_eco70313, w_eco70314, w_eco70315, w_eco70316, w_eco70317, w_eco70318, w_eco70319, w_eco70320, w_eco70321, w_eco70322, w_eco70323, w_eco70324, w_eco70325, w_eco70326, w_eco70327, w_eco70328, w_eco70329, w_eco70330, w_eco70331, w_eco70332, w_eco70333, w_eco70334, w_eco70335, w_eco70336, w_eco70337, w_eco70338, w_eco70339, w_eco70340, w_eco70341, w_eco70342, w_eco70343, w_eco70344, w_eco70345, w_eco70346, w_eco70347, w_eco70348, w_eco70349, w_eco70350, w_eco70351, w_eco70352, w_eco70353, w_eco70354, w_eco70355, w_eco70356, w_eco70357, w_eco70358, w_eco70359, w_eco70360, w_eco70361, w_eco70362, w_eco70363, w_eco70364, w_eco70365, w_eco70366, w_eco70367, w_eco70368, w_eco70369, w_eco70370, w_eco70371, w_eco70372, w_eco70373, w_eco70374, w_eco70375, w_eco70376, w_eco70377, w_eco70378, w_eco70379, w_eco70380, w_eco70381, w_eco70382, w_eco70383, w_eco70384, w_eco70385, w_eco70386, w_eco70387, w_eco70388, w_eco70389, w_eco70390, w_eco70391, w_eco70392, w_eco70393, w_eco70394, w_eco70395, w_eco70396, w_eco70397, w_eco70398, w_eco70399, w_eco70400, w_eco70401, w_eco70402, w_eco70403, w_eco70404, w_eco70405, w_eco70406, w_eco70407, w_eco70408, w_eco70409, w_eco70410, w_eco70411, w_eco70412, w_eco70413, w_eco70414, w_eco70415, w_eco70416, w_eco70417, w_eco70418, w_eco70419, w_eco70420, w_eco70421, w_eco70422, w_eco70423, w_eco70424, w_eco70425, w_eco70426, w_eco70427, w_eco70428, w_eco70429, w_eco70430, w_eco70431, w_eco70432, w_eco70433, w_eco70434, w_eco70435, w_eco70436, w_eco70437, w_eco70438, w_eco70439, w_eco70440, w_eco70441, w_eco70442, w_eco70443, w_eco70444, w_eco70445, w_eco70446, w_eco70447, w_eco70448, w_eco70449, w_eco70450, w_eco70451, w_eco70452, w_eco70453, w_eco70454, w_eco70455, w_eco70456, w_eco70457, w_eco70458, w_eco70459, w_eco70460, w_eco70461, w_eco70462, w_eco70463, w_eco70464, w_eco70465, w_eco70466, w_eco70467, w_eco70468, w_eco70469, w_eco70470, w_eco70471, w_eco70472, w_eco70473, w_eco70474, w_eco70475, w_eco70476, w_eco70477, w_eco70478, w_eco70479, w_eco70480, w_eco70481, w_eco70482, w_eco70483, w_eco70484, w_eco70485, w_eco70486, w_eco70487, w_eco70488, w_eco70489, w_eco70490, w_eco70491, w_eco70492, w_eco70493, w_eco70494, w_eco70495, w_eco70496, w_eco70497, w_eco70498, w_eco70499, w_eco70500, w_eco70501, w_eco70502, w_eco70503, w_eco70504, w_eco70505, w_eco70506, w_eco70507, w_eco70508, w_eco70509, w_eco70510, w_eco70511, w_eco70512, w_eco70513, w_eco70514, w_eco70515, w_eco70516, w_eco70517, w_eco70518, w_eco70519, w_eco70520, w_eco70521, w_eco70522, w_eco70523, w_eco70524, w_eco70525, w_eco70526, w_eco70527, w_eco70528, w_eco70529, w_eco70530, w_eco70531, w_eco70532, w_eco70533, w_eco70534, w_eco70535, w_eco70536, w_eco70537, w_eco70538, w_eco70539, w_eco70540, w_eco70541, w_eco70542, w_eco70543, w_eco70544, w_eco70545, w_eco70546, w_eco70547, w_eco70548, w_eco70549, w_eco70550, w_eco70551, w_eco70552, w_eco70553, w_eco70554, w_eco70555, w_eco70556, w_eco70557, w_eco70558, w_eco70559, w_eco70560, w_eco70561, w_eco70562, w_eco70563, w_eco70564, w_eco70565, w_eco70566, w_eco70567, w_eco70568, w_eco70569, w_eco70570, w_eco70571, w_eco70572, w_eco70573, w_eco70574, w_eco70575, w_eco70576, w_eco70577, w_eco70578, w_eco70579, w_eco70580, w_eco70581, w_eco70582, w_eco70583, w_eco70584, w_eco70585, w_eco70586, w_eco70587, w_eco70588, w_eco70589, w_eco70590, w_eco70591, w_eco70592, w_eco70593, w_eco70594, w_eco70595, w_eco70596, w_eco70597, w_eco70598, w_eco70599, w_eco70600, w_eco70601, w_eco70602, w_eco70603, w_eco70604, w_eco70605, w_eco70606, w_eco70607, w_eco70608, w_eco70609, w_eco70610, w_eco70611, w_eco70612, w_eco70613, w_eco70614, w_eco70615, w_eco70616, w_eco70617, w_eco70618, w_eco70619, w_eco70620, w_eco70621, w_eco70622, w_eco70623, w_eco70624, w_eco70625, w_eco70626, w_eco70627, w_eco70628, w_eco70629, w_eco70630, w_eco70631, w_eco70632, w_eco70633, w_eco70634, w_eco70635, w_eco70636, w_eco70637, w_eco70638, w_eco70639, w_eco70640, w_eco70641, w_eco70642, w_eco70643, w_eco70644, w_eco70645, w_eco70646, w_eco70647, w_eco70648, w_eco70649, w_eco70650, w_eco70651, w_eco70652, w_eco70653, w_eco70654, w_eco70655, w_eco70656, w_eco70657, w_eco70658, w_eco70659, w_eco70660, w_eco70661, w_eco70662, w_eco70663, w_eco70664, w_eco70665, w_eco70666, w_eco70667, w_eco70668, w_eco70669, w_eco70670, w_eco70671, w_eco70672, w_eco70673, w_eco70674, w_eco70675, w_eco70676, w_eco70677, w_eco70678, w_eco70679, w_eco70680, w_eco70681, w_eco70682, w_eco70683, w_eco70684, w_eco70685, w_eco70686, w_eco70687, w_eco70688, w_eco70689, w_eco70690, w_eco70691, w_eco70692, w_eco70693, w_eco70694, w_eco70695, w_eco70696, w_eco70697, w_eco70698, w_eco70699, w_eco70700, w_eco70701, w_eco70702, w_eco70703, w_eco70704, w_eco70705, w_eco70706, w_eco70707, w_eco70708, w_eco70709, w_eco70710, w_eco70711, w_eco70712, w_eco70713, w_eco70714, w_eco70715, w_eco70716, w_eco70717, w_eco70718, w_eco70719, w_eco70720, w_eco70721, w_eco70722, w_eco70723, w_eco70724, w_eco70725, w_eco70726, w_eco70727, w_eco70728, w_eco70729, w_eco70730, w_eco70731, w_eco70732, w_eco70733, w_eco70734, w_eco70735, w_eco70736, w_eco70737, w_eco70738, w_eco70739, w_eco70740, w_eco70741, w_eco70742, w_eco70743, w_eco70744, w_eco70745, w_eco70746, w_eco70747, w_eco70748, w_eco70749, w_eco70750, w_eco70751, w_eco70752, w_eco70753, w_eco70754, w_eco70755, w_eco70756, w_eco70757, w_eco70758, w_eco70759, w_eco70760, w_eco70761, w_eco70762, w_eco70763, w_eco70764, w_eco70765, w_eco70766, w_eco70767, w_eco70768, w_eco70769, w_eco70770, w_eco70771, w_eco70772, w_eco70773, w_eco70774, w_eco70775, w_eco70776, w_eco70777, w_eco70778, w_eco70779, w_eco70780, w_eco70781, w_eco70782, w_eco70783, w_eco70784, w_eco70785, w_eco70786, w_eco70787, w_eco70788, w_eco70789, w_eco70790, w_eco70791, w_eco70792, w_eco70793, w_eco70794, w_eco70795, w_eco70796, w_eco70797, w_eco70798, w_eco70799, w_eco70800, w_eco70801, w_eco70802, w_eco70803, w_eco70804, w_eco70805, w_eco70806, w_eco70807, w_eco70808, w_eco70809, w_eco70810, w_eco70811, w_eco70812, w_eco70813, w_eco70814, w_eco70815, w_eco70816, w_eco70817, w_eco70818, w_eco70819, w_eco70820, w_eco70821, w_eco70822, w_eco70823, w_eco70824, w_eco70825, w_eco70826, w_eco70827, w_eco70828, w_eco70829, w_eco70830, w_eco70831, w_eco70832, w_eco70833, w_eco70834, w_eco70835, w_eco70836, w_eco70837, w_eco70838, w_eco70839, w_eco70840, w_eco70841, w_eco70842, w_eco70843, w_eco70844, w_eco70845, w_eco70846, w_eco70847, w_eco70848, w_eco70849, w_eco70850, w_eco70851, w_eco70852, w_eco70853, w_eco70854, w_eco70855, w_eco70856, w_eco70857, w_eco70858, w_eco70859, w_eco70860, w_eco70861, w_eco70862, w_eco70863, w_eco70864, w_eco70865, w_eco70866, w_eco70867, w_eco70868, w_eco70869, w_eco70870, w_eco70871, w_eco70872, w_eco70873, w_eco70874, w_eco70875, w_eco70876, w_eco70877, w_eco70878, w_eco70879, w_eco70880, w_eco70881, w_eco70882, w_eco70883, w_eco70884, w_eco70885, w_eco70886, w_eco70887, w_eco70888, w_eco70889, w_eco70890, w_eco70891, w_eco70892, w_eco70893, w_eco70894, w_eco70895, w_eco70896, w_eco70897, w_eco70898, w_eco70899, w_eco70900, w_eco70901, w_eco70902, w_eco70903, w_eco70904, w_eco70905, w_eco70906, w_eco70907, w_eco70908, w_eco70909, w_eco70910, w_eco70911, w_eco70912, w_eco70913, w_eco70914, w_eco70915, w_eco70916, w_eco70917, w_eco70918, w_eco70919, w_eco70920, w_eco70921, w_eco70922, w_eco70923, w_eco70924, w_eco70925, w_eco70926, w_eco70927, w_eco70928, w_eco70929, w_eco70930, w_eco70931, w_eco70932, w_eco70933, w_eco70934, w_eco70935, w_eco70936, w_eco70937, w_eco70938, w_eco70939, w_eco70940, w_eco70941, w_eco70942, w_eco70943, w_eco70944, w_eco70945, w_eco70946, w_eco70947, w_eco70948, w_eco70949, w_eco70950, w_eco70951, w_eco70952, w_eco70953, w_eco70954, w_eco70955, w_eco70956, w_eco70957, w_eco70958, w_eco70959, w_eco70960, w_eco70961, w_eco70962, w_eco70963, w_eco70964, w_eco70965, w_eco70966, w_eco70967, w_eco70968, w_eco70969, w_eco70970, w_eco70971, w_eco70972, w_eco70973, w_eco70974, w_eco70975, w_eco70976, w_eco70977, w_eco70978, w_eco70979, w_eco70980, w_eco70981, w_eco70982, w_eco70983, w_eco70984, w_eco70985, w_eco70986, w_eco70987, w_eco70988, w_eco70989, w_eco70990, w_eco70991, w_eco70992, w_eco70993, w_eco70994, w_eco70995, w_eco70996, w_eco70997, w_eco70998, w_eco70999, w_eco71000, w_eco71001, w_eco71002, w_eco71003, w_eco71004, w_eco71005, w_eco71006, w_eco71007, w_eco71008, w_eco71009, w_eco71010, w_eco71011, w_eco71012, w_eco71013, w_eco71014, w_eco71015, w_eco71016, w_eco71017, w_eco71018, w_eco71019, w_eco71020, w_eco71021, w_eco71022, w_eco71023, w_eco71024, w_eco71025, w_eco71026, w_eco71027, w_eco71028, w_eco71029, w_eco71030, w_eco71031, w_eco71032, w_eco71033, w_eco71034, w_eco71035, w_eco71036, w_eco71037, w_eco71038, w_eco71039, w_eco71040, w_eco71041, w_eco71042, w_eco71043, w_eco71044, w_eco71045, w_eco71046, w_eco71047, w_eco71048, w_eco71049, w_eco71050, w_eco71051, w_eco71052, w_eco71053, w_eco71054, w_eco71055, w_eco71056, w_eco71057, w_eco71058, w_eco71059, w_eco71060, w_eco71061, w_eco71062, w_eco71063, w_eco71064, w_eco71065, w_eco71066, w_eco71067, w_eco71068, w_eco71069, w_eco71070, w_eco71071, w_eco71072, w_eco71073, w_eco71074, w_eco71075, w_eco71076, w_eco71077, w_eco71078, w_eco71079, w_eco71080, w_eco71081, w_eco71082, w_eco71083, w_eco71084, w_eco71085, w_eco71086, w_eco71087, w_eco71088, w_eco71089, w_eco71090, w_eco71091, w_eco71092, w_eco71093, w_eco71094, w_eco71095, w_eco71096, w_eco71097, w_eco71098, w_eco71099, w_eco71100, w_eco71101, w_eco71102, w_eco71103, w_eco71104, w_eco71105, w_eco71106, w_eco71107, w_eco71108, w_eco71109, w_eco71110, w_eco71111, w_eco71112, w_eco71113, w_eco71114, w_eco71115, w_eco71116, w_eco71117, w_eco71118, w_eco71119, w_eco71120, w_eco71121, w_eco71122, w_eco71123, w_eco71124, w_eco71125, w_eco71126, w_eco71127, w_eco71128, w_eco71129, w_eco71130, w_eco71131, w_eco71132, w_eco71133, w_eco71134, w_eco71135, w_eco71136, w_eco71137, w_eco71138, w_eco71139, w_eco71140, w_eco71141, w_eco71142, w_eco71143, w_eco71144, w_eco71145, w_eco71146, w_eco71147, w_eco71148, w_eco71149, w_eco71150, w_eco71151, w_eco71152, w_eco71153, w_eco71154, w_eco71155, w_eco71156, w_eco71157, w_eco71158, w_eco71159, w_eco71160, w_eco71161, w_eco71162, w_eco71163, w_eco71164, w_eco71165, w_eco71166, w_eco71167, w_eco71168, w_eco71169, w_eco71170, w_eco71171, w_eco71172, w_eco71173, w_eco71174, w_eco71175, w_eco71176, w_eco71177, w_eco71178, w_eco71179, w_eco71180, w_eco71181, w_eco71182, w_eco71183, w_eco71184, w_eco71185, w_eco71186, w_eco71187, w_eco71188, w_eco71189, w_eco71190, w_eco71191, w_eco71192, w_eco71193, w_eco71194, w_eco71195, w_eco71196, w_eco71197, w_eco71198, w_eco71199, w_eco71200, w_eco71201, w_eco71202, w_eco71203, w_eco71204, w_eco71205, w_eco71206, w_eco71207, w_eco71208, w_eco71209, w_eco71210, w_eco71211, w_eco71212, w_eco71213, w_eco71214, w_eco71215, w_eco71216, w_eco71217, w_eco71218, w_eco71219, w_eco71220, w_eco71221, w_eco71222, w_eco71223, w_eco71224, w_eco71225, w_eco71226, w_eco71227, w_eco71228, w_eco71229, w_eco71230, w_eco71231, w_eco71232, w_eco71233, w_eco71234, w_eco71235, w_eco71236, w_eco71237, w_eco71238, w_eco71239, w_eco71240, w_eco71241, w_eco71242, w_eco71243, w_eco71244, w_eco71245, w_eco71246, w_eco71247, w_eco71248, w_eco71249, w_eco71250, w_eco71251, w_eco71252, w_eco71253, w_eco71254, w_eco71255, w_eco71256, w_eco71257, w_eco71258, w_eco71259, w_eco71260, w_eco71261, w_eco71262, w_eco71263, w_eco71264, w_eco71265, w_eco71266, w_eco71267, w_eco71268, w_eco71269, w_eco71270, w_eco71271, w_eco71272, w_eco71273, w_eco71274, w_eco71275, w_eco71276, w_eco71277, w_eco71278, w_eco71279, w_eco71280, w_eco71281, w_eco71282, w_eco71283, w_eco71284, w_eco71285, w_eco71286, w_eco71287, w_eco71288, w_eco71289, w_eco71290, w_eco71291, w_eco71292, w_eco71293, w_eco71294, w_eco71295, w_eco71296, w_eco71297, w_eco71298, w_eco71299, w_eco71300, w_eco71301, w_eco71302, w_eco71303, w_eco71304, w_eco71305, w_eco71306, w_eco71307, w_eco71308, w_eco71309, w_eco71310, w_eco71311, w_eco71312, w_eco71313, w_eco71314, w_eco71315, w_eco71316, w_eco71317, w_eco71318, w_eco71319, w_eco71320, w_eco71321, w_eco71322, w_eco71323, w_eco71324, w_eco71325, w_eco71326, w_eco71327, w_eco71328, w_eco71329, w_eco71330, w_eco71331, w_eco71332, w_eco71333, w_eco71334, w_eco71335, w_eco71336, w_eco71337, w_eco71338, w_eco71339, w_eco71340, w_eco71341, w_eco71342, w_eco71343, w_eco71344, w_eco71345, w_eco71346, w_eco71347, w_eco71348, w_eco71349, w_eco71350, w_eco71351, w_eco71352, w_eco71353, w_eco71354, w_eco71355, w_eco71356, w_eco71357, w_eco71358, w_eco71359, w_eco71360, w_eco71361, w_eco71362, w_eco71363, w_eco71364, w_eco71365, w_eco71366, w_eco71367, w_eco71368, w_eco71369, w_eco71370, w_eco71371, w_eco71372, w_eco71373, w_eco71374, w_eco71375, w_eco71376, w_eco71377, w_eco71378, w_eco71379, w_eco71380, w_eco71381, w_eco71382, w_eco71383, w_eco71384, w_eco71385, w_eco71386, w_eco71387, w_eco71388, w_eco71389, w_eco71390, w_eco71391, w_eco71392, w_eco71393, w_eco71394, w_eco71395, w_eco71396, w_eco71397, w_eco71398, w_eco71399, w_eco71400, w_eco71401, w_eco71402, w_eco71403, w_eco71404, w_eco71405, w_eco71406, w_eco71407, w_eco71408, w_eco71409, w_eco71410, w_eco71411, w_eco71412, w_eco71413, w_eco71414, w_eco71415, w_eco71416, w_eco71417, w_eco71418, w_eco71419, w_eco71420, w_eco71421, w_eco71422, w_eco71423, w_eco71424, w_eco71425, w_eco71426, w_eco71427, w_eco71428, w_eco71429, w_eco71430, w_eco71431, w_eco71432, w_eco71433, w_eco71434, w_eco71435, w_eco71436, w_eco71437, w_eco71438, w_eco71439, w_eco71440, w_eco71441, w_eco71442, w_eco71443, w_eco71444, w_eco71445, w_eco71446, w_eco71447, w_eco71448, w_eco71449, w_eco71450, w_eco71451, w_eco71452, w_eco71453, w_eco71454, w_eco71455, w_eco71456, w_eco71457, w_eco71458, w_eco71459, w_eco71460, w_eco71461, w_eco71462, w_eco71463, w_eco71464, w_eco71465, w_eco71466, w_eco71467, w_eco71468, w_eco71469, w_eco71470, w_eco71471, w_eco71472, w_eco71473, w_eco71474, w_eco71475, w_eco71476, w_eco71477, w_eco71478, w_eco71479, w_eco71480, w_eco71481, w_eco71482, w_eco71483, w_eco71484, w_eco71485, w_eco71486, w_eco71487, w_eco71488, w_eco71489, w_eco71490, w_eco71491, w_eco71492, w_eco71493, w_eco71494, w_eco71495, w_eco71496, w_eco71497, w_eco71498, w_eco71499, w_eco71500, w_eco71501, w_eco71502, w_eco71503, w_eco71504, w_eco71505, w_eco71506, w_eco71507, w_eco71508, w_eco71509, w_eco71510, w_eco71511, w_eco71512, w_eco71513, w_eco71514, w_eco71515, w_eco71516, w_eco71517, w_eco71518, w_eco71519, w_eco71520, w_eco71521, w_eco71522, w_eco71523, w_eco71524, w_eco71525, w_eco71526, w_eco71527, w_eco71528, w_eco71529, w_eco71530, w_eco71531, w_eco71532, w_eco71533, w_eco71534, w_eco71535, w_eco71536, w_eco71537, w_eco71538, w_eco71539, w_eco71540, w_eco71541, w_eco71542, w_eco71543, w_eco71544, w_eco71545, w_eco71546, w_eco71547, w_eco71548, w_eco71549, w_eco71550, w_eco71551, w_eco71552, w_eco71553, w_eco71554, w_eco71555, w_eco71556, w_eco71557, w_eco71558, w_eco71559, w_eco71560, w_eco71561, w_eco71562, w_eco71563, w_eco71564, w_eco71565, w_eco71566, w_eco71567, w_eco71568, w_eco71569, w_eco71570, w_eco71571, w_eco71572, w_eco71573, w_eco71574, w_eco71575, w_eco71576, w_eco71577, w_eco71578, w_eco71579, w_eco71580, w_eco71581, w_eco71582, w_eco71583, w_eco71584, w_eco71585, w_eco71586, w_eco71587, w_eco71588, w_eco71589, w_eco71590, w_eco71591, w_eco71592, w_eco71593, w_eco71594, w_eco71595, w_eco71596, w_eco71597, w_eco71598, w_eco71599, w_eco71600, w_eco71601, w_eco71602, w_eco71603, w_eco71604, w_eco71605, w_eco71606, w_eco71607, w_eco71608, w_eco71609, w_eco71610, w_eco71611, w_eco71612, w_eco71613, w_eco71614, w_eco71615, w_eco71616, w_eco71617, w_eco71618, w_eco71619, w_eco71620, w_eco71621, w_eco71622, w_eco71623, w_eco71624, w_eco71625, w_eco71626, w_eco71627, w_eco71628, w_eco71629, w_eco71630, w_eco71631, w_eco71632, w_eco71633, w_eco71634, w_eco71635, w_eco71636, w_eco71637, w_eco71638, w_eco71639, w_eco71640, w_eco71641, w_eco71642, w_eco71643, w_eco71644, w_eco71645, w_eco71646, w_eco71647, w_eco71648, w_eco71649, w_eco71650, w_eco71651, w_eco71652, w_eco71653, w_eco71654, w_eco71655, w_eco71656, w_eco71657, w_eco71658, w_eco71659, w_eco71660, w_eco71661, w_eco71662, w_eco71663, w_eco71664, w_eco71665, w_eco71666, w_eco71667, w_eco71668, w_eco71669, w_eco71670, w_eco71671, w_eco71672, w_eco71673, w_eco71674, w_eco71675, w_eco71676, w_eco71677, w_eco71678, w_eco71679, w_eco71680, w_eco71681, w_eco71682, w_eco71683, w_eco71684, w_eco71685, w_eco71686, w_eco71687, w_eco71688, w_eco71689, w_eco71690, w_eco71691, w_eco71692, w_eco71693, w_eco71694, w_eco71695, w_eco71696, w_eco71697, w_eco71698, w_eco71699, w_eco71700, w_eco71701, w_eco71702, w_eco71703, w_eco71704, w_eco71705, w_eco71706, w_eco71707, w_eco71708, w_eco71709, w_eco71710, w_eco71711, w_eco71712, w_eco71713, w_eco71714, w_eco71715, w_eco71716, w_eco71717, w_eco71718, w_eco71719, w_eco71720, w_eco71721, w_eco71722, w_eco71723, w_eco71724, w_eco71725, w_eco71726, w_eco71727, w_eco71728, w_eco71729, w_eco71730, w_eco71731, w_eco71732, w_eco71733, w_eco71734, w_eco71735, w_eco71736, w_eco71737, w_eco71738, w_eco71739, w_eco71740, w_eco71741, w_eco71742, w_eco71743, w_eco71744, w_eco71745, w_eco71746, w_eco71747, w_eco71748, w_eco71749, w_eco71750, w_eco71751, w_eco71752, w_eco71753, w_eco71754, w_eco71755, w_eco71756, w_eco71757, w_eco71758, w_eco71759, w_eco71760, w_eco71761, w_eco71762, w_eco71763, w_eco71764, w_eco71765, w_eco71766, w_eco71767, w_eco71768, w_eco71769, w_eco71770, w_eco71771, w_eco71772, w_eco71773, w_eco71774, w_eco71775, w_eco71776, w_eco71777, w_eco71778, w_eco71779, w_eco71780, w_eco71781, w_eco71782, w_eco71783, w_eco71784, w_eco71785, w_eco71786, w_eco71787, w_eco71788, w_eco71789, w_eco71790, w_eco71791, w_eco71792, w_eco71793, w_eco71794, w_eco71795, w_eco71796, w_eco71797, w_eco71798, w_eco71799, w_eco71800, w_eco71801, w_eco71802, w_eco71803, w_eco71804, w_eco71805, w_eco71806, w_eco71807, w_eco71808, w_eco71809, w_eco71810, w_eco71811, w_eco71812, w_eco71813, w_eco71814, w_eco71815, w_eco71816, w_eco71817, w_eco71818, w_eco71819, w_eco71820, w_eco71821, w_eco71822, w_eco71823, w_eco71824, w_eco71825, w_eco71826, w_eco71827, w_eco71828, w_eco71829, w_eco71830, w_eco71831, w_eco71832, w_eco71833, w_eco71834, w_eco71835, w_eco71836, w_eco71837, w_eco71838, w_eco71839, w_eco71840, w_eco71841, w_eco71842, w_eco71843, w_eco71844, w_eco71845, w_eco71846, w_eco71847, w_eco71848, w_eco71849, w_eco71850, w_eco71851, w_eco71852, w_eco71853, w_eco71854, w_eco71855, w_eco71856, w_eco71857, w_eco71858, w_eco71859, w_eco71860, w_eco71861, w_eco71862, w_eco71863, w_eco71864, w_eco71865, w_eco71866, w_eco71867, w_eco71868, w_eco71869, w_eco71870, w_eco71871, w_eco71872, w_eco71873, w_eco71874, w_eco71875, w_eco71876, w_eco71877, w_eco71878, w_eco71879, w_eco71880, w_eco71881, w_eco71882, w_eco71883, w_eco71884, w_eco71885, w_eco71886, w_eco71887, w_eco71888, w_eco71889, w_eco71890, w_eco71891, w_eco71892, w_eco71893, w_eco71894, w_eco71895, w_eco71896, w_eco71897, w_eco71898, w_eco71899, w_eco71900, w_eco71901, w_eco71902, w_eco71903, w_eco71904, w_eco71905, w_eco71906, w_eco71907, w_eco71908, w_eco71909, w_eco71910, w_eco71911, w_eco71912, w_eco71913, w_eco71914, w_eco71915, w_eco71916, w_eco71917, w_eco71918, w_eco71919, w_eco71920, w_eco71921, w_eco71922, w_eco71923, w_eco71924, w_eco71925, w_eco71926, w_eco71927, w_eco71928, w_eco71929, w_eco71930, w_eco71931, w_eco71932, w_eco71933, w_eco71934, w_eco71935, w_eco71936, w_eco71937, w_eco71938, w_eco71939, w_eco71940, w_eco71941, w_eco71942, w_eco71943, w_eco71944, w_eco71945, w_eco71946, w_eco71947, w_eco71948, w_eco71949, w_eco71950, w_eco71951, w_eco71952, w_eco71953, w_eco71954, w_eco71955, w_eco71956, w_eco71957, w_eco71958, w_eco71959, w_eco71960, w_eco71961, w_eco71962, w_eco71963, w_eco71964, w_eco71965, w_eco71966, w_eco71967, w_eco71968, w_eco71969, w_eco71970, w_eco71971, w_eco71972, w_eco71973, w_eco71974, w_eco71975, w_eco71976, w_eco71977, w_eco71978, w_eco71979, w_eco71980, w_eco71981, w_eco71982, w_eco71983, w_eco71984, w_eco71985, w_eco71986, w_eco71987, w_eco71988, w_eco71989, w_eco71990, w_eco71991, w_eco71992, w_eco71993, w_eco71994, w_eco71995, w_eco71996, w_eco71997, w_eco71998, w_eco71999, w_eco72000, w_eco72001, w_eco72002, w_eco72003, w_eco72004, w_eco72005, w_eco72006, w_eco72007, w_eco72008, w_eco72009, w_eco72010, w_eco72011, w_eco72012, w_eco72013, w_eco72014, w_eco72015, w_eco72016, w_eco72017, w_eco72018, w_eco72019, w_eco72020, w_eco72021, w_eco72022, w_eco72023, w_eco72024, w_eco72025, w_eco72026, w_eco72027, w_eco72028, w_eco72029, w_eco72030, w_eco72031, w_eco72032, w_eco72033, w_eco72034, w_eco72035, w_eco72036, w_eco72037, w_eco72038, w_eco72039, w_eco72040, w_eco72041, w_eco72042, w_eco72043, w_eco72044, w_eco72045, w_eco72046, w_eco72047, w_eco72048, w_eco72049, w_eco72050, w_eco72051, w_eco72052, w_eco72053, w_eco72054, w_eco72055, w_eco72056, w_eco72057, w_eco72058, w_eco72059, w_eco72060, w_eco72061, w_eco72062, w_eco72063, w_eco72064, w_eco72065, w_eco72066, w_eco72067, w_eco72068, w_eco72069, w_eco72070, w_eco72071, w_eco72072, w_eco72073, w_eco72074, w_eco72075, w_eco72076, w_eco72077, w_eco72078, w_eco72079, w_eco72080, w_eco72081, w_eco72082, w_eco72083, w_eco72084, w_eco72085, w_eco72086, w_eco72087, w_eco72088, w_eco72089, w_eco72090, w_eco72091, w_eco72092, w_eco72093, w_eco72094, w_eco72095, w_eco72096, w_eco72097, w_eco72098, w_eco72099, w_eco72100, w_eco72101, w_eco72102, w_eco72103, w_eco72104, w_eco72105, w_eco72106, w_eco72107, w_eco72108, w_eco72109, w_eco72110, w_eco72111, w_eco72112, w_eco72113, w_eco72114, w_eco72115, w_eco72116, w_eco72117, w_eco72118, w_eco72119, w_eco72120, w_eco72121, w_eco72122, w_eco72123, w_eco72124, w_eco72125, w_eco72126, w_eco72127, w_eco72128, w_eco72129, w_eco72130, w_eco72131, w_eco72132, w_eco72133, w_eco72134, w_eco72135, w_eco72136, w_eco72137, w_eco72138, w_eco72139, w_eco72140, w_eco72141, w_eco72142, w_eco72143, w_eco72144, w_eco72145, w_eco72146, w_eco72147, w_eco72148, w_eco72149, w_eco72150, w_eco72151, w_eco72152, w_eco72153, w_eco72154, w_eco72155, w_eco72156, w_eco72157, w_eco72158, w_eco72159, w_eco72160, w_eco72161, w_eco72162, w_eco72163, w_eco72164, w_eco72165, w_eco72166, w_eco72167, w_eco72168, w_eco72169, w_eco72170, w_eco72171, w_eco72172, w_eco72173, w_eco72174, w_eco72175, w_eco72176, w_eco72177, w_eco72178, w_eco72179, w_eco72180, w_eco72181, w_eco72182, w_eco72183, w_eco72184, w_eco72185, w_eco72186, w_eco72187, w_eco72188, w_eco72189, w_eco72190, w_eco72191, w_eco72192, w_eco72193, w_eco72194, w_eco72195, w_eco72196, w_eco72197, w_eco72198, w_eco72199, w_eco72200, w_eco72201, w_eco72202, w_eco72203, w_eco72204, w_eco72205, w_eco72206, w_eco72207, w_eco72208, w_eco72209, w_eco72210, w_eco72211, w_eco72212, w_eco72213, w_eco72214, w_eco72215, w_eco72216, w_eco72217, w_eco72218, w_eco72219, w_eco72220, w_eco72221, w_eco72222, w_eco72223, w_eco72224, w_eco72225, w_eco72226, w_eco72227, w_eco72228, w_eco72229, w_eco72230, w_eco72231, w_eco72232, w_eco72233, w_eco72234, w_eco72235, w_eco72236, w_eco72237, w_eco72238, w_eco72239, w_eco72240, w_eco72241, w_eco72242, w_eco72243, w_eco72244, w_eco72245, w_eco72246, w_eco72247, w_eco72248, w_eco72249, w_eco72250, w_eco72251, w_eco72252, w_eco72253, w_eco72254, w_eco72255, w_eco72256, w_eco72257, w_eco72258, w_eco72259, w_eco72260, w_eco72261, w_eco72262, w_eco72263, w_eco72264, w_eco72265, w_eco72266, w_eco72267, w_eco72268, w_eco72269, w_eco72270, w_eco72271, w_eco72272, w_eco72273, w_eco72274, w_eco72275, w_eco72276, w_eco72277, w_eco72278, w_eco72279, w_eco72280, w_eco72281, w_eco72282, w_eco72283, w_eco72284, w_eco72285, w_eco72286, w_eco72287, w_eco72288, w_eco72289, w_eco72290, w_eco72291, w_eco72292, w_eco72293, w_eco72294, w_eco72295, w_eco72296, w_eco72297, w_eco72298, w_eco72299, w_eco72300, w_eco72301, w_eco72302, w_eco72303, w_eco72304, w_eco72305, w_eco72306, w_eco72307, w_eco72308, w_eco72309, w_eco72310, w_eco72311, w_eco72312, w_eco72313, w_eco72314, w_eco72315, w_eco72316, w_eco72317, w_eco72318, w_eco72319, w_eco72320, w_eco72321, w_eco72322, w_eco72323, w_eco72324, w_eco72325, w_eco72326, w_eco72327, w_eco72328, w_eco72329, w_eco72330, w_eco72331, w_eco72332, w_eco72333, w_eco72334, w_eco72335, w_eco72336, w_eco72337, w_eco72338, w_eco72339, w_eco72340, w_eco72341, w_eco72342, w_eco72343, w_eco72344, w_eco72345, w_eco72346, w_eco72347, w_eco72348, w_eco72349, w_eco72350, w_eco72351, w_eco72352, w_eco72353, w_eco72354, w_eco72355, w_eco72356, w_eco72357, w_eco72358, w_eco72359, w_eco72360, w_eco72361, w_eco72362, w_eco72363, w_eco72364, w_eco72365, w_eco72366, w_eco72367, w_eco72368, w_eco72369, w_eco72370, w_eco72371, w_eco72372, w_eco72373, w_eco72374, w_eco72375, w_eco72376, w_eco72377, w_eco72378, w_eco72379, w_eco72380, w_eco72381, w_eco72382, w_eco72383, w_eco72384, w_eco72385, w_eco72386, w_eco72387, w_eco72388, w_eco72389, w_eco72390, w_eco72391, w_eco72392, w_eco72393, w_eco72394, w_eco72395, w_eco72396, w_eco72397, w_eco72398, w_eco72399, w_eco72400, w_eco72401, w_eco72402, w_eco72403, w_eco72404, w_eco72405, w_eco72406, w_eco72407, w_eco72408, w_eco72409, w_eco72410, w_eco72411, w_eco72412, w_eco72413, w_eco72414, w_eco72415, w_eco72416, w_eco72417, w_eco72418, w_eco72419, w_eco72420, w_eco72421, w_eco72422, w_eco72423, w_eco72424, w_eco72425, w_eco72426, w_eco72427, w_eco72428, w_eco72429, w_eco72430, w_eco72431, w_eco72432, w_eco72433, w_eco72434, w_eco72435, w_eco72436, w_eco72437, w_eco72438, w_eco72439, w_eco72440, w_eco72441, w_eco72442, w_eco72443, w_eco72444, w_eco72445, w_eco72446, w_eco72447, w_eco72448, w_eco72449, w_eco72450, w_eco72451, w_eco72452, w_eco72453, w_eco72454, w_eco72455, w_eco72456, w_eco72457, w_eco72458, w_eco72459, w_eco72460, w_eco72461, w_eco72462, w_eco72463, w_eco72464, w_eco72465, w_eco72466, w_eco72467, w_eco72468, w_eco72469, w_eco72470, w_eco72471, w_eco72472, w_eco72473, w_eco72474, w_eco72475, w_eco72476, w_eco72477, w_eco72478, w_eco72479, w_eco72480, w_eco72481, w_eco72482, w_eco72483, w_eco72484, w_eco72485, w_eco72486, w_eco72487, w_eco72488, w_eco72489, w_eco72490, w_eco72491, w_eco72492, w_eco72493, w_eco72494, w_eco72495, w_eco72496, w_eco72497, w_eco72498, w_eco72499, w_eco72500, w_eco72501, w_eco72502, w_eco72503, w_eco72504, w_eco72505, w_eco72506, w_eco72507, w_eco72508, w_eco72509, w_eco72510, w_eco72511, w_eco72512, w_eco72513, w_eco72514, w_eco72515, w_eco72516, w_eco72517, w_eco72518, w_eco72519, w_eco72520, w_eco72521, w_eco72522, w_eco72523, w_eco72524, w_eco72525, w_eco72526, w_eco72527, w_eco72528, w_eco72529, w_eco72530, w_eco72531, w_eco72532, w_eco72533, w_eco72534, w_eco72535, w_eco72536, w_eco72537, w_eco72538, w_eco72539, w_eco72540, w_eco72541, w_eco72542, w_eco72543, w_eco72544, w_eco72545, w_eco72546, w_eco72547, w_eco72548, w_eco72549, w_eco72550, w_eco72551, w_eco72552, w_eco72553, w_eco72554, w_eco72555, w_eco72556, w_eco72557, w_eco72558, w_eco72559, w_eco72560, w_eco72561, w_eco72562, w_eco72563, w_eco72564, w_eco72565, w_eco72566, w_eco72567, w_eco72568, w_eco72569, w_eco72570, w_eco72571, w_eco72572, w_eco72573, w_eco72574, w_eco72575, w_eco72576, w_eco72577, w_eco72578, w_eco72579, w_eco72580, w_eco72581, w_eco72582, w_eco72583, w_eco72584, w_eco72585, w_eco72586, w_eco72587, w_eco72588, w_eco72589, w_eco72590, w_eco72591, w_eco72592, w_eco72593, w_eco72594, w_eco72595, w_eco72596, w_eco72597, w_eco72598, w_eco72599, w_eco72600, w_eco72601, w_eco72602, w_eco72603, w_eco72604, w_eco72605, w_eco72606, w_eco72607, w_eco72608, w_eco72609, w_eco72610, w_eco72611, w_eco72612, w_eco72613, w_eco72614, w_eco72615, w_eco72616, w_eco72617, w_eco72618, w_eco72619, w_eco72620, w_eco72621, w_eco72622, w_eco72623, w_eco72624, w_eco72625, w_eco72626, w_eco72627, w_eco72628, w_eco72629, w_eco72630, w_eco72631, w_eco72632, w_eco72633, w_eco72634, w_eco72635, w_eco72636, w_eco72637, w_eco72638, w_eco72639, w_eco72640, w_eco72641, w_eco72642, w_eco72643, w_eco72644, w_eco72645, w_eco72646, w_eco72647, w_eco72648, w_eco72649, w_eco72650, w_eco72651, w_eco72652, w_eco72653, w_eco72654, w_eco72655, w_eco72656, w_eco72657, w_eco72658, w_eco72659, w_eco72660, w_eco72661, w_eco72662, w_eco72663, w_eco72664, w_eco72665, w_eco72666, w_eco72667, w_eco72668, w_eco72669, w_eco72670, w_eco72671, w_eco72672, w_eco72673, w_eco72674, w_eco72675, w_eco72676, w_eco72677, w_eco72678, w_eco72679, w_eco72680, w_eco72681, w_eco72682, w_eco72683, w_eco72684, w_eco72685, w_eco72686, w_eco72687, w_eco72688, w_eco72689, w_eco72690, w_eco72691, w_eco72692, w_eco72693, w_eco72694, w_eco72695, w_eco72696, w_eco72697, w_eco72698, w_eco72699, w_eco72700, w_eco72701, w_eco72702, w_eco72703, w_eco72704, w_eco72705, w_eco72706, w_eco72707, w_eco72708, w_eco72709, w_eco72710, w_eco72711, w_eco72712, w_eco72713, w_eco72714, w_eco72715, w_eco72716, w_eco72717, w_eco72718, w_eco72719, w_eco72720, w_eco72721, w_eco72722, w_eco72723, w_eco72724, w_eco72725, w_eco72726, w_eco72727, w_eco72728, w_eco72729, w_eco72730, w_eco72731, w_eco72732, w_eco72733, w_eco72734, w_eco72735, w_eco72736, w_eco72737, w_eco72738, w_eco72739, w_eco72740, w_eco72741, w_eco72742, w_eco72743, w_eco72744, w_eco72745, w_eco72746, w_eco72747, w_eco72748, w_eco72749, w_eco72750, w_eco72751, w_eco72752, w_eco72753, w_eco72754, w_eco72755, w_eco72756, w_eco72757, w_eco72758, w_eco72759, w_eco72760, w_eco72761, w_eco72762, w_eco72763, w_eco72764, w_eco72765, w_eco72766, w_eco72767, w_eco72768, w_eco72769, w_eco72770, w_eco72771, w_eco72772, w_eco72773, w_eco72774, w_eco72775, w_eco72776, w_eco72777, w_eco72778, w_eco72779, w_eco72780, w_eco72781, w_eco72782, w_eco72783, w_eco72784, w_eco72785, w_eco72786, w_eco72787, w_eco72788, w_eco72789, w_eco72790, w_eco72791, w_eco72792, w_eco72793, w_eco72794, w_eco72795, w_eco72796, w_eco72797, w_eco72798, w_eco72799, w_eco72800, w_eco72801, w_eco72802, w_eco72803, w_eco72804, w_eco72805, w_eco72806, w_eco72807, w_eco72808, w_eco72809, w_eco72810, w_eco72811, w_eco72812, w_eco72813, w_eco72814, w_eco72815, w_eco72816, w_eco72817, w_eco72818, w_eco72819, w_eco72820, w_eco72821, w_eco72822, w_eco72823, w_eco72824, w_eco72825, w_eco72826, w_eco72827, w_eco72828, w_eco72829, w_eco72830, w_eco72831, w_eco72832, w_eco72833, w_eco72834, w_eco72835, w_eco72836, w_eco72837, w_eco72838, w_eco72839, w_eco72840, w_eco72841, w_eco72842, w_eco72843, w_eco72844, w_eco72845, w_eco72846, w_eco72847, w_eco72848, w_eco72849, w_eco72850, w_eco72851, w_eco72852, w_eco72853, w_eco72854, w_eco72855, w_eco72856, w_eco72857, w_eco72858, w_eco72859, w_eco72860, w_eco72861, w_eco72862, w_eco72863, w_eco72864, w_eco72865, w_eco72866, w_eco72867, w_eco72868, w_eco72869, w_eco72870, w_eco72871, w_eco72872, w_eco72873, w_eco72874, w_eco72875, w_eco72876, w_eco72877, w_eco72878, w_eco72879, w_eco72880, w_eco72881, w_eco72882, w_eco72883, w_eco72884, w_eco72885, w_eco72886, w_eco72887, w_eco72888, w_eco72889, w_eco72890, w_eco72891, w_eco72892, w_eco72893, w_eco72894, w_eco72895, w_eco72896, w_eco72897, w_eco72898, w_eco72899, w_eco72900, w_eco72901, w_eco72902, w_eco72903, w_eco72904, w_eco72905, w_eco72906, w_eco72907, w_eco72908, w_eco72909, w_eco72910, w_eco72911, w_eco72912, w_eco72913, w_eco72914, w_eco72915, w_eco72916, w_eco72917, w_eco72918, w_eco72919, w_eco72920, w_eco72921, w_eco72922, w_eco72923, w_eco72924, w_eco72925, w_eco72926, w_eco72927, w_eco72928, w_eco72929, w_eco72930, w_eco72931, w_eco72932, w_eco72933, w_eco72934, w_eco72935, w_eco72936, w_eco72937, w_eco72938, w_eco72939, w_eco72940, w_eco72941, w_eco72942, w_eco72943, w_eco72944, w_eco72945, w_eco72946, w_eco72947, w_eco72948, w_eco72949, w_eco72950, w_eco72951, w_eco72952, w_eco72953, w_eco72954, w_eco72955, w_eco72956, w_eco72957, w_eco72958, w_eco72959, w_eco72960, w_eco72961, w_eco72962, w_eco72963, w_eco72964, w_eco72965, w_eco72966, w_eco72967, w_eco72968, w_eco72969, w_eco72970, w_eco72971, w_eco72972, w_eco72973, w_eco72974, w_eco72975, w_eco72976, w_eco72977, w_eco72978, w_eco72979, w_eco72980, w_eco72981, w_eco72982, w_eco72983, w_eco72984, w_eco72985, w_eco72986, w_eco72987, w_eco72988, w_eco72989, w_eco72990, w_eco72991, w_eco72992, w_eco72993, w_eco72994, w_eco72995, w_eco72996, w_eco72997, w_eco72998, w_eco72999, w_eco73000, w_eco73001, w_eco73002, w_eco73003, w_eco73004, w_eco73005, w_eco73006, w_eco73007, w_eco73008, w_eco73009, w_eco73010, w_eco73011, w_eco73012, w_eco73013, w_eco73014, w_eco73015, w_eco73016, w_eco73017, w_eco73018, w_eco73019, w_eco73020, w_eco73021, w_eco73022, w_eco73023, w_eco73024, w_eco73025, w_eco73026, w_eco73027, w_eco73028, w_eco73029, w_eco73030, w_eco73031, w_eco73032, w_eco73033, w_eco73034, w_eco73035, w_eco73036, w_eco73037, w_eco73038, w_eco73039, w_eco73040, w_eco73041, w_eco73042, w_eco73043, w_eco73044, w_eco73045, w_eco73046, w_eco73047, w_eco73048, w_eco73049, w_eco73050, w_eco73051, w_eco73052, w_eco73053, w_eco73054, w_eco73055, w_eco73056, w_eco73057, w_eco73058, w_eco73059, w_eco73060, w_eco73061, w_eco73062, w_eco73063, w_eco73064, w_eco73065, w_eco73066, w_eco73067, w_eco73068, w_eco73069, w_eco73070, w_eco73071, w_eco73072, w_eco73073, w_eco73074, w_eco73075, w_eco73076, w_eco73077, w_eco73078, w_eco73079, w_eco73080, w_eco73081, w_eco73082, w_eco73083, w_eco73084, w_eco73085, w_eco73086, w_eco73087, w_eco73088, w_eco73089, w_eco73090, w_eco73091, w_eco73092, w_eco73093, w_eco73094, w_eco73095, w_eco73096, w_eco73097, w_eco73098, w_eco73099, w_eco73100, w_eco73101, w_eco73102, w_eco73103, w_eco73104, w_eco73105, w_eco73106, w_eco73107, w_eco73108, w_eco73109, w_eco73110, w_eco73111, w_eco73112, w_eco73113, w_eco73114, w_eco73115, w_eco73116, w_eco73117, w_eco73118, w_eco73119, w_eco73120, w_eco73121, w_eco73122, w_eco73123, w_eco73124, w_eco73125, w_eco73126, w_eco73127, w_eco73128, w_eco73129, w_eco73130, w_eco73131, w_eco73132, w_eco73133, w_eco73134, w_eco73135, w_eco73136, w_eco73137, w_eco73138, w_eco73139, w_eco73140, w_eco73141, w_eco73142, w_eco73143, w_eco73144, w_eco73145, w_eco73146, w_eco73147, w_eco73148, w_eco73149, w_eco73150, w_eco73151, w_eco73152, w_eco73153, w_eco73154, w_eco73155, w_eco73156, w_eco73157, w_eco73158, w_eco73159, w_eco73160, w_eco73161, w_eco73162, w_eco73163, w_eco73164, w_eco73165, w_eco73166, w_eco73167, w_eco73168, w_eco73169, w_eco73170, w_eco73171, w_eco73172, w_eco73173, w_eco73174, w_eco73175, w_eco73176, w_eco73177, w_eco73178, w_eco73179, w_eco73180, w_eco73181, w_eco73182, w_eco73183, w_eco73184, w_eco73185, w_eco73186, w_eco73187, w_eco73188, w_eco73189, w_eco73190, w_eco73191, w_eco73192, w_eco73193, w_eco73194, w_eco73195, w_eco73196, w_eco73197, w_eco73198, w_eco73199, w_eco73200, w_eco73201, w_eco73202, w_eco73203, w_eco73204, w_eco73205, w_eco73206, w_eco73207, w_eco73208, w_eco73209, w_eco73210, w_eco73211, w_eco73212, w_eco73213, w_eco73214, w_eco73215, w_eco73216, w_eco73217, w_eco73218, w_eco73219, w_eco73220, w_eco73221, w_eco73222, w_eco73223, w_eco73224, w_eco73225, w_eco73226, w_eco73227, w_eco73228, w_eco73229, w_eco73230, w_eco73231, w_eco73232, w_eco73233, w_eco73234, w_eco73235, w_eco73236, w_eco73237, w_eco73238, w_eco73239, w_eco73240, w_eco73241, w_eco73242, w_eco73243, w_eco73244, w_eco73245, w_eco73246, w_eco73247, w_eco73248, w_eco73249, w_eco73250, w_eco73251, w_eco73252, w_eco73253, w_eco73254, w_eco73255, w_eco73256, w_eco73257, w_eco73258, w_eco73259, w_eco73260, w_eco73261, w_eco73262, w_eco73263, w_eco73264, w_eco73265, w_eco73266, w_eco73267, w_eco73268, w_eco73269, w_eco73270, w_eco73271, w_eco73272, w_eco73273, w_eco73274, w_eco73275, w_eco73276, w_eco73277, w_eco73278, w_eco73279, w_eco73280, w_eco73281, w_eco73282, w_eco73283, w_eco73284, w_eco73285, w_eco73286, w_eco73287, w_eco73288, w_eco73289, w_eco73290, w_eco73291, w_eco73292, w_eco73293, w_eco73294, w_eco73295, w_eco73296, w_eco73297, w_eco73298, w_eco73299, w_eco73300, w_eco73301, w_eco73302, w_eco73303, w_eco73304, w_eco73305, w_eco73306, w_eco73307, w_eco73308, w_eco73309, w_eco73310, w_eco73311, w_eco73312, w_eco73313, w_eco73314, w_eco73315, w_eco73316, w_eco73317, w_eco73318, w_eco73319, w_eco73320, w_eco73321, w_eco73322, w_eco73323, w_eco73324, w_eco73325, w_eco73326, w_eco73327, w_eco73328, w_eco73329, w_eco73330, w_eco73331, w_eco73332, w_eco73333, w_eco73334, w_eco73335, w_eco73336, w_eco73337, w_eco73338, w_eco73339, w_eco73340, w_eco73341, w_eco73342, w_eco73343, w_eco73344, w_eco73345, w_eco73346, w_eco73347, w_eco73348, w_eco73349, w_eco73350, w_eco73351, w_eco73352, w_eco73353, w_eco73354, w_eco73355, w_eco73356, w_eco73357, w_eco73358, w_eco73359, w_eco73360, w_eco73361, w_eco73362, w_eco73363, w_eco73364, w_eco73365, w_eco73366, w_eco73367, w_eco73368, w_eco73369, w_eco73370, w_eco73371, w_eco73372, w_eco73373, w_eco73374, w_eco73375, w_eco73376, w_eco73377, w_eco73378, w_eco73379, w_eco73380, w_eco73381, w_eco73382, w_eco73383, w_eco73384, w_eco73385, w_eco73386, w_eco73387, w_eco73388, w_eco73389, w_eco73390, w_eco73391, w_eco73392, w_eco73393, w_eco73394, w_eco73395, w_eco73396, w_eco73397, w_eco73398, w_eco73399, w_eco73400, w_eco73401, w_eco73402, w_eco73403, w_eco73404, w_eco73405, w_eco73406, w_eco73407, w_eco73408, w_eco73409, w_eco73410, w_eco73411, w_eco73412, w_eco73413, w_eco73414, w_eco73415, w_eco73416, w_eco73417, w_eco73418, w_eco73419, w_eco73420, w_eco73421, w_eco73422, w_eco73423, w_eco73424, w_eco73425, w_eco73426, w_eco73427, w_eco73428, w_eco73429, w_eco73430, w_eco73431, w_eco73432, w_eco73433, w_eco73434, w_eco73435, w_eco73436, w_eco73437, w_eco73438, w_eco73439, w_eco73440, w_eco73441, w_eco73442, w_eco73443, w_eco73444, w_eco73445, w_eco73446, w_eco73447, w_eco73448, w_eco73449, w_eco73450, w_eco73451, w_eco73452, w_eco73453, w_eco73454, w_eco73455, w_eco73456, w_eco73457, w_eco73458, w_eco73459, w_eco73460, w_eco73461, w_eco73462, w_eco73463, w_eco73464, w_eco73465, w_eco73466, w_eco73467, w_eco73468, w_eco73469, w_eco73470, w_eco73471, w_eco73472, w_eco73473, w_eco73474, w_eco73475, w_eco73476, w_eco73477, w_eco73478, w_eco73479, w_eco73480, w_eco73481, w_eco73482, w_eco73483, w_eco73484, w_eco73485, w_eco73486, w_eco73487, w_eco73488, w_eco73489, w_eco73490, w_eco73491, w_eco73492, w_eco73493, w_eco73494, w_eco73495, w_eco73496, w_eco73497, w_eco73498, w_eco73499, w_eco73500, w_eco73501, w_eco73502, w_eco73503, w_eco73504, w_eco73505, w_eco73506, w_eco73507, w_eco73508, w_eco73509, w_eco73510, w_eco73511, w_eco73512, w_eco73513, w_eco73514, w_eco73515, w_eco73516, w_eco73517, w_eco73518, w_eco73519, w_eco73520, w_eco73521, w_eco73522, w_eco73523, w_eco73524, w_eco73525, w_eco73526, w_eco73527, w_eco73528, w_eco73529, w_eco73530, w_eco73531, w_eco73532, w_eco73533, w_eco73534, w_eco73535, w_eco73536, w_eco73537, w_eco73538, w_eco73539, w_eco73540, w_eco73541, w_eco73542, w_eco73543, w_eco73544, w_eco73545, w_eco73546, w_eco73547, w_eco73548, w_eco73549, w_eco73550, w_eco73551, w_eco73552, w_eco73553, w_eco73554, w_eco73555, w_eco73556, w_eco73557, w_eco73558, w_eco73559, w_eco73560, w_eco73561, w_eco73562, w_eco73563, w_eco73564, w_eco73565, w_eco73566, w_eco73567, w_eco73568, w_eco73569, w_eco73570, w_eco73571, w_eco73572, w_eco73573, w_eco73574, w_eco73575, w_eco73576, w_eco73577, w_eco73578, w_eco73579, w_eco73580, w_eco73581, w_eco73582, w_eco73583, w_eco73584, w_eco73585, w_eco73586, w_eco73587, w_eco73588, w_eco73589, w_eco73590, w_eco73591, w_eco73592, w_eco73593, w_eco73594, w_eco73595, w_eco73596, w_eco73597, w_eco73598, w_eco73599, w_eco73600, w_eco73601, w_eco73602, w_eco73603, w_eco73604, w_eco73605, w_eco73606, w_eco73607, w_eco73608, w_eco73609, w_eco73610, w_eco73611, w_eco73612, w_eco73613, w_eco73614, w_eco73615, w_eco73616, w_eco73617, w_eco73618, w_eco73619, w_eco73620, w_eco73621, w_eco73622, w_eco73623, w_eco73624, w_eco73625, w_eco73626, w_eco73627, w_eco73628, w_eco73629, w_eco73630, w_eco73631, w_eco73632, w_eco73633, w_eco73634, w_eco73635, w_eco73636, w_eco73637, w_eco73638, w_eco73639, w_eco73640, w_eco73641, w_eco73642, w_eco73643, w_eco73644, w_eco73645, w_eco73646, w_eco73647, w_eco73648, w_eco73649, w_eco73650, w_eco73651, w_eco73652, w_eco73653, w_eco73654, w_eco73655, w_eco73656, w_eco73657, w_eco73658, w_eco73659, w_eco73660, w_eco73661, w_eco73662, w_eco73663, w_eco73664, w_eco73665, w_eco73666, w_eco73667, w_eco73668, w_eco73669, w_eco73670, w_eco73671, w_eco73672, w_eco73673, w_eco73674, w_eco73675, w_eco73676, w_eco73677, w_eco73678, w_eco73679, w_eco73680, w_eco73681, w_eco73682, w_eco73683, w_eco73684, w_eco73685, w_eco73686, w_eco73687, w_eco73688, w_eco73689, w_eco73690, w_eco73691, w_eco73692, w_eco73693, w_eco73694, w_eco73695, w_eco73696, w_eco73697, w_eco73698, w_eco73699, w_eco73700, w_eco73701, w_eco73702, w_eco73703, w_eco73704, w_eco73705, w_eco73706, w_eco73707, w_eco73708, w_eco73709, w_eco73710, w_eco73711, w_eco73712, w_eco73713, w_eco73714, w_eco73715, w_eco73716, w_eco73717, w_eco73718, w_eco73719, w_eco73720, w_eco73721, w_eco73722, w_eco73723, w_eco73724, w_eco73725, w_eco73726, w_eco73727, w_eco73728, w_eco73729, w_eco73730, w_eco73731, w_eco73732, w_eco73733, w_eco73734, w_eco73735, w_eco73736, w_eco73737, w_eco73738, w_eco73739, w_eco73740, w_eco73741, w_eco73742, w_eco73743, w_eco73744, w_eco73745, w_eco73746, w_eco73747, w_eco73748, w_eco73749, w_eco73750, w_eco73751, w_eco73752, w_eco73753, w_eco73754, w_eco73755, w_eco73756, w_eco73757, w_eco73758, w_eco73759, w_eco73760, w_eco73761, w_eco73762, w_eco73763, w_eco73764, w_eco73765, w_eco73766, w_eco73767, w_eco73768, w_eco73769, w_eco73770, w_eco73771, w_eco73772, w_eco73773, w_eco73774, w_eco73775, w_eco73776, w_eco73777, w_eco73778, w_eco73779, w_eco73780, w_eco73781, w_eco73782, w_eco73783, w_eco73784, w_eco73785, w_eco73786, w_eco73787, w_eco73788, w_eco73789, w_eco73790, w_eco73791, w_eco73792, w_eco73793, w_eco73794, w_eco73795, w_eco73796, w_eco73797, w_eco73798, w_eco73799, w_eco73800, w_eco73801, w_eco73802, w_eco73803, w_eco73804, w_eco73805, w_eco73806, w_eco73807, w_eco73808, w_eco73809, w_eco73810, w_eco73811, w_eco73812, w_eco73813, w_eco73814, w_eco73815, w_eco73816, w_eco73817, w_eco73818, w_eco73819, w_eco73820, w_eco73821, w_eco73822, w_eco73823, w_eco73824, w_eco73825, w_eco73826, w_eco73827, w_eco73828, w_eco73829, w_eco73830, w_eco73831, w_eco73832, w_eco73833, w_eco73834, w_eco73835, w_eco73836, w_eco73837, w_eco73838, w_eco73839, w_eco73840, w_eco73841, w_eco73842, w_eco73843, w_eco73844, w_eco73845, w_eco73846, w_eco73847, w_eco73848, w_eco73849, w_eco73850, w_eco73851, w_eco73852, w_eco73853, w_eco73854, w_eco73855, w_eco73856, w_eco73857, w_eco73858, w_eco73859, w_eco73860, w_eco73861, w_eco73862, w_eco73863, w_eco73864, w_eco73865, w_eco73866, w_eco73867, w_eco73868, w_eco73869, w_eco73870, w_eco73871, w_eco73872, w_eco73873, w_eco73874, w_eco73875, w_eco73876, w_eco73877, w_eco73878, w_eco73879, w_eco73880, w_eco73881, w_eco73882, w_eco73883, w_eco73884, w_eco73885, w_eco73886, w_eco73887, w_eco73888, w_eco73889, w_eco73890, w_eco73891, w_eco73892, w_eco73893, w_eco73894, w_eco73895, w_eco73896, w_eco73897, w_eco73898, w_eco73899, w_eco73900, w_eco73901, w_eco73902, w_eco73903, w_eco73904, w_eco73905, w_eco73906, w_eco73907, w_eco73908, w_eco73909, w_eco73910, w_eco73911, w_eco73912, w_eco73913, w_eco73914, w_eco73915, w_eco73916, w_eco73917, w_eco73918, w_eco73919, w_eco73920, w_eco73921, w_eco73922, w_eco73923, w_eco73924, w_eco73925, w_eco73926, w_eco73927, w_eco73928, w_eco73929, w_eco73930, w_eco73931, w_eco73932, w_eco73933, w_eco73934, w_eco73935, w_eco73936, w_eco73937, w_eco73938, w_eco73939, w_eco73940, w_eco73941, w_eco73942, w_eco73943, w_eco73944, w_eco73945, w_eco73946, w_eco73947, w_eco73948, w_eco73949, w_eco73950, w_eco73951, w_eco73952, w_eco73953, w_eco73954, w_eco73955, w_eco73956, w_eco73957, w_eco73958, w_eco73959, w_eco73960, w_eco73961, w_eco73962, w_eco73963, w_eco73964, w_eco73965, w_eco73966, w_eco73967, w_eco73968, w_eco73969, w_eco73970, w_eco73971, w_eco73972, w_eco73973, w_eco73974, w_eco73975, w_eco73976, w_eco73977, w_eco73978, w_eco73979, w_eco73980, w_eco73981, w_eco73982, w_eco73983, w_eco73984, w_eco73985, w_eco73986, w_eco73987, w_eco73988, w_eco73989, w_eco73990, w_eco73991, w_eco73992, w_eco73993, w_eco73994, w_eco73995, w_eco73996, w_eco73997, w_eco73998, w_eco73999, w_eco74000, w_eco74001, w_eco74002, w_eco74003, w_eco74004, w_eco74005, w_eco74006, w_eco74007, w_eco74008, w_eco74009, w_eco74010, w_eco74011, w_eco74012, w_eco74013, w_eco74014, w_eco74015, w_eco74016, w_eco74017, w_eco74018, w_eco74019, w_eco74020, w_eco74021, w_eco74022, w_eco74023, w_eco74024, w_eco74025, w_eco74026, w_eco74027, w_eco74028, w_eco74029, w_eco74030, w_eco74031, w_eco74032, w_eco74033, w_eco74034, w_eco74035, w_eco74036, w_eco74037, w_eco74038, w_eco74039, w_eco74040, w_eco74041, w_eco74042, w_eco74043, w_eco74044, w_eco74045, w_eco74046, w_eco74047, w_eco74048, w_eco74049, w_eco74050, w_eco74051, w_eco74052, w_eco74053, w_eco74054, w_eco74055, w_eco74056, w_eco74057, w_eco74058, w_eco74059, w_eco74060, w_eco74061, w_eco74062, w_eco74063, w_eco74064, w_eco74065, w_eco74066, w_eco74067, w_eco74068, w_eco74069, w_eco74070, w_eco74071, w_eco74072, w_eco74073, w_eco74074, w_eco74075, w_eco74076, w_eco74077, w_eco74078, w_eco74079, w_eco74080, w_eco74081, w_eco74082, w_eco74083, w_eco74084, w_eco74085, w_eco74086, w_eco74087, w_eco74088, w_eco74089, w_eco74090, w_eco74091, w_eco74092, w_eco74093, w_eco74094, w_eco74095, w_eco74096, w_eco74097, w_eco74098, w_eco74099, w_eco74100, w_eco74101, w_eco74102, w_eco74103, w_eco74104, w_eco74105, w_eco74106, w_eco74107, w_eco74108, w_eco74109, w_eco74110, w_eco74111, w_eco74112, w_eco74113, w_eco74114, w_eco74115, w_eco74116, w_eco74117, w_eco74118, w_eco74119, w_eco74120, w_eco74121, w_eco74122, w_eco74123, w_eco74124, w_eco74125, w_eco74126, w_eco74127, w_eco74128, w_eco74129, w_eco74130, w_eco74131, w_eco74132, w_eco74133, w_eco74134, w_eco74135, w_eco74136, w_eco74137, w_eco74138, w_eco74139, w_eco74140, w_eco74141, w_eco74142, w_eco74143, w_eco74144, w_eco74145, w_eco74146, w_eco74147, w_eco74148, w_eco74149, w_eco74150, w_eco74151, w_eco74152, w_eco74153, w_eco74154, w_eco74155, w_eco74156, w_eco74157, w_eco74158, w_eco74159, w_eco74160, w_eco74161, w_eco74162, w_eco74163, w_eco74164, w_eco74165, w_eco74166, w_eco74167, w_eco74168, w_eco74169, w_eco74170, w_eco74171, w_eco74172, w_eco74173, w_eco74174, w_eco74175, w_eco74176, w_eco74177, w_eco74178, w_eco74179, w_eco74180, w_eco74181, w_eco74182, w_eco74183, w_eco74184, w_eco74185, w_eco74186, w_eco74187, w_eco74188, w_eco74189, w_eco74190, w_eco74191, w_eco74192, w_eco74193, w_eco74194, w_eco74195, w_eco74196, w_eco74197, w_eco74198, w_eco74199, w_eco74200, w_eco74201, w_eco74202, w_eco74203, w_eco74204, w_eco74205, w_eco74206, w_eco74207, w_eco74208, w_eco74209, w_eco74210, w_eco74211, w_eco74212, w_eco74213, w_eco74214, w_eco74215, w_eco74216, w_eco74217, w_eco74218, w_eco74219, w_eco74220, w_eco74221, w_eco74222, w_eco74223, w_eco74224, w_eco74225, w_eco74226, w_eco74227, w_eco74228, w_eco74229, w_eco74230, w_eco74231, w_eco74232, w_eco74233, w_eco74234, w_eco74235, w_eco74236, w_eco74237, w_eco74238, w_eco74239, w_eco74240, w_eco74241, w_eco74242, w_eco74243, w_eco74244, w_eco74245, w_eco74246, w_eco74247, w_eco74248, w_eco74249, w_eco74250, w_eco74251, w_eco74252, w_eco74253, w_eco74254, w_eco74255, w_eco74256, w_eco74257, w_eco74258, w_eco74259, w_eco74260, w_eco74261, w_eco74262, w_eco74263, w_eco74264, w_eco74265, w_eco74266, w_eco74267, w_eco74268, w_eco74269, w_eco74270, w_eco74271, w_eco74272, w_eco74273, w_eco74274, w_eco74275, w_eco74276, w_eco74277, w_eco74278, w_eco74279, w_eco74280, w_eco74281, w_eco74282, w_eco74283, w_eco74284, w_eco74285, w_eco74286, w_eco74287, w_eco74288, w_eco74289, w_eco74290, w_eco74291, w_eco74292, w_eco74293, w_eco74294, w_eco74295, w_eco74296, w_eco74297, w_eco74298, w_eco74299, w_eco74300, w_eco74301, w_eco74302, w_eco74303, w_eco74304, w_eco74305, w_eco74306, w_eco74307, w_eco74308, w_eco74309, w_eco74310, w_eco74311, w_eco74312, w_eco74313, w_eco74314, w_eco74315, w_eco74316, w_eco74317, w_eco74318, w_eco74319, w_eco74320, w_eco74321, w_eco74322, w_eco74323, w_eco74324, w_eco74325, w_eco74326, w_eco74327, w_eco74328, w_eco74329, w_eco74330, w_eco74331, w_eco74332, w_eco74333, w_eco74334, w_eco74335, w_eco74336, w_eco74337, w_eco74338, w_eco74339, w_eco74340, w_eco74341, w_eco74342, w_eco74343, w_eco74344, w_eco74345, w_eco74346, w_eco74347, w_eco74348, w_eco74349, w_eco74350, w_eco74351, w_eco74352, w_eco74353, w_eco74354, w_eco74355, w_eco74356, w_eco74357, w_eco74358, w_eco74359, w_eco74360, w_eco74361, w_eco74362, w_eco74363, w_eco74364, w_eco74365, w_eco74366, w_eco74367, w_eco74368, w_eco74369, w_eco74370, w_eco74371, w_eco74372, w_eco74373, w_eco74374, w_eco74375, w_eco74376, w_eco74377, w_eco74378, w_eco74379, w_eco74380, w_eco74381, w_eco74382, w_eco74383, w_eco74384, w_eco74385, w_eco74386, w_eco74387, w_eco74388, w_eco74389, w_eco74390, w_eco74391, w_eco74392, w_eco74393, w_eco74394, w_eco74395, w_eco74396, w_eco74397, w_eco74398, w_eco74399, w_eco74400, w_eco74401, w_eco74402, w_eco74403, w_eco74404, w_eco74405, w_eco74406, w_eco74407, w_eco74408, w_eco74409, w_eco74410, w_eco74411, w_eco74412, w_eco74413, w_eco74414, w_eco74415, w_eco74416, w_eco74417, w_eco74418, w_eco74419, w_eco74420, w_eco74421, w_eco74422, w_eco74423, w_eco74424, w_eco74425, w_eco74426, w_eco74427, w_eco74428, w_eco74429, w_eco74430, w_eco74431, w_eco74432, w_eco74433, w_eco74434, w_eco74435, w_eco74436, w_eco74437, w_eco74438, w_eco74439, w_eco74440, w_eco74441, w_eco74442, w_eco74443, w_eco74444, w_eco74445, w_eco74446, w_eco74447, w_eco74448, w_eco74449, w_eco74450, w_eco74451, w_eco74452, w_eco74453, w_eco74454, w_eco74455, w_eco74456, w_eco74457, w_eco74458, w_eco74459, w_eco74460, w_eco74461, w_eco74462, w_eco74463, w_eco74464, w_eco74465, w_eco74466, w_eco74467, w_eco74468, w_eco74469, w_eco74470, w_eco74471, w_eco74472, w_eco74473, w_eco74474, w_eco74475, w_eco74476, w_eco74477, w_eco74478, w_eco74479, w_eco74480, w_eco74481, w_eco74482, w_eco74483, w_eco74484, w_eco74485, w_eco74486, w_eco74487, w_eco74488, w_eco74489, w_eco74490, w_eco74491, w_eco74492, w_eco74493, w_eco74494, w_eco74495, w_eco74496, w_eco74497, w_eco74498, w_eco74499, w_eco74500, w_eco74501, w_eco74502, w_eco74503, w_eco74504, w_eco74505, w_eco74506, w_eco74507, w_eco74508, w_eco74509, w_eco74510, w_eco74511, w_eco74512, w_eco74513, w_eco74514, w_eco74515, w_eco74516, w_eco74517, w_eco74518, w_eco74519, w_eco74520, w_eco74521, w_eco74522, w_eco74523, w_eco74524, w_eco74525, w_eco74526, w_eco74527, w_eco74528, w_eco74529, w_eco74530, w_eco74531, w_eco74532, w_eco74533, w_eco74534, w_eco74535, w_eco74536, w_eco74537, w_eco74538, w_eco74539, w_eco74540, w_eco74541, w_eco74542, w_eco74543, w_eco74544, w_eco74545, w_eco74546, w_eco74547, w_eco74548, w_eco74549, w_eco74550, w_eco74551, w_eco74552, w_eco74553, w_eco74554, w_eco74555, w_eco74556, w_eco74557, w_eco74558, w_eco74559, w_eco74560, w_eco74561, w_eco74562, w_eco74563, w_eco74564, w_eco74565, w_eco74566, w_eco74567, w_eco74568, w_eco74569, w_eco74570, w_eco74571, w_eco74572, w_eco74573, w_eco74574, w_eco74575, w_eco74576, w_eco74577, w_eco74578, w_eco74579, w_eco74580, w_eco74581, w_eco74582, w_eco74583, w_eco74584, w_eco74585, w_eco74586, w_eco74587, w_eco74588, w_eco74589, w_eco74590, w_eco74591, w_eco74592, w_eco74593, w_eco74594, w_eco74595, w_eco74596, w_eco74597, w_eco74598, w_eco74599, w_eco74600, w_eco74601, w_eco74602, w_eco74603, w_eco74604, w_eco74605, w_eco74606, w_eco74607, w_eco74608, w_eco74609, w_eco74610, w_eco74611, w_eco74612, w_eco74613, w_eco74614, w_eco74615, w_eco74616, w_eco74617, w_eco74618, w_eco74619, w_eco74620, w_eco74621, w_eco74622, w_eco74623, w_eco74624, w_eco74625, w_eco74626, w_eco74627, w_eco74628, w_eco74629, w_eco74630, w_eco74631, w_eco74632, w_eco74633, w_eco74634, w_eco74635, w_eco74636, w_eco74637, w_eco74638, w_eco74639, w_eco74640, w_eco74641, w_eco74642, w_eco74643, w_eco74644, w_eco74645, w_eco74646, w_eco74647, w_eco74648, w_eco74649, w_eco74650, w_eco74651, w_eco74652, w_eco74653, w_eco74654, w_eco74655, w_eco74656, w_eco74657, w_eco74658, w_eco74659, w_eco74660, w_eco74661, w_eco74662, w_eco74663, w_eco74664, w_eco74665, w_eco74666, w_eco74667, w_eco74668, w_eco74669, w_eco74670, w_eco74671, w_eco74672, w_eco74673, w_eco74674, w_eco74675, w_eco74676, w_eco74677, w_eco74678, w_eco74679, w_eco74680, w_eco74681, w_eco74682, w_eco74683, w_eco74684, w_eco74685, w_eco74686, w_eco74687, w_eco74688, w_eco74689, w_eco74690, w_eco74691, w_eco74692, w_eco74693, w_eco74694, w_eco74695, w_eco74696, w_eco74697, w_eco74698, w_eco74699, w_eco74700, w_eco74701, w_eco74702, w_eco74703, w_eco74704, w_eco74705, w_eco74706, w_eco74707, w_eco74708, w_eco74709, w_eco74710, w_eco74711, w_eco74712, w_eco74713, w_eco74714, w_eco74715, w_eco74716, w_eco74717, w_eco74718, w_eco74719, w_eco74720, w_eco74721, w_eco74722, w_eco74723, w_eco74724, w_eco74725, w_eco74726, w_eco74727, w_eco74728, w_eco74729, w_eco74730, w_eco74731, w_eco74732, w_eco74733, w_eco74734, w_eco74735, w_eco74736, w_eco74737, w_eco74738, w_eco74739, w_eco74740, w_eco74741, w_eco74742, w_eco74743, w_eco74744, w_eco74745, w_eco74746, w_eco74747, w_eco74748, w_eco74749, w_eco74750, w_eco74751, w_eco74752, w_eco74753, w_eco74754, w_eco74755, w_eco74756, w_eco74757, w_eco74758, w_eco74759, w_eco74760, w_eco74761, w_eco74762, w_eco74763, w_eco74764, w_eco74765, w_eco74766, w_eco74767, w_eco74768, w_eco74769, w_eco74770, w_eco74771, w_eco74772, w_eco74773, w_eco74774, w_eco74775, w_eco74776, w_eco74777, w_eco74778, w_eco74779, w_eco74780, w_eco74781, w_eco74782, w_eco74783, w_eco74784, w_eco74785, w_eco74786, w_eco74787, w_eco74788, w_eco74789, w_eco74790, w_eco74791, w_eco74792, w_eco74793, w_eco74794, w_eco74795, w_eco74796, w_eco74797, w_eco74798, w_eco74799, w_eco74800, w_eco74801, w_eco74802, w_eco74803, w_eco74804, w_eco74805, w_eco74806, w_eco74807, w_eco74808, w_eco74809, w_eco74810, w_eco74811, w_eco74812, w_eco74813, w_eco74814, w_eco74815, w_eco74816, w_eco74817, w_eco74818, w_eco74819, w_eco74820, w_eco74821, w_eco74822, w_eco74823, w_eco74824, w_eco74825, w_eco74826, w_eco74827, w_eco74828, w_eco74829, w_eco74830, w_eco74831, w_eco74832, w_eco74833, w_eco74834, w_eco74835, w_eco74836, w_eco74837, w_eco74838, w_eco74839, w_eco74840, w_eco74841, w_eco74842, w_eco74843, w_eco74844, w_eco74845, w_eco74846, w_eco74847, w_eco74848, w_eco74849, w_eco74850, w_eco74851, w_eco74852, w_eco74853, w_eco74854, w_eco74855, w_eco74856, w_eco74857, w_eco74858, w_eco74859, w_eco74860, w_eco74861, w_eco74862, w_eco74863, w_eco74864, w_eco74865, w_eco74866, w_eco74867, w_eco74868, w_eco74869, w_eco74870, w_eco74871, w_eco74872, w_eco74873, w_eco74874, w_eco74875, w_eco74876, w_eco74877, w_eco74878, w_eco74879, w_eco74880, w_eco74881, w_eco74882, w_eco74883, w_eco74884, w_eco74885, w_eco74886, w_eco74887, w_eco74888, w_eco74889, w_eco74890, w_eco74891, w_eco74892, w_eco74893, w_eco74894, w_eco74895, w_eco74896, w_eco74897, w_eco74898, w_eco74899, w_eco74900, w_eco74901, w_eco74902, w_eco74903, w_eco74904, w_eco74905, w_eco74906, w_eco74907, w_eco74908, w_eco74909, w_eco74910, w_eco74911, w_eco74912, w_eco74913, w_eco74914, w_eco74915, w_eco74916, w_eco74917, w_eco74918, w_eco74919, w_eco74920, w_eco74921, w_eco74922, w_eco74923, w_eco74924, w_eco74925, w_eco74926, w_eco74927, w_eco74928, w_eco74929, w_eco74930, w_eco74931, w_eco74932, w_eco74933, w_eco74934, w_eco74935, w_eco74936, w_eco74937, w_eco74938, w_eco74939, w_eco74940, w_eco74941, w_eco74942, w_eco74943, w_eco74944, w_eco74945, w_eco74946, w_eco74947, w_eco74948, w_eco74949, w_eco74950, w_eco74951, w_eco74952, w_eco74953, w_eco74954, w_eco74955, w_eco74956, w_eco74957, w_eco74958, w_eco74959, w_eco74960, w_eco74961, w_eco74962, w_eco74963, w_eco74964, w_eco74965, w_eco74966, w_eco74967, w_eco74968, w_eco74969, w_eco74970, w_eco74971, w_eco74972, w_eco74973, w_eco74974, w_eco74975, w_eco74976, w_eco74977, w_eco74978, w_eco74979, w_eco74980, w_eco74981, w_eco74982, w_eco74983, w_eco74984, w_eco74985, w_eco74986, w_eco74987, w_eco74988, w_eco74989, w_eco74990, w_eco74991, w_eco74992, w_eco74993, w_eco74994, w_eco74995, w_eco74996, w_eco74997, w_eco74998, w_eco74999, w_eco75000, w_eco75001, w_eco75002, w_eco75003, w_eco75004, w_eco75005, w_eco75006, w_eco75007, w_eco75008, w_eco75009, w_eco75010, w_eco75011, w_eco75012, w_eco75013, w_eco75014, w_eco75015, w_eco75016, w_eco75017, w_eco75018, w_eco75019, w_eco75020, w_eco75021, w_eco75022, w_eco75023, w_eco75024, w_eco75025, w_eco75026, w_eco75027, w_eco75028, w_eco75029, w_eco75030, w_eco75031, w_eco75032, w_eco75033, w_eco75034, w_eco75035, w_eco75036, w_eco75037, w_eco75038, w_eco75039, w_eco75040, w_eco75041, w_eco75042, w_eco75043, w_eco75044, w_eco75045, w_eco75046, w_eco75047, w_eco75048, w_eco75049, w_eco75050, w_eco75051, w_eco75052, w_eco75053, w_eco75054, w_eco75055, w_eco75056, w_eco75057, w_eco75058, w_eco75059, w_eco75060, w_eco75061, w_eco75062, w_eco75063, w_eco75064, w_eco75065, w_eco75066, w_eco75067, w_eco75068, w_eco75069, w_eco75070, w_eco75071, w_eco75072, w_eco75073, w_eco75074, w_eco75075, w_eco75076, w_eco75077, w_eco75078, w_eco75079, w_eco75080, w_eco75081, w_eco75082, w_eco75083, w_eco75084, w_eco75085, w_eco75086, w_eco75087, w_eco75088, w_eco75089, w_eco75090, w_eco75091, w_eco75092, w_eco75093, w_eco75094, w_eco75095, w_eco75096, w_eco75097, w_eco75098, w_eco75099, w_eco75100, w_eco75101, w_eco75102, w_eco75103, w_eco75104, w_eco75105, w_eco75106, w_eco75107, w_eco75108, w_eco75109, w_eco75110, w_eco75111, w_eco75112, w_eco75113, w_eco75114, w_eco75115, w_eco75116, w_eco75117, w_eco75118, w_eco75119, w_eco75120, w_eco75121, w_eco75122, w_eco75123, w_eco75124, w_eco75125, w_eco75126, w_eco75127, w_eco75128, w_eco75129, w_eco75130, w_eco75131, w_eco75132, w_eco75133, w_eco75134, w_eco75135, w_eco75136, w_eco75137, w_eco75138, w_eco75139, w_eco75140, w_eco75141, w_eco75142, w_eco75143, w_eco75144, w_eco75145, w_eco75146, w_eco75147, w_eco75148, w_eco75149, w_eco75150, w_eco75151, w_eco75152, w_eco75153, w_eco75154, w_eco75155, w_eco75156, w_eco75157, w_eco75158, w_eco75159, w_eco75160, w_eco75161, w_eco75162, w_eco75163, w_eco75164, w_eco75165, w_eco75166, w_eco75167, w_eco75168, w_eco75169, w_eco75170, w_eco75171, w_eco75172, w_eco75173, w_eco75174, w_eco75175, w_eco75176, w_eco75177, w_eco75178, w_eco75179, w_eco75180, w_eco75181, w_eco75182, w_eco75183, w_eco75184, w_eco75185, w_eco75186, w_eco75187, w_eco75188, w_eco75189, w_eco75190, w_eco75191, w_eco75192, w_eco75193, w_eco75194, w_eco75195, w_eco75196, w_eco75197, w_eco75198, w_eco75199, w_eco75200, w_eco75201, w_eco75202, w_eco75203, w_eco75204, w_eco75205, w_eco75206, w_eco75207, w_eco75208, w_eco75209, w_eco75210, w_eco75211, w_eco75212, w_eco75213, w_eco75214, w_eco75215, w_eco75216, w_eco75217, w_eco75218, w_eco75219, w_eco75220, w_eco75221, w_eco75222, w_eco75223, w_eco75224, w_eco75225, w_eco75226, w_eco75227, w_eco75228, w_eco75229, w_eco75230, w_eco75231, w_eco75232, w_eco75233, w_eco75234, w_eco75235, w_eco75236, w_eco75237, w_eco75238, w_eco75239, w_eco75240, w_eco75241, w_eco75242, w_eco75243, w_eco75244, w_eco75245, w_eco75246, w_eco75247, w_eco75248, w_eco75249, w_eco75250, w_eco75251, w_eco75252, w_eco75253, w_eco75254, w_eco75255, w_eco75256, w_eco75257, w_eco75258, w_eco75259, w_eco75260, w_eco75261, w_eco75262, w_eco75263, w_eco75264, w_eco75265, w_eco75266, w_eco75267, w_eco75268, w_eco75269, w_eco75270, w_eco75271, w_eco75272, w_eco75273, w_eco75274, w_eco75275, w_eco75276, w_eco75277, w_eco75278, w_eco75279, w_eco75280, w_eco75281, w_eco75282, w_eco75283, w_eco75284, w_eco75285, w_eco75286, w_eco75287, w_eco75288, w_eco75289, w_eco75290, w_eco75291, w_eco75292, w_eco75293, w_eco75294, w_eco75295, w_eco75296, w_eco75297, w_eco75298, w_eco75299, w_eco75300, w_eco75301, w_eco75302, w_eco75303, w_eco75304, w_eco75305, w_eco75306, w_eco75307, w_eco75308, w_eco75309, w_eco75310, w_eco75311, w_eco75312, w_eco75313, w_eco75314, w_eco75315, w_eco75316, w_eco75317, w_eco75318, w_eco75319, w_eco75320, w_eco75321, w_eco75322, w_eco75323, w_eco75324, w_eco75325, w_eco75326, w_eco75327, w_eco75328, w_eco75329, w_eco75330, w_eco75331, w_eco75332, w_eco75333, w_eco75334, w_eco75335, w_eco75336, w_eco75337, w_eco75338, w_eco75339, w_eco75340, w_eco75341, w_eco75342, w_eco75343, w_eco75344, w_eco75345, w_eco75346, w_eco75347, w_eco75348, w_eco75349, w_eco75350, w_eco75351, w_eco75352, w_eco75353, w_eco75354, w_eco75355, w_eco75356, w_eco75357, w_eco75358, w_eco75359, w_eco75360, w_eco75361, w_eco75362, w_eco75363, w_eco75364, w_eco75365, w_eco75366, w_eco75367, w_eco75368, w_eco75369, w_eco75370, w_eco75371, w_eco75372, w_eco75373, w_eco75374, w_eco75375, w_eco75376, w_eco75377, w_eco75378, w_eco75379, w_eco75380, w_eco75381, w_eco75382, w_eco75383, w_eco75384, w_eco75385, w_eco75386, w_eco75387, w_eco75388, w_eco75389, w_eco75390, w_eco75391, w_eco75392, w_eco75393, w_eco75394, w_eco75395, w_eco75396, w_eco75397, w_eco75398, w_eco75399, w_eco75400, w_eco75401, w_eco75402, w_eco75403, w_eco75404, w_eco75405, w_eco75406, w_eco75407, w_eco75408, w_eco75409, w_eco75410, w_eco75411, w_eco75412, w_eco75413, w_eco75414, w_eco75415, w_eco75416, w_eco75417, w_eco75418, w_eco75419, w_eco75420, w_eco75421, w_eco75422, w_eco75423, w_eco75424, w_eco75425, w_eco75426, w_eco75427, w_eco75428, w_eco75429, w_eco75430, w_eco75431, w_eco75432, w_eco75433, w_eco75434, w_eco75435, w_eco75436, w_eco75437, w_eco75438, w_eco75439, w_eco75440, w_eco75441, w_eco75442, w_eco75443, w_eco75444, w_eco75445, w_eco75446, w_eco75447, w_eco75448, w_eco75449, w_eco75450, w_eco75451, w_eco75452, w_eco75453, w_eco75454, w_eco75455, w_eco75456, w_eco75457, w_eco75458, w_eco75459, w_eco75460, w_eco75461, w_eco75462, w_eco75463, w_eco75464, w_eco75465, w_eco75466, w_eco75467, w_eco75468, w_eco75469, w_eco75470, w_eco75471, w_eco75472, w_eco75473, w_eco75474, w_eco75475, w_eco75476, w_eco75477, w_eco75478, w_eco75479, w_eco75480, w_eco75481, w_eco75482, w_eco75483, w_eco75484, w_eco75485, w_eco75486, w_eco75487, w_eco75488, w_eco75489, w_eco75490, w_eco75491, w_eco75492, w_eco75493, w_eco75494, w_eco75495, w_eco75496, w_eco75497, w_eco75498, w_eco75499, w_eco75500, w_eco75501, w_eco75502, w_eco75503, w_eco75504, w_eco75505, w_eco75506, w_eco75507, w_eco75508, w_eco75509, w_eco75510, w_eco75511, w_eco75512, w_eco75513, w_eco75514, w_eco75515, w_eco75516, w_eco75517, w_eco75518, w_eco75519, w_eco75520, w_eco75521, w_eco75522, w_eco75523, w_eco75524, w_eco75525, w_eco75526, w_eco75527, w_eco75528, w_eco75529, w_eco75530, w_eco75531, w_eco75532, w_eco75533, w_eco75534, w_eco75535, w_eco75536, w_eco75537, w_eco75538, w_eco75539, w_eco75540, w_eco75541, w_eco75542, w_eco75543, w_eco75544, w_eco75545, w_eco75546, w_eco75547, w_eco75548, w_eco75549, w_eco75550, w_eco75551, w_eco75552, w_eco75553, w_eco75554, w_eco75555, w_eco75556, w_eco75557, w_eco75558, w_eco75559, w_eco75560, w_eco75561, w_eco75562, w_eco75563, w_eco75564, w_eco75565, w_eco75566, w_eco75567, w_eco75568, w_eco75569, w_eco75570, w_eco75571, w_eco75572, w_eco75573, w_eco75574, w_eco75575, w_eco75576, w_eco75577, w_eco75578, w_eco75579, w_eco75580, w_eco75581, w_eco75582, w_eco75583, w_eco75584, w_eco75585, w_eco75586, w_eco75587, w_eco75588, w_eco75589, w_eco75590, w_eco75591, w_eco75592, w_eco75593, w_eco75594, w_eco75595, w_eco75596, w_eco75597, w_eco75598, w_eco75599, w_eco75600, w_eco75601, w_eco75602, w_eco75603, w_eco75604, w_eco75605, w_eco75606, w_eco75607, w_eco75608, w_eco75609, w_eco75610, w_eco75611, w_eco75612, w_eco75613, w_eco75614, w_eco75615, w_eco75616, w_eco75617, w_eco75618, w_eco75619, w_eco75620, w_eco75621, w_eco75622, w_eco75623, w_eco75624, w_eco75625, w_eco75626, w_eco75627, w_eco75628, w_eco75629, w_eco75630, w_eco75631, w_eco75632, w_eco75633, w_eco75634, w_eco75635, w_eco75636, w_eco75637, w_eco75638, w_eco75639, w_eco75640, w_eco75641, w_eco75642, w_eco75643, w_eco75644, w_eco75645, w_eco75646, w_eco75647, w_eco75648, w_eco75649, w_eco75650, w_eco75651, w_eco75652, w_eco75653, w_eco75654, w_eco75655, w_eco75656, w_eco75657, w_eco75658, w_eco75659, w_eco75660, w_eco75661, w_eco75662, w_eco75663, w_eco75664, w_eco75665, w_eco75666, w_eco75667, w_eco75668, w_eco75669, w_eco75670, w_eco75671, w_eco75672, w_eco75673, w_eco75674, w_eco75675, w_eco75676, w_eco75677, w_eco75678, w_eco75679, w_eco75680, w_eco75681, w_eco75682, w_eco75683, w_eco75684, w_eco75685, w_eco75686, w_eco75687, w_eco75688, w_eco75689, w_eco75690, w_eco75691, w_eco75692, w_eco75693, w_eco75694, w_eco75695, w_eco75696, w_eco75697, w_eco75698, w_eco75699, w_eco75700, w_eco75701, w_eco75702, w_eco75703, w_eco75704, w_eco75705, w_eco75706, w_eco75707, w_eco75708, w_eco75709, w_eco75710, w_eco75711, w_eco75712, w_eco75713, w_eco75714, w_eco75715, w_eco75716, w_eco75717, w_eco75718, w_eco75719, w_eco75720, w_eco75721, w_eco75722, w_eco75723, w_eco75724, w_eco75725, w_eco75726, w_eco75727, w_eco75728, w_eco75729, w_eco75730, w_eco75731, w_eco75732, w_eco75733, w_eco75734, w_eco75735, w_eco75736, w_eco75737, w_eco75738, w_eco75739, w_eco75740, w_eco75741, w_eco75742, w_eco75743, w_eco75744, w_eco75745, w_eco75746, w_eco75747, w_eco75748, w_eco75749, w_eco75750, w_eco75751, w_eco75752, w_eco75753, w_eco75754, w_eco75755, w_eco75756, w_eco75757, w_eco75758, w_eco75759, w_eco75760, w_eco75761, w_eco75762, w_eco75763, w_eco75764, w_eco75765, w_eco75766, w_eco75767, w_eco75768, w_eco75769, w_eco75770, w_eco75771, w_eco75772, w_eco75773, w_eco75774, w_eco75775, w_eco75776, w_eco75777, w_eco75778, w_eco75779, w_eco75780, w_eco75781, w_eco75782, w_eco75783, w_eco75784, w_eco75785, w_eco75786, w_eco75787, w_eco75788, w_eco75789, w_eco75790, w_eco75791, w_eco75792, w_eco75793, w_eco75794, w_eco75795, w_eco75796, w_eco75797, w_eco75798, w_eco75799, w_eco75800, w_eco75801, w_eco75802, w_eco75803, w_eco75804, w_eco75805, w_eco75806, w_eco75807, w_eco75808, w_eco75809, w_eco75810, w_eco75811, w_eco75812, w_eco75813, w_eco75814, w_eco75815, w_eco75816, w_eco75817, w_eco75818, w_eco75819, w_eco75820, w_eco75821, w_eco75822, w_eco75823, w_eco75824, w_eco75825, w_eco75826, w_eco75827, w_eco75828, w_eco75829, w_eco75830, w_eco75831, w_eco75832, w_eco75833, w_eco75834, w_eco75835, w_eco75836, w_eco75837, w_eco75838, w_eco75839, w_eco75840, w_eco75841, w_eco75842, w_eco75843, w_eco75844, w_eco75845, w_eco75846, w_eco75847, w_eco75848, w_eco75849, w_eco75850, w_eco75851, w_eco75852, w_eco75853, w_eco75854, w_eco75855, w_eco75856, w_eco75857, w_eco75858, w_eco75859, w_eco75860, w_eco75861, w_eco75862, w_eco75863, w_eco75864, w_eco75865, w_eco75866, w_eco75867, w_eco75868, w_eco75869, w_eco75870, w_eco75871, w_eco75872, w_eco75873, w_eco75874, w_eco75875, w_eco75876, w_eco75877, w_eco75878, w_eco75879, w_eco75880, w_eco75881, w_eco75882, w_eco75883, w_eco75884, w_eco75885, w_eco75886, w_eco75887, w_eco75888, w_eco75889, w_eco75890, w_eco75891, w_eco75892, w_eco75893, w_eco75894, w_eco75895, w_eco75896, w_eco75897, w_eco75898, w_eco75899, w_eco75900, w_eco75901, w_eco75902, w_eco75903, w_eco75904, w_eco75905, w_eco75906, w_eco75907, w_eco75908, w_eco75909, w_eco75910, w_eco75911, w_eco75912, w_eco75913, w_eco75914, w_eco75915, w_eco75916, w_eco75917, w_eco75918, w_eco75919, w_eco75920, w_eco75921, w_eco75922, w_eco75923, w_eco75924, w_eco75925, w_eco75926, w_eco75927, w_eco75928, w_eco75929, w_eco75930, w_eco75931, w_eco75932, w_eco75933, w_eco75934, w_eco75935, w_eco75936, w_eco75937, w_eco75938, w_eco75939, w_eco75940, w_eco75941, w_eco75942, w_eco75943, w_eco75944, w_eco75945, w_eco75946, w_eco75947, w_eco75948, w_eco75949, w_eco75950, w_eco75951, w_eco75952, w_eco75953, w_eco75954, w_eco75955, w_eco75956, w_eco75957, w_eco75958, w_eco75959, w_eco75960, w_eco75961, w_eco75962, w_eco75963, w_eco75964, w_eco75965, w_eco75966, w_eco75967, w_eco75968, w_eco75969, w_eco75970, w_eco75971, w_eco75972, w_eco75973, w_eco75974, w_eco75975, w_eco75976, w_eco75977, w_eco75978, w_eco75979, w_eco75980, w_eco75981, w_eco75982, w_eco75983, w_eco75984, w_eco75985, w_eco75986, w_eco75987, w_eco75988, w_eco75989, w_eco75990, w_eco75991, w_eco75992, w_eco75993, w_eco75994, w_eco75995, w_eco75996, w_eco75997, w_eco75998, w_eco75999, w_eco76000, w_eco76001, w_eco76002, w_eco76003, w_eco76004, w_eco76005, w_eco76006, w_eco76007, w_eco76008, w_eco76009, w_eco76010, w_eco76011, w_eco76012, w_eco76013, w_eco76014, w_eco76015, w_eco76016, w_eco76017, w_eco76018, w_eco76019, w_eco76020, w_eco76021, w_eco76022, w_eco76023, w_eco76024, w_eco76025, w_eco76026, w_eco76027, w_eco76028, w_eco76029, w_eco76030, w_eco76031, w_eco76032, w_eco76033, w_eco76034, w_eco76035, w_eco76036, w_eco76037, w_eco76038, w_eco76039, w_eco76040, w_eco76041, w_eco76042, w_eco76043, w_eco76044, w_eco76045, w_eco76046, w_eco76047, w_eco76048, w_eco76049, w_eco76050, w_eco76051, w_eco76052, w_eco76053, w_eco76054, w_eco76055, w_eco76056, w_eco76057, w_eco76058, w_eco76059, w_eco76060, w_eco76061, w_eco76062, w_eco76063, w_eco76064, w_eco76065, w_eco76066, w_eco76067, w_eco76068, w_eco76069, w_eco76070, w_eco76071, w_eco76072, w_eco76073, w_eco76074, w_eco76075, w_eco76076, w_eco76077, w_eco76078, w_eco76079, w_eco76080, w_eco76081, w_eco76082, w_eco76083, w_eco76084, w_eco76085, w_eco76086, w_eco76087, w_eco76088, w_eco76089, w_eco76090, w_eco76091, w_eco76092, w_eco76093, w_eco76094, w_eco76095, w_eco76096, w_eco76097, w_eco76098, w_eco76099, w_eco76100, w_eco76101, w_eco76102, w_eco76103, w_eco76104, w_eco76105, w_eco76106, w_eco76107, w_eco76108, w_eco76109, w_eco76110, w_eco76111, w_eco76112, w_eco76113, w_eco76114, w_eco76115, w_eco76116, w_eco76117, w_eco76118, w_eco76119, w_eco76120, w_eco76121, w_eco76122, w_eco76123, w_eco76124, w_eco76125, w_eco76126, w_eco76127, w_eco76128, w_eco76129, w_eco76130, w_eco76131, w_eco76132, w_eco76133, w_eco76134, w_eco76135, w_eco76136, w_eco76137, w_eco76138, w_eco76139, w_eco76140, w_eco76141, w_eco76142, w_eco76143, w_eco76144, w_eco76145, w_eco76146, w_eco76147, w_eco76148, w_eco76149, w_eco76150, w_eco76151, w_eco76152, w_eco76153, w_eco76154, w_eco76155, w_eco76156, w_eco76157, w_eco76158, w_eco76159, w_eco76160, w_eco76161, w_eco76162, w_eco76163, w_eco76164, w_eco76165, w_eco76166, w_eco76167, w_eco76168, w_eco76169, w_eco76170, w_eco76171, w_eco76172, w_eco76173, w_eco76174, w_eco76175, w_eco76176, w_eco76177, w_eco76178, w_eco76179, w_eco76180, w_eco76181, w_eco76182, w_eco76183, w_eco76184, w_eco76185, w_eco76186, w_eco76187, w_eco76188, w_eco76189, w_eco76190, w_eco76191, w_eco76192, w_eco76193, w_eco76194, w_eco76195, w_eco76196, w_eco76197, w_eco76198, w_eco76199, w_eco76200, w_eco76201, w_eco76202, w_eco76203, w_eco76204, w_eco76205, w_eco76206, w_eco76207, w_eco76208, w_eco76209, w_eco76210, w_eco76211, w_eco76212, w_eco76213, w_eco76214, w_eco76215, w_eco76216, w_eco76217, w_eco76218, w_eco76219, w_eco76220, w_eco76221, w_eco76222, w_eco76223, w_eco76224, w_eco76225, w_eco76226, w_eco76227, w_eco76228, w_eco76229, w_eco76230, w_eco76231, w_eco76232, w_eco76233, w_eco76234, w_eco76235, w_eco76236, w_eco76237, w_eco76238, w_eco76239, w_eco76240, w_eco76241, w_eco76242, w_eco76243, w_eco76244, w_eco76245, w_eco76246, w_eco76247, w_eco76248, w_eco76249, w_eco76250, w_eco76251, w_eco76252, w_eco76253, w_eco76254, w_eco76255, w_eco76256, w_eco76257, w_eco76258, w_eco76259, w_eco76260, w_eco76261, w_eco76262, w_eco76263, w_eco76264, w_eco76265, w_eco76266, w_eco76267, w_eco76268, w_eco76269, w_eco76270, w_eco76271, w_eco76272, w_eco76273, w_eco76274, w_eco76275, w_eco76276, w_eco76277, w_eco76278, w_eco76279, w_eco76280, w_eco76281, w_eco76282, w_eco76283, w_eco76284, w_eco76285, w_eco76286, w_eco76287, w_eco76288, w_eco76289, w_eco76290, w_eco76291, w_eco76292, w_eco76293, w_eco76294, w_eco76295, w_eco76296, w_eco76297, w_eco76298, w_eco76299, w_eco76300, w_eco76301, w_eco76302, w_eco76303, w_eco76304, w_eco76305, w_eco76306, w_eco76307, w_eco76308, w_eco76309, w_eco76310, w_eco76311, w_eco76312, w_eco76313, w_eco76314, w_eco76315, w_eco76316, w_eco76317, w_eco76318, w_eco76319, w_eco76320, w_eco76321, w_eco76322, w_eco76323, w_eco76324, w_eco76325, w_eco76326, w_eco76327, w_eco76328, w_eco76329, w_eco76330, w_eco76331, w_eco76332, w_eco76333, w_eco76334, w_eco76335, w_eco76336, w_eco76337, w_eco76338, w_eco76339, w_eco76340, w_eco76341, w_eco76342, w_eco76343, w_eco76344, w_eco76345, w_eco76346, w_eco76347, w_eco76348, w_eco76349, w_eco76350, w_eco76351, w_eco76352, w_eco76353, w_eco76354, w_eco76355, w_eco76356, w_eco76357, w_eco76358, w_eco76359, w_eco76360, w_eco76361, w_eco76362, w_eco76363, w_eco76364, w_eco76365, w_eco76366, w_eco76367, w_eco76368, w_eco76369, w_eco76370, w_eco76371, w_eco76372, w_eco76373, w_eco76374, w_eco76375, w_eco76376, w_eco76377, w_eco76378, w_eco76379, w_eco76380, w_eco76381, w_eco76382, w_eco76383, w_eco76384, w_eco76385, w_eco76386, w_eco76387, w_eco76388, w_eco76389, w_eco76390, w_eco76391, w_eco76392, w_eco76393, w_eco76394, w_eco76395, w_eco76396, w_eco76397, w_eco76398, w_eco76399, w_eco76400, w_eco76401, w_eco76402, w_eco76403, w_eco76404, w_eco76405, w_eco76406, w_eco76407, w_eco76408, w_eco76409, w_eco76410, w_eco76411, w_eco76412, w_eco76413, w_eco76414, w_eco76415, w_eco76416, w_eco76417, w_eco76418, w_eco76419, w_eco76420, w_eco76421, w_eco76422, w_eco76423, w_eco76424, w_eco76425, w_eco76426, w_eco76427, w_eco76428, w_eco76429, w_eco76430, w_eco76431, w_eco76432, w_eco76433, w_eco76434, w_eco76435, w_eco76436, w_eco76437, w_eco76438, w_eco76439, w_eco76440, w_eco76441, w_eco76442, w_eco76443, w_eco76444, w_eco76445, w_eco76446, w_eco76447, w_eco76448, w_eco76449, w_eco76450, w_eco76451, w_eco76452, w_eco76453, w_eco76454, w_eco76455, w_eco76456, w_eco76457, w_eco76458, w_eco76459, w_eco76460, w_eco76461, w_eco76462, w_eco76463, w_eco76464, w_eco76465, w_eco76466, w_eco76467, w_eco76468, w_eco76469, w_eco76470, w_eco76471, w_eco76472, w_eco76473, w_eco76474, w_eco76475, w_eco76476, w_eco76477, w_eco76478, w_eco76479, w_eco76480, w_eco76481, w_eco76482, w_eco76483, w_eco76484, w_eco76485, w_eco76486, w_eco76487, w_eco76488, w_eco76489, w_eco76490, w_eco76491, w_eco76492, w_eco76493, w_eco76494, w_eco76495, w_eco76496, w_eco76497, w_eco76498, w_eco76499, w_eco76500, w_eco76501, w_eco76502, w_eco76503, w_eco76504, w_eco76505, w_eco76506, w_eco76507, w_eco76508, w_eco76509, w_eco76510, w_eco76511, w_eco76512, w_eco76513, w_eco76514, w_eco76515, w_eco76516, w_eco76517, w_eco76518, w_eco76519, w_eco76520, w_eco76521, w_eco76522, w_eco76523, w_eco76524, w_eco76525, w_eco76526, w_eco76527, w_eco76528, w_eco76529, w_eco76530, w_eco76531, w_eco76532, w_eco76533, w_eco76534, w_eco76535, w_eco76536, w_eco76537, w_eco76538, w_eco76539, w_eco76540, w_eco76541, w_eco76542, w_eco76543, w_eco76544, w_eco76545, w_eco76546, w_eco76547, w_eco76548, w_eco76549, w_eco76550, w_eco76551, w_eco76552, w_eco76553, w_eco76554, w_eco76555, w_eco76556, w_eco76557, w_eco76558, w_eco76559, w_eco76560, w_eco76561, w_eco76562, w_eco76563, w_eco76564, w_eco76565, w_eco76566, w_eco76567, w_eco76568, w_eco76569, w_eco76570, w_eco76571, w_eco76572, w_eco76573, w_eco76574, w_eco76575, w_eco76576, w_eco76577, w_eco76578, w_eco76579, w_eco76580, w_eco76581, w_eco76582, w_eco76583, w_eco76584, w_eco76585, w_eco76586, w_eco76587, w_eco76588, w_eco76589, w_eco76590, w_eco76591, w_eco76592, w_eco76593, w_eco76594, w_eco76595, w_eco76596, w_eco76597, w_eco76598, w_eco76599, w_eco76600, w_eco76601, w_eco76602, w_eco76603, w_eco76604, w_eco76605, w_eco76606, w_eco76607, w_eco76608, w_eco76609, w_eco76610, w_eco76611, w_eco76612, w_eco76613, w_eco76614, w_eco76615, w_eco76616, w_eco76617, w_eco76618, w_eco76619, w_eco76620, w_eco76621, w_eco76622, w_eco76623, w_eco76624, w_eco76625, w_eco76626, w_eco76627, w_eco76628, w_eco76629, w_eco76630, w_eco76631, w_eco76632, w_eco76633, w_eco76634, w_eco76635, w_eco76636, w_eco76637, w_eco76638, w_eco76639, w_eco76640, w_eco76641, w_eco76642, w_eco76643, w_eco76644, w_eco76645, w_eco76646, w_eco76647, w_eco76648, w_eco76649, w_eco76650, w_eco76651, w_eco76652, w_eco76653, w_eco76654, w_eco76655, w_eco76656, w_eco76657, w_eco76658, w_eco76659, w_eco76660, w_eco76661, w_eco76662, w_eco76663, w_eco76664, w_eco76665, w_eco76666, w_eco76667, w_eco76668, w_eco76669, w_eco76670, w_eco76671, w_eco76672, w_eco76673, w_eco76674, w_eco76675, w_eco76676, w_eco76677, w_eco76678, w_eco76679, w_eco76680, w_eco76681, w_eco76682, w_eco76683, w_eco76684, w_eco76685, w_eco76686, w_eco76687, w_eco76688, w_eco76689, w_eco76690, w_eco76691, w_eco76692, w_eco76693, w_eco76694, w_eco76695, w_eco76696, w_eco76697, w_eco76698, w_eco76699, w_eco76700, w_eco76701, w_eco76702, w_eco76703, w_eco76704, w_eco76705, w_eco76706, w_eco76707, w_eco76708, w_eco76709, w_eco76710, w_eco76711, w_eco76712, w_eco76713, w_eco76714, w_eco76715, w_eco76716, w_eco76717, w_eco76718, w_eco76719, w_eco76720, w_eco76721, w_eco76722, w_eco76723, w_eco76724, w_eco76725, w_eco76726, w_eco76727, w_eco76728, w_eco76729, w_eco76730, w_eco76731, w_eco76732, w_eco76733, w_eco76734, w_eco76735, w_eco76736, w_eco76737, w_eco76738, w_eco76739, w_eco76740, w_eco76741, w_eco76742, w_eco76743, w_eco76744, w_eco76745, w_eco76746, w_eco76747, w_eco76748, w_eco76749, w_eco76750, w_eco76751, w_eco76752, w_eco76753, w_eco76754, w_eco76755, w_eco76756, w_eco76757, w_eco76758, w_eco76759, w_eco76760, w_eco76761, w_eco76762, w_eco76763, w_eco76764, w_eco76765, w_eco76766, w_eco76767, w_eco76768, w_eco76769, w_eco76770, w_eco76771, w_eco76772, w_eco76773, w_eco76774, w_eco76775, w_eco76776, w_eco76777, w_eco76778, w_eco76779, w_eco76780, w_eco76781, w_eco76782, w_eco76783, w_eco76784, w_eco76785, w_eco76786, w_eco76787, w_eco76788, w_eco76789, w_eco76790, w_eco76791, w_eco76792, w_eco76793, w_eco76794, w_eco76795, w_eco76796, w_eco76797, w_eco76798, w_eco76799, w_eco76800, w_eco76801, w_eco76802, w_eco76803, w_eco76804, w_eco76805, w_eco76806, w_eco76807, w_eco76808, w_eco76809, w_eco76810, w_eco76811, w_eco76812, w_eco76813, w_eco76814, w_eco76815, w_eco76816, w_eco76817, w_eco76818, w_eco76819, w_eco76820, w_eco76821, w_eco76822, w_eco76823, w_eco76824, w_eco76825, w_eco76826, w_eco76827, w_eco76828, w_eco76829, w_eco76830, w_eco76831, w_eco76832, w_eco76833, w_eco76834, w_eco76835, w_eco76836, w_eco76837, w_eco76838, w_eco76839, w_eco76840, w_eco76841, w_eco76842, w_eco76843, w_eco76844, w_eco76845, w_eco76846, w_eco76847, w_eco76848, w_eco76849, w_eco76850, w_eco76851, w_eco76852, w_eco76853, w_eco76854, w_eco76855, w_eco76856, w_eco76857, w_eco76858, w_eco76859, w_eco76860, w_eco76861, w_eco76862, w_eco76863, w_eco76864, w_eco76865, w_eco76866, w_eco76867, w_eco76868, w_eco76869, w_eco76870, w_eco76871, w_eco76872, w_eco76873, w_eco76874, w_eco76875, w_eco76876, w_eco76877, w_eco76878, w_eco76879, w_eco76880, w_eco76881, w_eco76882, w_eco76883, w_eco76884, w_eco76885, w_eco76886, w_eco76887, w_eco76888, w_eco76889, w_eco76890, w_eco76891, w_eco76892, w_eco76893, w_eco76894, w_eco76895, w_eco76896, w_eco76897, w_eco76898, w_eco76899, w_eco76900, w_eco76901, w_eco76902, w_eco76903, w_eco76904, w_eco76905, w_eco76906, w_eco76907, w_eco76908, w_eco76909, w_eco76910, w_eco76911, w_eco76912, w_eco76913, w_eco76914, w_eco76915, w_eco76916, w_eco76917, w_eco76918, w_eco76919, w_eco76920, w_eco76921, w_eco76922, w_eco76923, w_eco76924, w_eco76925, w_eco76926, w_eco76927, w_eco76928, w_eco76929, w_eco76930, w_eco76931, w_eco76932, w_eco76933, w_eco76934, w_eco76935, w_eco76936, w_eco76937, w_eco76938, w_eco76939, w_eco76940, w_eco76941, w_eco76942, w_eco76943, w_eco76944, w_eco76945, w_eco76946, w_eco76947, w_eco76948, w_eco76949, w_eco76950, w_eco76951, w_eco76952, w_eco76953, w_eco76954, w_eco76955, w_eco76956, w_eco76957, w_eco76958, w_eco76959, w_eco76960, w_eco76961, w_eco76962, w_eco76963, w_eco76964, w_eco76965, w_eco76966, w_eco76967, w_eco76968, w_eco76969, w_eco76970, w_eco76971, w_eco76972, w_eco76973, w_eco76974, w_eco76975, w_eco76976, w_eco76977, w_eco76978, w_eco76979, w_eco76980, w_eco76981, w_eco76982, w_eco76983, w_eco76984, w_eco76985, w_eco76986, w_eco76987, w_eco76988, w_eco76989, w_eco76990, w_eco76991, w_eco76992, w_eco76993, w_eco76994, w_eco76995, w_eco76996, w_eco76997, w_eco76998, w_eco76999, w_eco77000, w_eco77001, w_eco77002, w_eco77003, w_eco77004, w_eco77005, w_eco77006, w_eco77007, w_eco77008, w_eco77009, w_eco77010, w_eco77011, w_eco77012, w_eco77013, w_eco77014, w_eco77015, w_eco77016, w_eco77017, w_eco77018, w_eco77019, w_eco77020, w_eco77021, w_eco77022, w_eco77023, w_eco77024, w_eco77025, w_eco77026, w_eco77027, w_eco77028, w_eco77029, w_eco77030, w_eco77031, w_eco77032, w_eco77033, w_eco77034, w_eco77035, w_eco77036, w_eco77037, w_eco77038, w_eco77039, w_eco77040, w_eco77041, w_eco77042, w_eco77043, w_eco77044, w_eco77045, w_eco77046, w_eco77047, w_eco77048, w_eco77049, w_eco77050, w_eco77051, w_eco77052, w_eco77053, w_eco77054, w_eco77055, w_eco77056, w_eco77057, w_eco77058, w_eco77059, w_eco77060, w_eco77061, w_eco77062, w_eco77063, w_eco77064, w_eco77065, w_eco77066, w_eco77067, w_eco77068, w_eco77069, w_eco77070, w_eco77071, w_eco77072, w_eco77073, w_eco77074, w_eco77075, w_eco77076, w_eco77077, w_eco77078, w_eco77079, w_eco77080, w_eco77081, w_eco77082, w_eco77083, w_eco77084, w_eco77085, w_eco77086, w_eco77087, w_eco77088, w_eco77089, w_eco77090, w_eco77091, w_eco77092, w_eco77093, w_eco77094, w_eco77095, w_eco77096, w_eco77097, w_eco77098, w_eco77099, w_eco77100, w_eco77101, w_eco77102, w_eco77103, w_eco77104, w_eco77105, w_eco77106, w_eco77107, w_eco77108, w_eco77109, w_eco77110, w_eco77111, w_eco77112, w_eco77113, w_eco77114, w_eco77115, w_eco77116, w_eco77117, w_eco77118, w_eco77119, w_eco77120, w_eco77121, w_eco77122, w_eco77123, w_eco77124, w_eco77125, w_eco77126, w_eco77127, w_eco77128, w_eco77129, w_eco77130, w_eco77131, w_eco77132, w_eco77133, w_eco77134, w_eco77135, w_eco77136, w_eco77137, w_eco77138, w_eco77139, w_eco77140, w_eco77141, w_eco77142, w_eco77143, w_eco77144, w_eco77145, w_eco77146, w_eco77147, w_eco77148, w_eco77149, w_eco77150, w_eco77151, w_eco77152, w_eco77153, w_eco77154, w_eco77155, w_eco77156, w_eco77157, w_eco77158, w_eco77159, w_eco77160, w_eco77161, w_eco77162, w_eco77163, w_eco77164, w_eco77165, w_eco77166, w_eco77167, w_eco77168, w_eco77169, w_eco77170, w_eco77171, w_eco77172, w_eco77173, w_eco77174, w_eco77175, w_eco77176, w_eco77177, w_eco77178, w_eco77179, w_eco77180, w_eco77181, w_eco77182, w_eco77183, w_eco77184, w_eco77185, w_eco77186, w_eco77187, w_eco77188, w_eco77189, w_eco77190, w_eco77191, w_eco77192, w_eco77193, w_eco77194, w_eco77195, w_eco77196, w_eco77197, w_eco77198, w_eco77199, w_eco77200, w_eco77201, w_eco77202, w_eco77203, w_eco77204, w_eco77205, w_eco77206, w_eco77207, w_eco77208, w_eco77209, w_eco77210, w_eco77211, w_eco77212, w_eco77213, w_eco77214, w_eco77215, w_eco77216, w_eco77217, w_eco77218, w_eco77219, w_eco77220, w_eco77221, w_eco77222, w_eco77223, w_eco77224, w_eco77225, w_eco77226, w_eco77227, w_eco77228, w_eco77229, w_eco77230, w_eco77231, w_eco77232, w_eco77233, w_eco77234, w_eco77235, w_eco77236, w_eco77237, w_eco77238, w_eco77239, w_eco77240, w_eco77241, w_eco77242, w_eco77243, w_eco77244, w_eco77245, w_eco77246, w_eco77247, w_eco77248, w_eco77249, w_eco77250, w_eco77251, w_eco77252, w_eco77253, w_eco77254, w_eco77255, w_eco77256, w_eco77257, w_eco77258, w_eco77259, w_eco77260, w_eco77261, w_eco77262, w_eco77263, w_eco77264, w_eco77265, w_eco77266, w_eco77267, w_eco77268, w_eco77269, w_eco77270, w_eco77271, w_eco77272, w_eco77273, w_eco77274, w_eco77275, w_eco77276, w_eco77277, w_eco77278, w_eco77279, w_eco77280, w_eco77281, w_eco77282, w_eco77283, w_eco77284, w_eco77285, w_eco77286, w_eco77287, w_eco77288, w_eco77289, w_eco77290, w_eco77291, w_eco77292, w_eco77293, w_eco77294, w_eco77295, w_eco77296, w_eco77297, w_eco77298, w_eco77299, w_eco77300, w_eco77301, w_eco77302, w_eco77303, w_eco77304, w_eco77305, w_eco77306, w_eco77307, w_eco77308, w_eco77309, w_eco77310, w_eco77311, w_eco77312, w_eco77313, w_eco77314, w_eco77315, w_eco77316, w_eco77317, w_eco77318, w_eco77319, w_eco77320, w_eco77321, w_eco77322, w_eco77323, w_eco77324, w_eco77325, w_eco77326, w_eco77327, w_eco77328, w_eco77329, w_eco77330, w_eco77331, w_eco77332, w_eco77333, w_eco77334, w_eco77335, w_eco77336, w_eco77337, w_eco77338, w_eco77339, w_eco77340, w_eco77341, w_eco77342, w_eco77343, w_eco77344, w_eco77345, w_eco77346, w_eco77347, w_eco77348, w_eco77349, w_eco77350, w_eco77351, w_eco77352, w_eco77353, w_eco77354, w_eco77355, w_eco77356, w_eco77357, w_eco77358, w_eco77359, w_eco77360, w_eco77361, w_eco77362, w_eco77363, w_eco77364, w_eco77365, w_eco77366, w_eco77367, w_eco77368, w_eco77369, w_eco77370, w_eco77371, w_eco77372, w_eco77373, w_eco77374, w_eco77375, w_eco77376, w_eco77377, w_eco77378, w_eco77379, w_eco77380, w_eco77381, w_eco77382, w_eco77383, w_eco77384, w_eco77385, w_eco77386, w_eco77387, w_eco77388, w_eco77389, w_eco77390, w_eco77391, w_eco77392, w_eco77393, w_eco77394, w_eco77395, w_eco77396, w_eco77397, w_eco77398, w_eco77399, w_eco77400, w_eco77401, w_eco77402, w_eco77403, w_eco77404, w_eco77405, w_eco77406, w_eco77407, w_eco77408, w_eco77409, w_eco77410, w_eco77411, w_eco77412, w_eco77413, w_eco77414, w_eco77415, w_eco77416, w_eco77417, w_eco77418, w_eco77419, w_eco77420, w_eco77421, w_eco77422, w_eco77423, w_eco77424, w_eco77425, w_eco77426, w_eco77427, w_eco77428, w_eco77429, w_eco77430, w_eco77431, w_eco77432, w_eco77433, w_eco77434, w_eco77435, w_eco77436, w_eco77437, w_eco77438, w_eco77439, w_eco77440, w_eco77441, w_eco77442, w_eco77443, w_eco77444, w_eco77445, w_eco77446, w_eco77447, w_eco77448, w_eco77449, w_eco77450, w_eco77451, w_eco77452, w_eco77453, w_eco77454, w_eco77455, w_eco77456, w_eco77457, w_eco77458, w_eco77459, w_eco77460, w_eco77461, w_eco77462, w_eco77463, w_eco77464, w_eco77465, w_eco77466, w_eco77467, w_eco77468, w_eco77469, w_eco77470, w_eco77471, w_eco77472, w_eco77473, w_eco77474, w_eco77475, w_eco77476, w_eco77477, w_eco77478, w_eco77479, w_eco77480, w_eco77481, w_eco77482, w_eco77483, w_eco77484, w_eco77485, w_eco77486, w_eco77487, w_eco77488, w_eco77489, w_eco77490, w_eco77491, w_eco77492, w_eco77493, w_eco77494, w_eco77495, w_eco77496, w_eco77497, w_eco77498, w_eco77499, w_eco77500, w_eco77501, w_eco77502, w_eco77503, w_eco77504, w_eco77505, w_eco77506, w_eco77507, w_eco77508, w_eco77509, w_eco77510, w_eco77511, w_eco77512, w_eco77513, w_eco77514, w_eco77515, w_eco77516, w_eco77517, w_eco77518, w_eco77519, w_eco77520, w_eco77521, w_eco77522, w_eco77523, w_eco77524, w_eco77525, w_eco77526, w_eco77527, w_eco77528, w_eco77529, w_eco77530, w_eco77531, w_eco77532, w_eco77533, w_eco77534, w_eco77535, w_eco77536, w_eco77537, w_eco77538, w_eco77539, w_eco77540, w_eco77541, w_eco77542, w_eco77543, w_eco77544, w_eco77545, w_eco77546, w_eco77547, w_eco77548, w_eco77549, w_eco77550, w_eco77551, w_eco77552, w_eco77553, w_eco77554, w_eco77555, w_eco77556, w_eco77557, w_eco77558, w_eco77559, w_eco77560, w_eco77561, w_eco77562, w_eco77563, w_eco77564, w_eco77565, w_eco77566, w_eco77567, w_eco77568, w_eco77569, w_eco77570, w_eco77571, w_eco77572, w_eco77573, w_eco77574, w_eco77575, w_eco77576, w_eco77577, w_eco77578, w_eco77579, w_eco77580, w_eco77581, w_eco77582, w_eco77583, w_eco77584, w_eco77585, w_eco77586, w_eco77587, w_eco77588, w_eco77589, w_eco77590, w_eco77591, w_eco77592, w_eco77593, w_eco77594, w_eco77595, w_eco77596, w_eco77597, w_eco77598, w_eco77599, w_eco77600, w_eco77601, w_eco77602, w_eco77603, w_eco77604, w_eco77605, w_eco77606, w_eco77607, w_eco77608, w_eco77609, w_eco77610, w_eco77611, w_eco77612, w_eco77613, w_eco77614, w_eco77615, w_eco77616, w_eco77617, w_eco77618, w_eco77619, w_eco77620, w_eco77621, w_eco77622, w_eco77623, w_eco77624, w_eco77625, w_eco77626, w_eco77627, w_eco77628, w_eco77629, w_eco77630, w_eco77631, w_eco77632, w_eco77633, w_eco77634, w_eco77635, w_eco77636, w_eco77637, w_eco77638, w_eco77639, w_eco77640, w_eco77641, w_eco77642, w_eco77643, w_eco77644, w_eco77645, w_eco77646, w_eco77647, w_eco77648, w_eco77649, w_eco77650, w_eco77651, w_eco77652, w_eco77653, w_eco77654, w_eco77655, w_eco77656, w_eco77657, w_eco77658, w_eco77659, w_eco77660, w_eco77661, w_eco77662, w_eco77663, w_eco77664, w_eco77665, w_eco77666, w_eco77667, w_eco77668, w_eco77669, w_eco77670, w_eco77671, w_eco77672, w_eco77673, w_eco77674, w_eco77675, w_eco77676, w_eco77677, w_eco77678, w_eco77679, w_eco77680, w_eco77681, w_eco77682, w_eco77683, w_eco77684, w_eco77685, w_eco77686, w_eco77687, w_eco77688, w_eco77689, w_eco77690, w_eco77691, w_eco77692, w_eco77693, w_eco77694, w_eco77695, w_eco77696, w_eco77697, w_eco77698, w_eco77699, w_eco77700, w_eco77701, w_eco77702, w_eco77703, w_eco77704, w_eco77705, w_eco77706, w_eco77707, w_eco77708, w_eco77709, w_eco77710, w_eco77711, w_eco77712, w_eco77713, w_eco77714, w_eco77715, w_eco77716, w_eco77717, w_eco77718, w_eco77719, w_eco77720, w_eco77721, w_eco77722, w_eco77723, w_eco77724, w_eco77725, w_eco77726, w_eco77727, w_eco77728, w_eco77729, w_eco77730, w_eco77731, w_eco77732, w_eco77733, w_eco77734, w_eco77735, w_eco77736, w_eco77737, w_eco77738, w_eco77739, w_eco77740, w_eco77741, w_eco77742, w_eco77743, w_eco77744, w_eco77745, w_eco77746, w_eco77747, w_eco77748, w_eco77749, w_eco77750, w_eco77751, w_eco77752, w_eco77753, w_eco77754, w_eco77755, w_eco77756, w_eco77757, w_eco77758, w_eco77759, w_eco77760, w_eco77761, w_eco77762, w_eco77763, w_eco77764, w_eco77765, w_eco77766, w_eco77767, w_eco77768, w_eco77769, w_eco77770, w_eco77771, w_eco77772, w_eco77773, w_eco77774, w_eco77775, w_eco77776, w_eco77777, w_eco77778, w_eco77779, w_eco77780, w_eco77781, w_eco77782, w_eco77783, w_eco77784, w_eco77785, w_eco77786, w_eco77787, w_eco77788, w_eco77789, w_eco77790, w_eco77791, w_eco77792, w_eco77793, w_eco77794, w_eco77795, w_eco77796, w_eco77797, w_eco77798, w_eco77799, w_eco77800, w_eco77801, w_eco77802, w_eco77803, w_eco77804, w_eco77805, w_eco77806, w_eco77807, w_eco77808, w_eco77809, w_eco77810, w_eco77811, w_eco77812, w_eco77813, w_eco77814, w_eco77815, w_eco77816, w_eco77817, w_eco77818, w_eco77819, w_eco77820, w_eco77821, w_eco77822, w_eco77823, w_eco77824, w_eco77825, w_eco77826, w_eco77827, w_eco77828, w_eco77829, w_eco77830, w_eco77831, w_eco77832, w_eco77833, w_eco77834, w_eco77835, w_eco77836, w_eco77837, w_eco77838, w_eco77839, w_eco77840, w_eco77841, w_eco77842, w_eco77843, w_eco77844, w_eco77845, w_eco77846, w_eco77847, w_eco77848, w_eco77849, w_eco77850, w_eco77851, w_eco77852, w_eco77853, w_eco77854, w_eco77855, w_eco77856, w_eco77857, w_eco77858, w_eco77859, w_eco77860, w_eco77861, w_eco77862, w_eco77863, w_eco77864, w_eco77865, w_eco77866, w_eco77867, w_eco77868, w_eco77869, w_eco77870, w_eco77871, w_eco77872, w_eco77873, w_eco77874, w_eco77875, w_eco77876, w_eco77877, w_eco77878, w_eco77879, w_eco77880, w_eco77881, w_eco77882, w_eco77883, w_eco77884, w_eco77885, w_eco77886, w_eco77887, w_eco77888, w_eco77889, w_eco77890, w_eco77891, w_eco77892, w_eco77893, w_eco77894, w_eco77895, w_eco77896, w_eco77897, w_eco77898, w_eco77899, w_eco77900, w_eco77901, w_eco77902, w_eco77903, w_eco77904, w_eco77905, w_eco77906, w_eco77907, w_eco77908, w_eco77909, w_eco77910, w_eco77911, w_eco77912, w_eco77913, w_eco77914, w_eco77915, w_eco77916, w_eco77917, w_eco77918, w_eco77919, w_eco77920, w_eco77921, w_eco77922, w_eco77923, w_eco77924, w_eco77925, w_eco77926, w_eco77927, w_eco77928, w_eco77929, w_eco77930, w_eco77931, w_eco77932, w_eco77933, w_eco77934, w_eco77935, w_eco77936, w_eco77937, w_eco77938, w_eco77939, w_eco77940, w_eco77941, w_eco77942, w_eco77943, w_eco77944, w_eco77945, w_eco77946, w_eco77947, w_eco77948, w_eco77949, w_eco77950, w_eco77951, w_eco77952, w_eco77953, w_eco77954, w_eco77955, w_eco77956, w_eco77957, w_eco77958, w_eco77959, w_eco77960, w_eco77961, w_eco77962, w_eco77963, w_eco77964, w_eco77965, w_eco77966, w_eco77967, w_eco77968, w_eco77969, w_eco77970, w_eco77971, w_eco77972, w_eco77973, w_eco77974, w_eco77975, w_eco77976, w_eco77977, w_eco77978, w_eco77979, w_eco77980, w_eco77981, w_eco77982, w_eco77983, w_eco77984, w_eco77985, w_eco77986, w_eco77987, w_eco77988, w_eco77989, w_eco77990, w_eco77991, w_eco77992, w_eco77993, w_eco77994, w_eco77995, w_eco77996, w_eco77997, w_eco77998, w_eco77999, w_eco78000, w_eco78001, w_eco78002, w_eco78003, w_eco78004, w_eco78005, w_eco78006, w_eco78007, w_eco78008, w_eco78009, w_eco78010, w_eco78011, w_eco78012, w_eco78013, w_eco78014, w_eco78015, w_eco78016, w_eco78017, w_eco78018, w_eco78019, w_eco78020, w_eco78021, w_eco78022, w_eco78023, w_eco78024, w_eco78025, w_eco78026, w_eco78027, w_eco78028, w_eco78029, w_eco78030, w_eco78031, w_eco78032, w_eco78033, w_eco78034, w_eco78035, w_eco78036, w_eco78037, w_eco78038, w_eco78039, w_eco78040, w_eco78041, w_eco78042, w_eco78043, w_eco78044, w_eco78045, w_eco78046, w_eco78047, w_eco78048, w_eco78049, w_eco78050, w_eco78051, w_eco78052, w_eco78053, w_eco78054, w_eco78055, w_eco78056, w_eco78057, w_eco78058, w_eco78059, w_eco78060, w_eco78061, w_eco78062, w_eco78063, w_eco78064, w_eco78065, w_eco78066, w_eco78067, w_eco78068, w_eco78069, w_eco78070, w_eco78071, w_eco78072, w_eco78073, w_eco78074, w_eco78075, w_eco78076, w_eco78077, w_eco78078, w_eco78079, w_eco78080, w_eco78081, w_eco78082, w_eco78083, w_eco78084, w_eco78085, w_eco78086, w_eco78087, w_eco78088, w_eco78089, w_eco78090, w_eco78091, w_eco78092, w_eco78093, w_eco78094, w_eco78095, w_eco78096, w_eco78097, w_eco78098, w_eco78099, w_eco78100, w_eco78101, w_eco78102, w_eco78103, w_eco78104, w_eco78105, w_eco78106, w_eco78107, w_eco78108, w_eco78109, w_eco78110, w_eco78111, w_eco78112, w_eco78113, w_eco78114, w_eco78115, w_eco78116, w_eco78117, w_eco78118, w_eco78119, w_eco78120, w_eco78121, w_eco78122, w_eco78123, w_eco78124, w_eco78125, w_eco78126, w_eco78127, w_eco78128, w_eco78129, w_eco78130, w_eco78131, w_eco78132, w_eco78133, w_eco78134, w_eco78135, w_eco78136, w_eco78137, w_eco78138, w_eco78139, w_eco78140, w_eco78141, w_eco78142, w_eco78143, w_eco78144, w_eco78145, w_eco78146, w_eco78147, w_eco78148, w_eco78149, w_eco78150, w_eco78151, w_eco78152, w_eco78153, w_eco78154, w_eco78155, w_eco78156, w_eco78157, w_eco78158, w_eco78159, w_eco78160, w_eco78161, w_eco78162, w_eco78163, w_eco78164, w_eco78165, w_eco78166, w_eco78167, w_eco78168, w_eco78169, w_eco78170, w_eco78171, w_eco78172, w_eco78173, w_eco78174, w_eco78175, w_eco78176, w_eco78177, w_eco78178, w_eco78179, w_eco78180, w_eco78181, w_eco78182, w_eco78183, w_eco78184, w_eco78185, w_eco78186, w_eco78187, w_eco78188, w_eco78189, w_eco78190, w_eco78191, w_eco78192, w_eco78193, w_eco78194, w_eco78195, w_eco78196, w_eco78197, w_eco78198, w_eco78199, w_eco78200, w_eco78201, w_eco78202, w_eco78203, w_eco78204, w_eco78205, w_eco78206, w_eco78207, w_eco78208, w_eco78209, w_eco78210, w_eco78211, w_eco78212, w_eco78213, w_eco78214, w_eco78215, w_eco78216, w_eco78217, w_eco78218, w_eco78219, w_eco78220, w_eco78221, w_eco78222, w_eco78223, w_eco78224, w_eco78225, w_eco78226, w_eco78227, w_eco78228, w_eco78229, w_eco78230, w_eco78231, w_eco78232, w_eco78233, w_eco78234, w_eco78235, w_eco78236, w_eco78237, w_eco78238, w_eco78239, w_eco78240, w_eco78241, w_eco78242, w_eco78243, w_eco78244, w_eco78245, w_eco78246, w_eco78247, w_eco78248, w_eco78249, w_eco78250, w_eco78251, w_eco78252, w_eco78253, w_eco78254, w_eco78255, w_eco78256, w_eco78257, w_eco78258, w_eco78259, w_eco78260, w_eco78261, w_eco78262, w_eco78263, w_eco78264, w_eco78265, w_eco78266, w_eco78267, w_eco78268, w_eco78269, w_eco78270, w_eco78271, w_eco78272, w_eco78273, w_eco78274, w_eco78275, w_eco78276, w_eco78277, w_eco78278, w_eco78279, w_eco78280, w_eco78281, w_eco78282, w_eco78283, w_eco78284, w_eco78285, w_eco78286, w_eco78287, w_eco78288, w_eco78289, w_eco78290, w_eco78291, w_eco78292, w_eco78293, w_eco78294, w_eco78295, w_eco78296, w_eco78297, w_eco78298, w_eco78299, w_eco78300, w_eco78301, w_eco78302, w_eco78303, w_eco78304, w_eco78305, w_eco78306, w_eco78307, w_eco78308, w_eco78309, w_eco78310, w_eco78311, w_eco78312, w_eco78313, w_eco78314, w_eco78315, w_eco78316, w_eco78317, w_eco78318, w_eco78319, w_eco78320, w_eco78321, w_eco78322, w_eco78323, w_eco78324, w_eco78325, w_eco78326, w_eco78327, w_eco78328, w_eco78329, w_eco78330, w_eco78331, w_eco78332, w_eco78333, w_eco78334, w_eco78335, w_eco78336, w_eco78337, w_eco78338, w_eco78339, w_eco78340, w_eco78341, w_eco78342, w_eco78343, w_eco78344, w_eco78345, w_eco78346, w_eco78347, w_eco78348, w_eco78349, w_eco78350, w_eco78351, w_eco78352, w_eco78353, w_eco78354, w_eco78355, w_eco78356, w_eco78357, w_eco78358, w_eco78359, w_eco78360, w_eco78361, w_eco78362, w_eco78363, w_eco78364, w_eco78365, w_eco78366, w_eco78367, w_eco78368, w_eco78369, w_eco78370, w_eco78371, w_eco78372, w_eco78373, w_eco78374, w_eco78375, w_eco78376, w_eco78377, w_eco78378, w_eco78379, w_eco78380, w_eco78381, w_eco78382, w_eco78383, w_eco78384, w_eco78385, w_eco78386, w_eco78387, w_eco78388, w_eco78389, w_eco78390, w_eco78391, w_eco78392, w_eco78393, w_eco78394, w_eco78395, w_eco78396, w_eco78397, w_eco78398, w_eco78399, w_eco78400, w_eco78401, w_eco78402, w_eco78403, w_eco78404, w_eco78405, w_eco78406, w_eco78407, w_eco78408, w_eco78409, w_eco78410, w_eco78411, w_eco78412, w_eco78413, w_eco78414, w_eco78415, w_eco78416, w_eco78417, w_eco78418, w_eco78419, w_eco78420, w_eco78421, w_eco78422, w_eco78423, w_eco78424, w_eco78425, w_eco78426, w_eco78427, w_eco78428, w_eco78429, w_eco78430, w_eco78431, w_eco78432, w_eco78433, w_eco78434, w_eco78435, w_eco78436, w_eco78437, w_eco78438, w_eco78439, w_eco78440, w_eco78441, w_eco78442, w_eco78443, w_eco78444, w_eco78445, w_eco78446, w_eco78447, w_eco78448, w_eco78449, w_eco78450, w_eco78451, w_eco78452, w_eco78453, w_eco78454, w_eco78455, w_eco78456, w_eco78457, w_eco78458, w_eco78459, w_eco78460, w_eco78461, w_eco78462, w_eco78463, w_eco78464, w_eco78465, w_eco78466, w_eco78467, w_eco78468, w_eco78469, w_eco78470, w_eco78471, w_eco78472, w_eco78473, w_eco78474, w_eco78475, w_eco78476, w_eco78477, w_eco78478, w_eco78479, w_eco78480, w_eco78481, w_eco78482, w_eco78483, w_eco78484, w_eco78485, w_eco78486, w_eco78487, w_eco78488, w_eco78489, w_eco78490, w_eco78491, w_eco78492, w_eco78493, w_eco78494, w_eco78495, w_eco78496, w_eco78497, w_eco78498, w_eco78499, w_eco78500, w_eco78501, w_eco78502, w_eco78503, w_eco78504, w_eco78505, w_eco78506, w_eco78507, w_eco78508, w_eco78509, w_eco78510, w_eco78511, w_eco78512, w_eco78513, w_eco78514, w_eco78515, w_eco78516, w_eco78517, w_eco78518, w_eco78519, w_eco78520, w_eco78521, w_eco78522, w_eco78523, w_eco78524, w_eco78525, w_eco78526, w_eco78527, w_eco78528, w_eco78529, w_eco78530, w_eco78531, w_eco78532, w_eco78533, w_eco78534, w_eco78535, w_eco78536, w_eco78537, w_eco78538, w_eco78539, w_eco78540, w_eco78541, w_eco78542, w_eco78543, w_eco78544, w_eco78545, w_eco78546, w_eco78547, w_eco78548, w_eco78549, w_eco78550, w_eco78551, w_eco78552, w_eco78553, w_eco78554, w_eco78555, w_eco78556, w_eco78557, w_eco78558, w_eco78559, w_eco78560, w_eco78561, w_eco78562, w_eco78563, w_eco78564, w_eco78565, w_eco78566, w_eco78567, w_eco78568, w_eco78569, w_eco78570, w_eco78571, w_eco78572, w_eco78573, w_eco78574, w_eco78575, w_eco78576, w_eco78577, w_eco78578, w_eco78579, w_eco78580, w_eco78581, w_eco78582, w_eco78583, w_eco78584, w_eco78585, w_eco78586, w_eco78587, w_eco78588, w_eco78589, w_eco78590, w_eco78591, w_eco78592, w_eco78593, w_eco78594, w_eco78595, w_eco78596, w_eco78597, w_eco78598, w_eco78599, w_eco78600, w_eco78601, w_eco78602, w_eco78603, w_eco78604, w_eco78605, w_eco78606, w_eco78607, w_eco78608, w_eco78609, w_eco78610, w_eco78611, w_eco78612, w_eco78613, w_eco78614, w_eco78615, w_eco78616, w_eco78617, w_eco78618, w_eco78619, w_eco78620, w_eco78621, w_eco78622, w_eco78623, w_eco78624, w_eco78625, w_eco78626, w_eco78627, w_eco78628, w_eco78629, w_eco78630, w_eco78631, w_eco78632, w_eco78633, w_eco78634, w_eco78635, w_eco78636, w_eco78637, w_eco78638, w_eco78639, w_eco78640, w_eco78641, w_eco78642, w_eco78643, w_eco78644, w_eco78645, w_eco78646, w_eco78647, w_eco78648, w_eco78649, w_eco78650, w_eco78651, w_eco78652, w_eco78653, w_eco78654, w_eco78655, w_eco78656, w_eco78657, w_eco78658, w_eco78659, w_eco78660, w_eco78661, w_eco78662, w_eco78663, w_eco78664, w_eco78665, w_eco78666, w_eco78667, w_eco78668, w_eco78669, w_eco78670, w_eco78671, w_eco78672, w_eco78673, w_eco78674, w_eco78675, w_eco78676, w_eco78677, w_eco78678, w_eco78679, w_eco78680, w_eco78681, w_eco78682, w_eco78683, w_eco78684, w_eco78685, w_eco78686, w_eco78687, w_eco78688, w_eco78689, w_eco78690, w_eco78691, w_eco78692, w_eco78693, w_eco78694, w_eco78695, w_eco78696, w_eco78697, w_eco78698, w_eco78699, w_eco78700, w_eco78701, w_eco78702, w_eco78703, w_eco78704, w_eco78705, w_eco78706, w_eco78707, w_eco78708, w_eco78709, w_eco78710, w_eco78711, w_eco78712, w_eco78713, w_eco78714, w_eco78715, w_eco78716, w_eco78717, w_eco78718, w_eco78719, w_eco78720, w_eco78721, w_eco78722, w_eco78723, w_eco78724, w_eco78725, w_eco78726, w_eco78727, w_eco78728, w_eco78729, w_eco78730, w_eco78731, w_eco78732, w_eco78733, w_eco78734, w_eco78735, w_eco78736, w_eco78737, w_eco78738, w_eco78739, w_eco78740, w_eco78741, w_eco78742, w_eco78743, w_eco78744, w_eco78745, w_eco78746, w_eco78747, w_eco78748, w_eco78749, w_eco78750, w_eco78751, w_eco78752, w_eco78753, w_eco78754, w_eco78755, w_eco78756, w_eco78757, w_eco78758, w_eco78759, w_eco78760, w_eco78761, w_eco78762, w_eco78763, w_eco78764, w_eco78765, w_eco78766, w_eco78767, w_eco78768, w_eco78769, w_eco78770, w_eco78771, w_eco78772, w_eco78773, w_eco78774, w_eco78775, w_eco78776, w_eco78777, w_eco78778, w_eco78779, w_eco78780, w_eco78781, w_eco78782, w_eco78783, w_eco78784, w_eco78785, w_eco78786, w_eco78787, w_eco78788, w_eco78789, w_eco78790, w_eco78791, w_eco78792, w_eco78793, w_eco78794, w_eco78795, w_eco78796, w_eco78797, w_eco78798, w_eco78799, w_eco78800, w_eco78801, w_eco78802, w_eco78803, w_eco78804, w_eco78805, w_eco78806, w_eco78807, w_eco78808, w_eco78809, w_eco78810, w_eco78811, w_eco78812, w_eco78813, w_eco78814, w_eco78815, w_eco78816, w_eco78817, w_eco78818, w_eco78819, w_eco78820, w_eco78821, w_eco78822, w_eco78823, w_eco78824, w_eco78825, w_eco78826, w_eco78827, w_eco78828, w_eco78829, w_eco78830, w_eco78831, w_eco78832, w_eco78833, w_eco78834, w_eco78835, w_eco78836, w_eco78837, w_eco78838, w_eco78839, w_eco78840, w_eco78841, w_eco78842, w_eco78843, w_eco78844, w_eco78845, w_eco78846, w_eco78847, w_eco78848, w_eco78849, w_eco78850, w_eco78851, w_eco78852, w_eco78853, w_eco78854, w_eco78855, w_eco78856, w_eco78857, w_eco78858, w_eco78859, w_eco78860, w_eco78861, w_eco78862, w_eco78863, w_eco78864, w_eco78865, w_eco78866, w_eco78867, w_eco78868, w_eco78869, w_eco78870, w_eco78871, w_eco78872, w_eco78873, w_eco78874, w_eco78875, w_eco78876, w_eco78877, w_eco78878, w_eco78879, w_eco78880, w_eco78881, w_eco78882, w_eco78883, w_eco78884, w_eco78885, w_eco78886, w_eco78887, w_eco78888, w_eco78889, w_eco78890, w_eco78891, w_eco78892, w_eco78893, w_eco78894, w_eco78895, w_eco78896, w_eco78897, w_eco78898, w_eco78899, w_eco78900, w_eco78901, w_eco78902, w_eco78903, w_eco78904, w_eco78905, w_eco78906, w_eco78907, w_eco78908, w_eco78909, w_eco78910, w_eco78911, w_eco78912, w_eco78913, w_eco78914, w_eco78915, w_eco78916, w_eco78917, w_eco78918, w_eco78919, w_eco78920, w_eco78921, w_eco78922, w_eco78923, w_eco78924, w_eco78925, w_eco78926, w_eco78927, w_eco78928, w_eco78929, w_eco78930, w_eco78931, w_eco78932, w_eco78933, w_eco78934, w_eco78935, w_eco78936, w_eco78937, w_eco78938, w_eco78939, w_eco78940, w_eco78941, w_eco78942, w_eco78943, w_eco78944, w_eco78945, w_eco78946, w_eco78947, w_eco78948, w_eco78949, w_eco78950, w_eco78951, w_eco78952, w_eco78953, w_eco78954, w_eco78955, w_eco78956, w_eco78957, w_eco78958, w_eco78959, w_eco78960, w_eco78961, w_eco78962, w_eco78963, w_eco78964, w_eco78965, w_eco78966, w_eco78967, w_eco78968, w_eco78969, w_eco78970, w_eco78971, w_eco78972, w_eco78973, w_eco78974, w_eco78975, w_eco78976, w_eco78977, w_eco78978, w_eco78979, w_eco78980, w_eco78981, w_eco78982, w_eco78983, w_eco78984, w_eco78985, w_eco78986, w_eco78987, w_eco78988, w_eco78989, w_eco78990, w_eco78991, w_eco78992, w_eco78993, w_eco78994, w_eco78995, w_eco78996, w_eco78997, w_eco78998, w_eco78999, w_eco79000, w_eco79001, w_eco79002, w_eco79003, w_eco79004, w_eco79005, w_eco79006, w_eco79007, w_eco79008, w_eco79009, w_eco79010, w_eco79011, w_eco79012, w_eco79013, w_eco79014, w_eco79015, w_eco79016, w_eco79017, w_eco79018, w_eco79019, w_eco79020, w_eco79021, w_eco79022, w_eco79023, w_eco79024, w_eco79025, w_eco79026, w_eco79027, w_eco79028, w_eco79029, w_eco79030, w_eco79031, w_eco79032, w_eco79033, w_eco79034, w_eco79035, w_eco79036, w_eco79037, w_eco79038, w_eco79039, w_eco79040, w_eco79041, w_eco79042, w_eco79043, w_eco79044, w_eco79045, w_eco79046, w_eco79047, w_eco79048, w_eco79049, w_eco79050, w_eco79051, w_eco79052, w_eco79053, w_eco79054, w_eco79055, w_eco79056, w_eco79057, w_eco79058, w_eco79059, w_eco79060, w_eco79061, w_eco79062, w_eco79063, w_eco79064, w_eco79065, w_eco79066, w_eco79067, w_eco79068, w_eco79069, w_eco79070, w_eco79071, w_eco79072, w_eco79073, w_eco79074, w_eco79075, w_eco79076, w_eco79077, w_eco79078, w_eco79079, w_eco79080, w_eco79081, w_eco79082, w_eco79083, w_eco79084, w_eco79085, w_eco79086, w_eco79087, w_eco79088, w_eco79089, w_eco79090, w_eco79091, w_eco79092, w_eco79093, w_eco79094, w_eco79095, w_eco79096, w_eco79097, w_eco79098, w_eco79099, w_eco79100, w_eco79101, w_eco79102, w_eco79103, w_eco79104, w_eco79105, w_eco79106, w_eco79107, w_eco79108, w_eco79109, w_eco79110, w_eco79111, w_eco79112, w_eco79113, w_eco79114, w_eco79115, w_eco79116, w_eco79117, w_eco79118, w_eco79119, w_eco79120, w_eco79121, w_eco79122, w_eco79123, w_eco79124, w_eco79125, w_eco79126, w_eco79127, w_eco79128, w_eco79129, w_eco79130, w_eco79131, w_eco79132, w_eco79133, w_eco79134, w_eco79135, w_eco79136, w_eco79137, w_eco79138, w_eco79139, w_eco79140, w_eco79141, w_eco79142, w_eco79143, w_eco79144, w_eco79145, w_eco79146, w_eco79147, w_eco79148, w_eco79149, w_eco79150, w_eco79151, w_eco79152, w_eco79153, w_eco79154, w_eco79155, w_eco79156, w_eco79157, w_eco79158, w_eco79159, w_eco79160, w_eco79161, w_eco79162, w_eco79163, w_eco79164, w_eco79165, w_eco79166, w_eco79167, w_eco79168, w_eco79169, w_eco79170, w_eco79171, w_eco79172, w_eco79173, w_eco79174, w_eco79175, w_eco79176, w_eco79177, w_eco79178, w_eco79179, w_eco79180, w_eco79181, w_eco79182, w_eco79183, w_eco79184, w_eco79185, w_eco79186, w_eco79187, w_eco79188, w_eco79189, w_eco79190, w_eco79191, w_eco79192, w_eco79193, w_eco79194, w_eco79195, w_eco79196, w_eco79197, w_eco79198, w_eco79199, w_eco79200, w_eco79201, w_eco79202, w_eco79203, w_eco79204, w_eco79205, w_eco79206, w_eco79207, w_eco79208, w_eco79209, w_eco79210, w_eco79211, w_eco79212, w_eco79213, w_eco79214, w_eco79215, w_eco79216, w_eco79217, w_eco79218, w_eco79219, w_eco79220, w_eco79221, w_eco79222, w_eco79223, w_eco79224, w_eco79225, w_eco79226, w_eco79227, w_eco79228, w_eco79229, w_eco79230, w_eco79231, w_eco79232, w_eco79233, w_eco79234, w_eco79235, w_eco79236, w_eco79237, w_eco79238, w_eco79239, w_eco79240, w_eco79241, w_eco79242, w_eco79243, w_eco79244, w_eco79245, w_eco79246, w_eco79247, w_eco79248, w_eco79249, w_eco79250, w_eco79251, w_eco79252, w_eco79253, w_eco79254, w_eco79255, w_eco79256, w_eco79257, w_eco79258, w_eco79259, w_eco79260, w_eco79261, w_eco79262, w_eco79263, w_eco79264, w_eco79265, w_eco79266, w_eco79267, w_eco79268, w_eco79269, w_eco79270, w_eco79271, w_eco79272, w_eco79273, w_eco79274, w_eco79275, w_eco79276, w_eco79277, w_eco79278, w_eco79279, w_eco79280, w_eco79281, w_eco79282, w_eco79283, w_eco79284, w_eco79285, w_eco79286, w_eco79287, w_eco79288, w_eco79289, w_eco79290, w_eco79291, w_eco79292, w_eco79293, w_eco79294, w_eco79295, w_eco79296, w_eco79297, w_eco79298, w_eco79299, w_eco79300, w_eco79301, w_eco79302, w_eco79303, w_eco79304, w_eco79305, w_eco79306, w_eco79307, w_eco79308, w_eco79309, w_eco79310, w_eco79311, w_eco79312, w_eco79313, w_eco79314, w_eco79315, w_eco79316, w_eco79317, w_eco79318, w_eco79319, w_eco79320, w_eco79321, w_eco79322, w_eco79323, w_eco79324, w_eco79325, w_eco79326, w_eco79327, w_eco79328, w_eco79329, w_eco79330, w_eco79331, w_eco79332, w_eco79333, w_eco79334, w_eco79335, w_eco79336, w_eco79337, w_eco79338, w_eco79339, w_eco79340, w_eco79341, w_eco79342, w_eco79343, w_eco79344, w_eco79345, w_eco79346, w_eco79347, w_eco79348, w_eco79349, w_eco79350, w_eco79351, w_eco79352, w_eco79353, w_eco79354, w_eco79355, w_eco79356, w_eco79357, w_eco79358, w_eco79359, w_eco79360, w_eco79361, w_eco79362, w_eco79363, w_eco79364, w_eco79365, w_eco79366, w_eco79367, w_eco79368, w_eco79369, w_eco79370, w_eco79371, w_eco79372, w_eco79373, w_eco79374, w_eco79375, w_eco79376, w_eco79377, w_eco79378, w_eco79379, w_eco79380, w_eco79381, w_eco79382, w_eco79383, w_eco79384, w_eco79385, w_eco79386, w_eco79387, w_eco79388, w_eco79389, w_eco79390, w_eco79391, w_eco79392, w_eco79393, w_eco79394, w_eco79395, w_eco79396, w_eco79397, w_eco79398, w_eco79399, w_eco79400, w_eco79401, w_eco79402, w_eco79403, w_eco79404, w_eco79405, w_eco79406, w_eco79407, w_eco79408, w_eco79409, w_eco79410, w_eco79411, w_eco79412, w_eco79413, w_eco79414, w_eco79415, w_eco79416, w_eco79417, w_eco79418, w_eco79419, w_eco79420, w_eco79421, w_eco79422, w_eco79423, w_eco79424, w_eco79425, w_eco79426, w_eco79427, w_eco79428, w_eco79429, w_eco79430, w_eco79431, w_eco79432, w_eco79433, w_eco79434, w_eco79435, w_eco79436, w_eco79437, w_eco79438, w_eco79439, w_eco79440, w_eco79441, w_eco79442, w_eco79443, w_eco79444, w_eco79445, w_eco79446, w_eco79447, w_eco79448, w_eco79449, w_eco79450, w_eco79451, w_eco79452, w_eco79453, w_eco79454, w_eco79455, w_eco79456, w_eco79457, w_eco79458, w_eco79459, w_eco79460, w_eco79461, w_eco79462, w_eco79463, w_eco79464, w_eco79465, w_eco79466, w_eco79467, w_eco79468, w_eco79469, w_eco79470, w_eco79471, w_eco79472, w_eco79473, w_eco79474, w_eco79475, w_eco79476, w_eco79477, w_eco79478, w_eco79479, w_eco79480, w_eco79481, w_eco79482, w_eco79483, w_eco79484, w_eco79485, w_eco79486, w_eco79487, w_eco79488, w_eco79489, w_eco79490, w_eco79491, w_eco79492, w_eco79493, w_eco79494, w_eco79495, w_eco79496, w_eco79497, w_eco79498, w_eco79499, w_eco79500, w_eco79501, w_eco79502, w_eco79503, w_eco79504, w_eco79505, w_eco79506, w_eco79507, w_eco79508, w_eco79509, w_eco79510, w_eco79511, w_eco79512, w_eco79513, w_eco79514, w_eco79515, w_eco79516, w_eco79517, w_eco79518, w_eco79519, w_eco79520, w_eco79521, w_eco79522, w_eco79523, w_eco79524, w_eco79525, w_eco79526, w_eco79527, w_eco79528, w_eco79529, w_eco79530, w_eco79531, w_eco79532, w_eco79533, w_eco79534, w_eco79535, w_eco79536, w_eco79537, w_eco79538, w_eco79539, w_eco79540, w_eco79541, w_eco79542, w_eco79543, w_eco79544, w_eco79545, w_eco79546, w_eco79547, w_eco79548, w_eco79549, w_eco79550, w_eco79551, w_eco79552, w_eco79553, w_eco79554, w_eco79555, w_eco79556, w_eco79557, w_eco79558, w_eco79559, w_eco79560, w_eco79561, w_eco79562, w_eco79563, w_eco79564, w_eco79565, w_eco79566, w_eco79567, w_eco79568, w_eco79569, w_eco79570, w_eco79571, w_eco79572, w_eco79573, w_eco79574, w_eco79575, w_eco79576, w_eco79577, w_eco79578, w_eco79579, w_eco79580, w_eco79581, w_eco79582, w_eco79583, w_eco79584, w_eco79585, w_eco79586, w_eco79587, w_eco79588, w_eco79589, w_eco79590, w_eco79591, w_eco79592, w_eco79593, w_eco79594, w_eco79595, w_eco79596, w_eco79597, w_eco79598, w_eco79599, w_eco79600, w_eco79601, w_eco79602, w_eco79603, w_eco79604, w_eco79605, w_eco79606, w_eco79607, w_eco79608, w_eco79609, w_eco79610, w_eco79611, w_eco79612, w_eco79613, w_eco79614, w_eco79615, w_eco79616, w_eco79617, w_eco79618, w_eco79619, w_eco79620, w_eco79621, w_eco79622, w_eco79623, w_eco79624, w_eco79625, w_eco79626, w_eco79627, w_eco79628, w_eco79629, w_eco79630, w_eco79631, w_eco79632, w_eco79633, w_eco79634, w_eco79635, w_eco79636, w_eco79637, w_eco79638, w_eco79639, w_eco79640, w_eco79641, w_eco79642, w_eco79643, w_eco79644, w_eco79645, w_eco79646, w_eco79647, w_eco79648, w_eco79649, w_eco79650, w_eco79651, w_eco79652, w_eco79653, w_eco79654, w_eco79655, w_eco79656, w_eco79657, w_eco79658, w_eco79659, w_eco79660, w_eco79661, w_eco79662, w_eco79663, w_eco79664, w_eco79665, w_eco79666, w_eco79667, w_eco79668, w_eco79669, w_eco79670, w_eco79671, w_eco79672, w_eco79673, w_eco79674, w_eco79675, w_eco79676, w_eco79677, w_eco79678, w_eco79679, w_eco79680, w_eco79681, w_eco79682, w_eco79683, w_eco79684, w_eco79685, w_eco79686, w_eco79687, w_eco79688, w_eco79689, w_eco79690, w_eco79691, w_eco79692, w_eco79693, w_eco79694, w_eco79695, w_eco79696, w_eco79697, w_eco79698, w_eco79699, w_eco79700, w_eco79701, w_eco79702, w_eco79703, w_eco79704, w_eco79705, w_eco79706, w_eco79707, w_eco79708, w_eco79709, w_eco79710, w_eco79711, w_eco79712, w_eco79713, w_eco79714, w_eco79715, w_eco79716, w_eco79717, w_eco79718, w_eco79719, w_eco79720, w_eco79721, w_eco79722, w_eco79723, w_eco79724, w_eco79725, w_eco79726, w_eco79727, w_eco79728, w_eco79729, w_eco79730, w_eco79731, w_eco79732, w_eco79733, w_eco79734, w_eco79735, w_eco79736, w_eco79737, w_eco79738, w_eco79739, w_eco79740, w_eco79741, w_eco79742, w_eco79743, w_eco79744, w_eco79745, w_eco79746, w_eco79747, w_eco79748, w_eco79749, w_eco79750, w_eco79751, w_eco79752, w_eco79753, w_eco79754, w_eco79755, w_eco79756, w_eco79757, w_eco79758, w_eco79759, w_eco79760, w_eco79761, w_eco79762, w_eco79763, w_eco79764, w_eco79765, w_eco79766, w_eco79767, w_eco79768, w_eco79769, w_eco79770, w_eco79771, w_eco79772, w_eco79773, w_eco79774, w_eco79775, w_eco79776, w_eco79777, w_eco79778, w_eco79779, w_eco79780, w_eco79781, w_eco79782, w_eco79783, w_eco79784, w_eco79785, w_eco79786, w_eco79787, w_eco79788, w_eco79789, w_eco79790, w_eco79791, w_eco79792, w_eco79793, w_eco79794, w_eco79795, w_eco79796, w_eco79797, w_eco79798, w_eco79799, w_eco79800, w_eco79801, w_eco79802, w_eco79803, w_eco79804, w_eco79805, w_eco79806, w_eco79807, w_eco79808, w_eco79809, w_eco79810, w_eco79811, w_eco79812, w_eco79813, w_eco79814, w_eco79815, w_eco79816, w_eco79817, w_eco79818, w_eco79819, w_eco79820, w_eco79821, w_eco79822, w_eco79823, w_eco79824, w_eco79825, w_eco79826, w_eco79827, w_eco79828, w_eco79829, w_eco79830, w_eco79831, w_eco79832, w_eco79833, w_eco79834, w_eco79835, w_eco79836, w_eco79837, w_eco79838, w_eco79839, w_eco79840, w_eco79841, w_eco79842, w_eco79843, w_eco79844, w_eco79845, w_eco79846, w_eco79847, w_eco79848, w_eco79849, w_eco79850, w_eco79851, w_eco79852, w_eco79853, w_eco79854, w_eco79855, w_eco79856, w_eco79857, w_eco79858, w_eco79859, w_eco79860, w_eco79861, w_eco79862, w_eco79863, w_eco79864, w_eco79865, w_eco79866, w_eco79867, w_eco79868, w_eco79869, w_eco79870, w_eco79871, w_eco79872, w_eco79873, w_eco79874, w_eco79875, w_eco79876, w_eco79877, w_eco79878, w_eco79879, w_eco79880, w_eco79881, w_eco79882, w_eco79883, w_eco79884, w_eco79885, w_eco79886, w_eco79887, w_eco79888, w_eco79889, w_eco79890, w_eco79891, w_eco79892, w_eco79893, w_eco79894, w_eco79895, w_eco79896, w_eco79897, w_eco79898, w_eco79899, w_eco79900, w_eco79901, w_eco79902, w_eco79903, w_eco79904, w_eco79905, w_eco79906, w_eco79907, w_eco79908, w_eco79909, w_eco79910, w_eco79911, w_eco79912, w_eco79913, w_eco79914, w_eco79915, w_eco79916, w_eco79917, w_eco79918, w_eco79919, w_eco79920, w_eco79921, w_eco79922, w_eco79923, w_eco79924, w_eco79925, w_eco79926, w_eco79927, w_eco79928, w_eco79929, w_eco79930, w_eco79931, w_eco79932, w_eco79933, w_eco79934, w_eco79935, w_eco79936, w_eco79937, w_eco79938, w_eco79939, w_eco79940, w_eco79941, w_eco79942, w_eco79943, w_eco79944, w_eco79945, w_eco79946, w_eco79947, w_eco79948, w_eco79949, w_eco79950, w_eco79951, w_eco79952, w_eco79953, w_eco79954, w_eco79955, w_eco79956, w_eco79957, w_eco79958, w_eco79959, w_eco79960, w_eco79961, w_eco79962, w_eco79963, w_eco79964, w_eco79965, w_eco79966, w_eco79967, w_eco79968, w_eco79969, w_eco79970, w_eco79971, w_eco79972, w_eco79973, w_eco79974, w_eco79975, w_eco79976, w_eco79977, w_eco79978, w_eco79979, w_eco79980, w_eco79981, w_eco79982, w_eco79983, w_eco79984, w_eco79985, w_eco79986, w_eco79987, w_eco79988, w_eco79989, w_eco79990, w_eco79991, w_eco79992, w_eco79993, w_eco79994, w_eco79995, w_eco79996, w_eco79997, w_eco79998, w_eco79999, w_eco80000, w_eco80001, w_eco80002, w_eco80003, w_eco80004, w_eco80005, w_eco80006, w_eco80007, w_eco80008, w_eco80009, w_eco80010, w_eco80011, w_eco80012, w_eco80013, w_eco80014, w_eco80015, w_eco80016, w_eco80017, w_eco80018, w_eco80019, w_eco80020, w_eco80021, w_eco80022, w_eco80023, w_eco80024, w_eco80025, w_eco80026, w_eco80027, w_eco80028, w_eco80029, w_eco80030, w_eco80031, w_eco80032, w_eco80033, w_eco80034, w_eco80035, w_eco80036, w_eco80037, w_eco80038, w_eco80039, w_eco80040, w_eco80041, w_eco80042, w_eco80043, w_eco80044, w_eco80045, w_eco80046, w_eco80047, w_eco80048, w_eco80049, w_eco80050, w_eco80051, w_eco80052, w_eco80053, w_eco80054, w_eco80055, w_eco80056, w_eco80057, w_eco80058, w_eco80059, w_eco80060, w_eco80061, w_eco80062, w_eco80063, w_eco80064, w_eco80065, w_eco80066, w_eco80067, w_eco80068, w_eco80069, w_eco80070, w_eco80071, w_eco80072, w_eco80073, w_eco80074, w_eco80075, w_eco80076, w_eco80077, w_eco80078, w_eco80079, w_eco80080, w_eco80081, w_eco80082, w_eco80083, w_eco80084, w_eco80085, w_eco80086, w_eco80087, w_eco80088, w_eco80089, w_eco80090, w_eco80091, w_eco80092, w_eco80093, w_eco80094, w_eco80095, w_eco80096, w_eco80097, w_eco80098, w_eco80099, w_eco80100, w_eco80101, w_eco80102, w_eco80103, w_eco80104, w_eco80105, w_eco80106, w_eco80107, w_eco80108, w_eco80109, w_eco80110, w_eco80111, w_eco80112, w_eco80113, w_eco80114, w_eco80115, w_eco80116, w_eco80117, w_eco80118, w_eco80119, w_eco80120, w_eco80121, w_eco80122, w_eco80123, w_eco80124, w_eco80125, w_eco80126, w_eco80127, w_eco80128, w_eco80129, w_eco80130, w_eco80131, w_eco80132, w_eco80133, w_eco80134, w_eco80135, w_eco80136, w_eco80137, w_eco80138, w_eco80139, w_eco80140, w_eco80141, w_eco80142, w_eco80143, w_eco80144, w_eco80145, w_eco80146, w_eco80147, w_eco80148, w_eco80149, w_eco80150, w_eco80151, w_eco80152, w_eco80153, w_eco80154, w_eco80155, w_eco80156, w_eco80157, w_eco80158, w_eco80159, w_eco80160, w_eco80161, w_eco80162, w_eco80163, w_eco80164, w_eco80165, w_eco80166, w_eco80167, w_eco80168, w_eco80169, w_eco80170, w_eco80171, w_eco80172, w_eco80173, w_eco80174, w_eco80175, w_eco80176, w_eco80177, w_eco80178, w_eco80179, w_eco80180, w_eco80181, w_eco80182, w_eco80183, w_eco80184, w_eco80185, w_eco80186, w_eco80187, w_eco80188, w_eco80189, w_eco80190, w_eco80191, w_eco80192, w_eco80193, w_eco80194, w_eco80195, w_eco80196, w_eco80197, w_eco80198, w_eco80199, w_eco80200, w_eco80201, w_eco80202, w_eco80203, w_eco80204, w_eco80205, w_eco80206, w_eco80207, w_eco80208, w_eco80209, w_eco80210, w_eco80211, w_eco80212, w_eco80213, w_eco80214, w_eco80215, w_eco80216, w_eco80217, w_eco80218, w_eco80219, w_eco80220, w_eco80221, w_eco80222, w_eco80223, w_eco80224, w_eco80225, w_eco80226, w_eco80227, w_eco80228, w_eco80229, w_eco80230, w_eco80231, w_eco80232, w_eco80233, w_eco80234, w_eco80235, w_eco80236, w_eco80237, w_eco80238, w_eco80239, w_eco80240, w_eco80241, w_eco80242, w_eco80243, w_eco80244, w_eco80245, w_eco80246, w_eco80247, w_eco80248, w_eco80249, w_eco80250, w_eco80251, w_eco80252, w_eco80253, w_eco80254, w_eco80255, w_eco80256, w_eco80257, w_eco80258, w_eco80259, w_eco80260, w_eco80261, w_eco80262, w_eco80263, w_eco80264, w_eco80265, w_eco80266, w_eco80267, w_eco80268, w_eco80269, w_eco80270, w_eco80271, w_eco80272, w_eco80273, w_eco80274, w_eco80275, w_eco80276, w_eco80277, w_eco80278, w_eco80279, w_eco80280, w_eco80281, w_eco80282, w_eco80283, w_eco80284, w_eco80285, w_eco80286, w_eco80287, w_eco80288, w_eco80289, w_eco80290, w_eco80291, w_eco80292, w_eco80293, w_eco80294, w_eco80295, w_eco80296, w_eco80297, w_eco80298, w_eco80299, w_eco80300, w_eco80301, w_eco80302, w_eco80303, w_eco80304, w_eco80305, w_eco80306, w_eco80307, w_eco80308, w_eco80309, w_eco80310, w_eco80311, w_eco80312, w_eco80313, w_eco80314, w_eco80315, w_eco80316, w_eco80317, w_eco80318, w_eco80319, w_eco80320, w_eco80321, w_eco80322, w_eco80323, w_eco80324, w_eco80325, w_eco80326, w_eco80327, w_eco80328, w_eco80329, w_eco80330, w_eco80331, w_eco80332, w_eco80333, w_eco80334, w_eco80335, w_eco80336, w_eco80337, w_eco80338, w_eco80339, w_eco80340, w_eco80341, w_eco80342, w_eco80343, w_eco80344, w_eco80345, w_eco80346, w_eco80347, w_eco80348, w_eco80349, w_eco80350, w_eco80351, w_eco80352, w_eco80353, w_eco80354, w_eco80355, w_eco80356, w_eco80357, w_eco80358, w_eco80359, w_eco80360, w_eco80361, w_eco80362, w_eco80363, w_eco80364, w_eco80365, w_eco80366, w_eco80367, w_eco80368, w_eco80369, w_eco80370, w_eco80371, w_eco80372, w_eco80373, w_eco80374, w_eco80375, w_eco80376, w_eco80377, w_eco80378, w_eco80379, w_eco80380, w_eco80381, w_eco80382, w_eco80383, w_eco80384, w_eco80385, w_eco80386, w_eco80387, w_eco80388, w_eco80389, w_eco80390, w_eco80391, w_eco80392, w_eco80393, w_eco80394, w_eco80395, w_eco80396, w_eco80397, w_eco80398, w_eco80399, w_eco80400, w_eco80401, w_eco80402, w_eco80403, w_eco80404, w_eco80405, w_eco80406, w_eco80407, w_eco80408, w_eco80409, w_eco80410, w_eco80411, w_eco80412, w_eco80413, w_eco80414, w_eco80415, w_eco80416, w_eco80417, w_eco80418, w_eco80419, w_eco80420, w_eco80421, w_eco80422, w_eco80423, w_eco80424, w_eco80425, w_eco80426, w_eco80427, w_eco80428, w_eco80429, w_eco80430, w_eco80431, w_eco80432, w_eco80433, w_eco80434, w_eco80435, w_eco80436, w_eco80437, w_eco80438, w_eco80439, w_eco80440, w_eco80441, w_eco80442, w_eco80443, w_eco80444, w_eco80445, w_eco80446, w_eco80447, w_eco80448, w_eco80449, w_eco80450, w_eco80451, w_eco80452, w_eco80453, w_eco80454, w_eco80455, w_eco80456, w_eco80457, w_eco80458, w_eco80459, w_eco80460, w_eco80461, w_eco80462, w_eco80463, w_eco80464, w_eco80465, w_eco80466, w_eco80467, w_eco80468, w_eco80469, w_eco80470, w_eco80471, w_eco80472, w_eco80473, w_eco80474, w_eco80475, w_eco80476, w_eco80477, w_eco80478, w_eco80479, w_eco80480, w_eco80481, w_eco80482, w_eco80483, w_eco80484, w_eco80485, w_eco80486, w_eco80487, w_eco80488, w_eco80489, w_eco80490, w_eco80491, w_eco80492, w_eco80493, w_eco80494, w_eco80495, w_eco80496, w_eco80497, w_eco80498, w_eco80499, w_eco80500, w_eco80501, w_eco80502, w_eco80503, w_eco80504, w_eco80505, w_eco80506, w_eco80507, w_eco80508, w_eco80509, w_eco80510, w_eco80511, w_eco80512, w_eco80513, w_eco80514, w_eco80515, w_eco80516, w_eco80517, w_eco80518, w_eco80519, w_eco80520, w_eco80521, w_eco80522, w_eco80523, w_eco80524, w_eco80525, w_eco80526, w_eco80527, w_eco80528, w_eco80529, w_eco80530, w_eco80531, w_eco80532, w_eco80533, w_eco80534, w_eco80535, w_eco80536, w_eco80537, w_eco80538, w_eco80539, w_eco80540, w_eco80541, w_eco80542, w_eco80543, w_eco80544, w_eco80545, w_eco80546, w_eco80547, w_eco80548, w_eco80549, w_eco80550, w_eco80551, w_eco80552, w_eco80553, w_eco80554, w_eco80555, w_eco80556, w_eco80557, w_eco80558, w_eco80559, w_eco80560, w_eco80561, w_eco80562, w_eco80563, w_eco80564, w_eco80565, w_eco80566, w_eco80567, w_eco80568, w_eco80569, w_eco80570, w_eco80571, w_eco80572, w_eco80573, w_eco80574, w_eco80575, w_eco80576, w_eco80577, w_eco80578, w_eco80579, w_eco80580, w_eco80581, w_eco80582, w_eco80583, w_eco80584, w_eco80585, w_eco80586, w_eco80587, w_eco80588, w_eco80589, w_eco80590, w_eco80591, w_eco80592, w_eco80593, w_eco80594, w_eco80595, w_eco80596, w_eco80597, w_eco80598, w_eco80599, w_eco80600, w_eco80601, w_eco80602, w_eco80603, w_eco80604, w_eco80605, w_eco80606, w_eco80607, w_eco80608, w_eco80609, w_eco80610, w_eco80611, w_eco80612, w_eco80613, w_eco80614, w_eco80615, w_eco80616, w_eco80617, w_eco80618, w_eco80619, w_eco80620, w_eco80621, w_eco80622, w_eco80623, w_eco80624, w_eco80625, w_eco80626, w_eco80627, w_eco80628, w_eco80629, w_eco80630, w_eco80631, w_eco80632, w_eco80633, w_eco80634, w_eco80635, w_eco80636, w_eco80637, w_eco80638, w_eco80639, w_eco80640, w_eco80641, w_eco80642, w_eco80643, w_eco80644, w_eco80645, w_eco80646, w_eco80647, w_eco80648, w_eco80649, w_eco80650, w_eco80651, w_eco80652, w_eco80653, w_eco80654, w_eco80655, w_eco80656, w_eco80657, w_eco80658, w_eco80659, w_eco80660, w_eco80661, w_eco80662, w_eco80663, w_eco80664, w_eco80665, w_eco80666, w_eco80667, w_eco80668, w_eco80669, w_eco80670, w_eco80671, w_eco80672, w_eco80673, w_eco80674, w_eco80675, w_eco80676, w_eco80677, w_eco80678, w_eco80679, w_eco80680, w_eco80681, w_eco80682, w_eco80683, w_eco80684, w_eco80685, w_eco80686, w_eco80687, w_eco80688, w_eco80689, w_eco80690, w_eco80691, w_eco80692, w_eco80693, w_eco80694, w_eco80695, w_eco80696, w_eco80697, w_eco80698, w_eco80699, w_eco80700, w_eco80701, w_eco80702, w_eco80703, w_eco80704, w_eco80705, w_eco80706, w_eco80707, w_eco80708, w_eco80709, w_eco80710, w_eco80711, w_eco80712, w_eco80713, w_eco80714, w_eco80715, w_eco80716, w_eco80717, w_eco80718, w_eco80719, w_eco80720, w_eco80721, w_eco80722, w_eco80723, w_eco80724, w_eco80725, w_eco80726, w_eco80727, w_eco80728, w_eco80729, w_eco80730, w_eco80731, w_eco80732, w_eco80733, w_eco80734, w_eco80735, w_eco80736, w_eco80737, w_eco80738, w_eco80739, w_eco80740, w_eco80741, w_eco80742, w_eco80743, w_eco80744, w_eco80745, w_eco80746, w_eco80747, w_eco80748, w_eco80749, w_eco80750, w_eco80751, w_eco80752, w_eco80753, w_eco80754, w_eco80755, w_eco80756, w_eco80757, w_eco80758, w_eco80759, w_eco80760, w_eco80761, w_eco80762, w_eco80763, w_eco80764, w_eco80765, w_eco80766, w_eco80767, w_eco80768, w_eco80769, w_eco80770, w_eco80771, w_eco80772, w_eco80773, w_eco80774, w_eco80775, w_eco80776, w_eco80777, w_eco80778, w_eco80779, w_eco80780, w_eco80781, w_eco80782, w_eco80783, w_eco80784, w_eco80785, w_eco80786, w_eco80787, w_eco80788, w_eco80789, w_eco80790, w_eco80791, w_eco80792, w_eco80793, w_eco80794, w_eco80795, w_eco80796, w_eco80797, w_eco80798, w_eco80799, w_eco80800, w_eco80801, w_eco80802, w_eco80803, w_eco80804, w_eco80805, w_eco80806, w_eco80807, w_eco80808, w_eco80809, w_eco80810, w_eco80811, w_eco80812, w_eco80813, w_eco80814, w_eco80815, w_eco80816, w_eco80817, w_eco80818, w_eco80819, w_eco80820, w_eco80821, w_eco80822, w_eco80823, w_eco80824, w_eco80825, w_eco80826, w_eco80827, w_eco80828, w_eco80829, w_eco80830, w_eco80831, w_eco80832, w_eco80833, w_eco80834, w_eco80835, w_eco80836, w_eco80837, w_eco80838, w_eco80839, w_eco80840, w_eco80841, w_eco80842, w_eco80843, w_eco80844, w_eco80845, w_eco80846, w_eco80847, w_eco80848, w_eco80849, w_eco80850, w_eco80851, w_eco80852, w_eco80853, w_eco80854, w_eco80855, w_eco80856, w_eco80857, w_eco80858, w_eco80859, w_eco80860, w_eco80861, w_eco80862, w_eco80863, w_eco80864, w_eco80865, w_eco80866, w_eco80867, w_eco80868, w_eco80869, w_eco80870, w_eco80871, w_eco80872, w_eco80873, w_eco80874, w_eco80875, w_eco80876, w_eco80877, w_eco80878, w_eco80879, w_eco80880, w_eco80881, w_eco80882, w_eco80883, w_eco80884, w_eco80885, w_eco80886, w_eco80887, w_eco80888, w_eco80889, w_eco80890, w_eco80891, w_eco80892, w_eco80893, w_eco80894, w_eco80895, w_eco80896, w_eco80897, w_eco80898, w_eco80899, w_eco80900, w_eco80901, w_eco80902, w_eco80903, w_eco80904, w_eco80905, w_eco80906, w_eco80907, w_eco80908, w_eco80909, w_eco80910, w_eco80911, w_eco80912, w_eco80913, w_eco80914, w_eco80915, w_eco80916, w_eco80917, w_eco80918, w_eco80919, w_eco80920, w_eco80921, w_eco80922, w_eco80923, w_eco80924, w_eco80925, w_eco80926, w_eco80927, w_eco80928, w_eco80929, w_eco80930, w_eco80931, w_eco80932, w_eco80933, w_eco80934, w_eco80935, w_eco80936, w_eco80937, w_eco80938, w_eco80939, w_eco80940, w_eco80941, w_eco80942, w_eco80943, w_eco80944, w_eco80945, w_eco80946, w_eco80947, w_eco80948, w_eco80949, w_eco80950, w_eco80951, w_eco80952, w_eco80953, w_eco80954, w_eco80955, w_eco80956, w_eco80957, w_eco80958, w_eco80959, w_eco80960, w_eco80961, w_eco80962, w_eco80963, w_eco80964, w_eco80965, w_eco80966, w_eco80967, w_eco80968, w_eco80969, w_eco80970, w_eco80971, w_eco80972, w_eco80973, w_eco80974, w_eco80975, w_eco80976, w_eco80977, w_eco80978, w_eco80979, w_eco80980, w_eco80981, w_eco80982, w_eco80983, w_eco80984, w_eco80985, w_eco80986, w_eco80987, w_eco80988, w_eco80989, w_eco80990, w_eco80991, w_eco80992, w_eco80993, w_eco80994, w_eco80995, w_eco80996, w_eco80997, w_eco80998, w_eco80999, w_eco81000, w_eco81001, w_eco81002, w_eco81003, w_eco81004, w_eco81005, w_eco81006, w_eco81007, w_eco81008, w_eco81009, w_eco81010, w_eco81011, w_eco81012, w_eco81013, w_eco81014, w_eco81015, w_eco81016, w_eco81017, w_eco81018, w_eco81019, w_eco81020, w_eco81021, w_eco81022, w_eco81023, w_eco81024, w_eco81025, w_eco81026, w_eco81027, w_eco81028, w_eco81029, w_eco81030, w_eco81031, w_eco81032, w_eco81033, w_eco81034, w_eco81035, w_eco81036, w_eco81037, w_eco81038, w_eco81039, w_eco81040, w_eco81041, w_eco81042, w_eco81043, w_eco81044, w_eco81045, w_eco81046, w_eco81047, w_eco81048, w_eco81049, w_eco81050, w_eco81051, w_eco81052, w_eco81053, w_eco81054, w_eco81055, w_eco81056, w_eco81057, w_eco81058, w_eco81059, w_eco81060, w_eco81061, w_eco81062, w_eco81063, w_eco81064, w_eco81065, w_eco81066, w_eco81067, w_eco81068, w_eco81069, w_eco81070, w_eco81071, w_eco81072, w_eco81073, w_eco81074, w_eco81075, w_eco81076, w_eco81077, w_eco81078, w_eco81079, w_eco81080, w_eco81081, w_eco81082, w_eco81083, w_eco81084, w_eco81085, w_eco81086, w_eco81087, w_eco81088, w_eco81089, w_eco81090, w_eco81091, w_eco81092, w_eco81093, w_eco81094, w_eco81095, w_eco81096, w_eco81097, w_eco81098, w_eco81099, w_eco81100, w_eco81101, w_eco81102, w_eco81103, w_eco81104, w_eco81105, w_eco81106, w_eco81107, w_eco81108, w_eco81109, w_eco81110, w_eco81111, w_eco81112, w_eco81113, w_eco81114, w_eco81115, w_eco81116, w_eco81117, w_eco81118, w_eco81119, w_eco81120, w_eco81121, w_eco81122, w_eco81123, w_eco81124, w_eco81125, w_eco81126, w_eco81127, w_eco81128, w_eco81129, w_eco81130, w_eco81131, w_eco81132, w_eco81133, w_eco81134, w_eco81135, w_eco81136, w_eco81137, w_eco81138, w_eco81139, w_eco81140, w_eco81141, w_eco81142, w_eco81143, w_eco81144, w_eco81145, w_eco81146, w_eco81147, w_eco81148, w_eco81149, w_eco81150, w_eco81151, w_eco81152, w_eco81153, w_eco81154, w_eco81155, w_eco81156, w_eco81157, w_eco81158, w_eco81159, w_eco81160, w_eco81161, w_eco81162, w_eco81163, w_eco81164, w_eco81165, w_eco81166, w_eco81167, w_eco81168, w_eco81169, w_eco81170, w_eco81171, w_eco81172, w_eco81173, w_eco81174, w_eco81175, w_eco81176, w_eco81177, w_eco81178, w_eco81179, w_eco81180, w_eco81181, w_eco81182, w_eco81183, w_eco81184, w_eco81185, w_eco81186, w_eco81187, w_eco81188, w_eco81189, w_eco81190, w_eco81191, w_eco81192, w_eco81193, w_eco81194, w_eco81195, w_eco81196, w_eco81197, w_eco81198, w_eco81199, w_eco81200, w_eco81201, w_eco81202, w_eco81203, w_eco81204, w_eco81205, w_eco81206, w_eco81207, w_eco81208, w_eco81209, w_eco81210, w_eco81211, w_eco81212, w_eco81213, w_eco81214, w_eco81215, w_eco81216, w_eco81217, w_eco81218, w_eco81219, w_eco81220, w_eco81221, w_eco81222, w_eco81223, w_eco81224, w_eco81225, w_eco81226, w_eco81227, w_eco81228, w_eco81229, w_eco81230, w_eco81231, w_eco81232, w_eco81233, w_eco81234, w_eco81235, w_eco81236, w_eco81237, w_eco81238, w_eco81239, w_eco81240, w_eco81241, w_eco81242, w_eco81243, w_eco81244, w_eco81245, w_eco81246, w_eco81247, w_eco81248, w_eco81249, w_eco81250, w_eco81251, w_eco81252, w_eco81253, w_eco81254, w_eco81255, w_eco81256, w_eco81257, w_eco81258, w_eco81259, w_eco81260, w_eco81261, w_eco81262, w_eco81263, w_eco81264, w_eco81265, w_eco81266, w_eco81267, w_eco81268, w_eco81269, w_eco81270, w_eco81271, w_eco81272, w_eco81273, w_eco81274, w_eco81275, w_eco81276, w_eco81277, w_eco81278, w_eco81279, w_eco81280, w_eco81281, w_eco81282, w_eco81283, w_eco81284, w_eco81285, w_eco81286, w_eco81287, w_eco81288, w_eco81289, w_eco81290, w_eco81291, w_eco81292, w_eco81293, w_eco81294, w_eco81295, w_eco81296, w_eco81297, w_eco81298, w_eco81299, w_eco81300, w_eco81301, w_eco81302, w_eco81303, w_eco81304, w_eco81305, w_eco81306, w_eco81307, w_eco81308, w_eco81309, w_eco81310, w_eco81311, w_eco81312, w_eco81313, w_eco81314, w_eco81315, w_eco81316, w_eco81317, w_eco81318, w_eco81319, w_eco81320, w_eco81321, w_eco81322, w_eco81323, w_eco81324, w_eco81325, w_eco81326, w_eco81327, w_eco81328, w_eco81329, w_eco81330, w_eco81331, w_eco81332, w_eco81333, w_eco81334, w_eco81335, w_eco81336, w_eco81337, w_eco81338, w_eco81339, w_eco81340, w_eco81341, w_eco81342, w_eco81343, w_eco81344, w_eco81345, w_eco81346, w_eco81347, w_eco81348, w_eco81349, w_eco81350, w_eco81351, w_eco81352, w_eco81353, w_eco81354, w_eco81355, w_eco81356, w_eco81357, w_eco81358, w_eco81359, w_eco81360, w_eco81361, w_eco81362, w_eco81363, w_eco81364, w_eco81365, w_eco81366, w_eco81367, w_eco81368, w_eco81369, w_eco81370, w_eco81371, w_eco81372, w_eco81373, w_eco81374, w_eco81375, w_eco81376, w_eco81377, w_eco81378, w_eco81379, w_eco81380, w_eco81381, w_eco81382, w_eco81383, w_eco81384, w_eco81385, w_eco81386, w_eco81387, w_eco81388, w_eco81389, w_eco81390, w_eco81391, w_eco81392, w_eco81393, w_eco81394, w_eco81395, w_eco81396, w_eco81397, w_eco81398, w_eco81399, w_eco81400, w_eco81401, w_eco81402, w_eco81403, w_eco81404, w_eco81405, w_eco81406, w_eco81407, w_eco81408, w_eco81409, w_eco81410, w_eco81411, w_eco81412, w_eco81413, w_eco81414, w_eco81415, w_eco81416, w_eco81417, w_eco81418, w_eco81419, w_eco81420, w_eco81421, w_eco81422, w_eco81423, w_eco81424, w_eco81425, w_eco81426, w_eco81427, w_eco81428, w_eco81429, w_eco81430, w_eco81431, w_eco81432, w_eco81433, w_eco81434, w_eco81435, w_eco81436, w_eco81437, w_eco81438, w_eco81439, w_eco81440, w_eco81441, w_eco81442, w_eco81443, w_eco81444, w_eco81445, w_eco81446, w_eco81447, w_eco81448, w_eco81449, w_eco81450, w_eco81451, w_eco81452, w_eco81453, w_eco81454, w_eco81455, w_eco81456, w_eco81457, w_eco81458, w_eco81459, w_eco81460, w_eco81461, w_eco81462, w_eco81463, w_eco81464, w_eco81465, w_eco81466, w_eco81467, w_eco81468, w_eco81469, w_eco81470, w_eco81471, w_eco81472, w_eco81473, w_eco81474, w_eco81475, w_eco81476, w_eco81477, w_eco81478, w_eco81479, w_eco81480, w_eco81481, w_eco81482, w_eco81483, w_eco81484, w_eco81485, w_eco81486, w_eco81487, w_eco81488, w_eco81489, w_eco81490, w_eco81491, w_eco81492, w_eco81493, w_eco81494, w_eco81495, w_eco81496, w_eco81497, w_eco81498, w_eco81499, w_eco81500, w_eco81501, w_eco81502, w_eco81503, w_eco81504, w_eco81505, w_eco81506, w_eco81507, w_eco81508, w_eco81509, w_eco81510, w_eco81511, w_eco81512, w_eco81513, w_eco81514, w_eco81515, w_eco81516, w_eco81517, w_eco81518, w_eco81519, w_eco81520, w_eco81521, w_eco81522, w_eco81523, w_eco81524, w_eco81525, w_eco81526, w_eco81527, w_eco81528, w_eco81529, w_eco81530, w_eco81531, w_eco81532, w_eco81533, w_eco81534, w_eco81535, w_eco81536, w_eco81537, w_eco81538, w_eco81539, w_eco81540, w_eco81541, w_eco81542, w_eco81543, w_eco81544, w_eco81545, w_eco81546, w_eco81547, w_eco81548, w_eco81549, w_eco81550, w_eco81551, w_eco81552, w_eco81553, w_eco81554, w_eco81555, w_eco81556, w_eco81557, w_eco81558, w_eco81559, w_eco81560, w_eco81561, w_eco81562, w_eco81563, w_eco81564, w_eco81565, w_eco81566, w_eco81567, w_eco81568, w_eco81569, w_eco81570, w_eco81571, w_eco81572, w_eco81573, w_eco81574, w_eco81575, w_eco81576, w_eco81577, w_eco81578, w_eco81579, w_eco81580, w_eco81581, w_eco81582, w_eco81583, w_eco81584, w_eco81585, w_eco81586, w_eco81587, w_eco81588, w_eco81589, w_eco81590, w_eco81591, w_eco81592, w_eco81593, w_eco81594, w_eco81595, w_eco81596, w_eco81597, w_eco81598, w_eco81599, w_eco81600, w_eco81601, w_eco81602, w_eco81603, w_eco81604, w_eco81605, w_eco81606, w_eco81607, w_eco81608, w_eco81609, w_eco81610, w_eco81611, w_eco81612, w_eco81613, w_eco81614, w_eco81615, w_eco81616, w_eco81617, w_eco81618, w_eco81619, w_eco81620, w_eco81621, w_eco81622, w_eco81623, w_eco81624, w_eco81625, w_eco81626, w_eco81627, w_eco81628, w_eco81629, w_eco81630, w_eco81631, w_eco81632, w_eco81633, w_eco81634, w_eco81635, w_eco81636, w_eco81637, w_eco81638, w_eco81639, w_eco81640, w_eco81641, w_eco81642, w_eco81643, w_eco81644, w_eco81645, w_eco81646, w_eco81647, w_eco81648, w_eco81649, w_eco81650, w_eco81651, w_eco81652, w_eco81653, w_eco81654, w_eco81655, w_eco81656, w_eco81657, w_eco81658, w_eco81659, w_eco81660, w_eco81661, w_eco81662, w_eco81663, w_eco81664, w_eco81665, w_eco81666, w_eco81667, w_eco81668, w_eco81669, w_eco81670, w_eco81671, w_eco81672, w_eco81673, w_eco81674, w_eco81675, w_eco81676, w_eco81677, w_eco81678, w_eco81679, w_eco81680, w_eco81681, w_eco81682, w_eco81683, w_eco81684, w_eco81685, w_eco81686, w_eco81687, w_eco81688, w_eco81689, w_eco81690, w_eco81691, w_eco81692, w_eco81693, w_eco81694, w_eco81695, w_eco81696, w_eco81697, w_eco81698, w_eco81699, w_eco81700, w_eco81701, w_eco81702, w_eco81703, w_eco81704, w_eco81705, w_eco81706, w_eco81707, w_eco81708, w_eco81709, w_eco81710, w_eco81711, w_eco81712, w_eco81713, w_eco81714, w_eco81715, w_eco81716, w_eco81717, w_eco81718, w_eco81719, w_eco81720, w_eco81721, w_eco81722, w_eco81723, w_eco81724, w_eco81725, w_eco81726, w_eco81727, w_eco81728, w_eco81729, w_eco81730, w_eco81731, w_eco81732, w_eco81733, w_eco81734, w_eco81735, w_eco81736, w_eco81737, w_eco81738, w_eco81739, w_eco81740, w_eco81741, w_eco81742, w_eco81743, w_eco81744, w_eco81745, w_eco81746, w_eco81747, w_eco81748, w_eco81749, w_eco81750, w_eco81751, w_eco81752, w_eco81753, w_eco81754, w_eco81755, w_eco81756, w_eco81757, w_eco81758, w_eco81759, w_eco81760, w_eco81761, w_eco81762, w_eco81763, w_eco81764, w_eco81765, w_eco81766, w_eco81767, w_eco81768, w_eco81769, w_eco81770, w_eco81771, w_eco81772, w_eco81773, w_eco81774, w_eco81775, w_eco81776, w_eco81777, w_eco81778, w_eco81779, w_eco81780, w_eco81781, w_eco81782, w_eco81783, w_eco81784, w_eco81785, w_eco81786, w_eco81787, w_eco81788, w_eco81789, w_eco81790, w_eco81791, w_eco81792, w_eco81793, w_eco81794, w_eco81795, w_eco81796, w_eco81797, w_eco81798, w_eco81799, w_eco81800, w_eco81801, w_eco81802, w_eco81803, w_eco81804, w_eco81805, w_eco81806, w_eco81807, w_eco81808, w_eco81809, w_eco81810, w_eco81811, w_eco81812, w_eco81813, w_eco81814, w_eco81815, w_eco81816, w_eco81817, w_eco81818, w_eco81819, w_eco81820, w_eco81821, w_eco81822, w_eco81823, w_eco81824, w_eco81825, w_eco81826, w_eco81827, w_eco81828, w_eco81829, w_eco81830, w_eco81831, w_eco81832, w_eco81833, w_eco81834, w_eco81835, w_eco81836, w_eco81837, w_eco81838, w_eco81839, w_eco81840, w_eco81841, w_eco81842, w_eco81843, w_eco81844, w_eco81845, w_eco81846, w_eco81847, w_eco81848, w_eco81849, w_eco81850, w_eco81851, w_eco81852, w_eco81853, w_eco81854, w_eco81855, w_eco81856, w_eco81857, w_eco81858, w_eco81859, w_eco81860, w_eco81861, w_eco81862, w_eco81863, w_eco81864, w_eco81865, w_eco81866, w_eco81867, w_eco81868, w_eco81869, w_eco81870, w_eco81871, w_eco81872, w_eco81873, w_eco81874, w_eco81875, w_eco81876, w_eco81877, w_eco81878, w_eco81879, w_eco81880, w_eco81881, w_eco81882, w_eco81883, w_eco81884, w_eco81885, w_eco81886, w_eco81887, w_eco81888, w_eco81889, w_eco81890, w_eco81891, w_eco81892, w_eco81893, w_eco81894, w_eco81895, w_eco81896, w_eco81897, w_eco81898, w_eco81899, w_eco81900, w_eco81901, w_eco81902, w_eco81903, w_eco81904, w_eco81905, w_eco81906, w_eco81907, w_eco81908, w_eco81909, w_eco81910, w_eco81911, w_eco81912, w_eco81913, w_eco81914, w_eco81915, w_eco81916, w_eco81917, w_eco81918, w_eco81919, w_eco81920, w_eco81921, w_eco81922, w_eco81923, w_eco81924, w_eco81925, w_eco81926, w_eco81927, w_eco81928, w_eco81929, w_eco81930, w_eco81931, w_eco81932, w_eco81933, w_eco81934, w_eco81935, w_eco81936, w_eco81937, w_eco81938, w_eco81939, w_eco81940, w_eco81941, w_eco81942, w_eco81943, w_eco81944, w_eco81945, w_eco81946, w_eco81947, w_eco81948, w_eco81949, w_eco81950, w_eco81951, w_eco81952, w_eco81953, w_eco81954, w_eco81955, w_eco81956, w_eco81957, w_eco81958, w_eco81959, w_eco81960, w_eco81961, w_eco81962, w_eco81963, w_eco81964, w_eco81965, w_eco81966, w_eco81967, w_eco81968, w_eco81969, w_eco81970, w_eco81971, w_eco81972, w_eco81973, w_eco81974, w_eco81975, w_eco81976, w_eco81977, w_eco81978, w_eco81979, w_eco81980, w_eco81981, w_eco81982, w_eco81983, w_eco81984, w_eco81985, w_eco81986, w_eco81987, w_eco81988, w_eco81989, w_eco81990, w_eco81991, w_eco81992, w_eco81993, w_eco81994, w_eco81995, w_eco81996, w_eco81997, w_eco81998, w_eco81999, w_eco82000, w_eco82001, w_eco82002, w_eco82003, w_eco82004, w_eco82005, w_eco82006, w_eco82007, w_eco82008, w_eco82009, w_eco82010, w_eco82011, w_eco82012, w_eco82013, w_eco82014, w_eco82015, w_eco82016, w_eco82017, w_eco82018, w_eco82019, w_eco82020, w_eco82021, w_eco82022, w_eco82023, w_eco82024, w_eco82025, w_eco82026, w_eco82027, w_eco82028, w_eco82029, w_eco82030, w_eco82031, w_eco82032, w_eco82033, w_eco82034, w_eco82035, w_eco82036, w_eco82037, w_eco82038, w_eco82039, w_eco82040, w_eco82041, w_eco82042, w_eco82043, w_eco82044, w_eco82045, w_eco82046, w_eco82047, w_eco82048, w_eco82049, w_eco82050, w_eco82051, w_eco82052, w_eco82053, w_eco82054, w_eco82055, w_eco82056, w_eco82057, w_eco82058, w_eco82059, w_eco82060, w_eco82061, w_eco82062, w_eco82063, w_eco82064, w_eco82065, w_eco82066, w_eco82067, w_eco82068, w_eco82069, w_eco82070, w_eco82071, w_eco82072, w_eco82073, w_eco82074, w_eco82075, w_eco82076, w_eco82077, w_eco82078, w_eco82079, w_eco82080, w_eco82081, w_eco82082, w_eco82083, w_eco82084, w_eco82085, w_eco82086, w_eco82087, w_eco82088, w_eco82089, w_eco82090, w_eco82091, w_eco82092, w_eco82093, w_eco82094, w_eco82095, w_eco82096, w_eco82097, w_eco82098, w_eco82099, w_eco82100, w_eco82101, w_eco82102, w_eco82103, w_eco82104, w_eco82105, w_eco82106, w_eco82107, w_eco82108, w_eco82109, w_eco82110, w_eco82111, w_eco82112, w_eco82113, w_eco82114, w_eco82115, w_eco82116, w_eco82117, w_eco82118, w_eco82119, w_eco82120, w_eco82121, w_eco82122, w_eco82123, w_eco82124, w_eco82125, w_eco82126, w_eco82127, w_eco82128, w_eco82129, w_eco82130, w_eco82131, w_eco82132, w_eco82133, w_eco82134, w_eco82135, w_eco82136, w_eco82137, w_eco82138, w_eco82139, w_eco82140, w_eco82141, w_eco82142, w_eco82143, w_eco82144, w_eco82145, w_eco82146, w_eco82147, w_eco82148, w_eco82149, w_eco82150, w_eco82151, w_eco82152, w_eco82153, w_eco82154, w_eco82155, w_eco82156, w_eco82157, w_eco82158, w_eco82159, w_eco82160, w_eco82161, w_eco82162, w_eco82163, w_eco82164, w_eco82165, w_eco82166, w_eco82167, w_eco82168, w_eco82169, w_eco82170, w_eco82171, w_eco82172, w_eco82173, w_eco82174, w_eco82175, w_eco82176, w_eco82177, w_eco82178, w_eco82179, w_eco82180, w_eco82181, w_eco82182, w_eco82183, w_eco82184, w_eco82185, w_eco82186, w_eco82187, w_eco82188, w_eco82189, w_eco82190, w_eco82191, w_eco82192, w_eco82193, w_eco82194, w_eco82195, w_eco82196, w_eco82197, w_eco82198, w_eco82199, w_eco82200, w_eco82201, w_eco82202, w_eco82203, w_eco82204, w_eco82205, w_eco82206, w_eco82207, w_eco82208, w_eco82209, w_eco82210, w_eco82211, w_eco82212, w_eco82213, w_eco82214, w_eco82215, w_eco82216, w_eco82217, w_eco82218, w_eco82219, w_eco82220, w_eco82221, w_eco82222, w_eco82223, w_eco82224, w_eco82225, w_eco82226, w_eco82227, w_eco82228, w_eco82229, w_eco82230, w_eco82231, w_eco82232, w_eco82233, w_eco82234, w_eco82235, w_eco82236, w_eco82237, w_eco82238, w_eco82239, w_eco82240, w_eco82241, w_eco82242, w_eco82243, w_eco82244, w_eco82245, w_eco82246, w_eco82247, w_eco82248, w_eco82249, w_eco82250, w_eco82251, w_eco82252, w_eco82253, w_eco82254, w_eco82255, w_eco82256, w_eco82257, w_eco82258, w_eco82259, w_eco82260, w_eco82261, w_eco82262, w_eco82263, w_eco82264, w_eco82265, w_eco82266, w_eco82267, w_eco82268, w_eco82269, w_eco82270, w_eco82271, w_eco82272, w_eco82273, w_eco82274, w_eco82275, w_eco82276, w_eco82277, w_eco82278, w_eco82279, w_eco82280, w_eco82281, w_eco82282, w_eco82283, w_eco82284, w_eco82285, w_eco82286, w_eco82287, w_eco82288, w_eco82289, w_eco82290, w_eco82291, w_eco82292, w_eco82293, w_eco82294, w_eco82295, w_eco82296, w_eco82297, w_eco82298, w_eco82299, w_eco82300, w_eco82301, w_eco82302, w_eco82303, w_eco82304, w_eco82305, w_eco82306, w_eco82307, w_eco82308, w_eco82309, w_eco82310, w_eco82311, w_eco82312, w_eco82313, w_eco82314, w_eco82315, w_eco82316, w_eco82317, w_eco82318, w_eco82319, w_eco82320, w_eco82321, w_eco82322, w_eco82323, w_eco82324, w_eco82325, w_eco82326, w_eco82327, w_eco82328, w_eco82329, w_eco82330, w_eco82331, w_eco82332, w_eco82333, w_eco82334, w_eco82335, w_eco82336, w_eco82337, w_eco82338, w_eco82339, w_eco82340, w_eco82341, w_eco82342, w_eco82343, w_eco82344, w_eco82345, w_eco82346, w_eco82347, w_eco82348, w_eco82349, w_eco82350, w_eco82351, w_eco82352, w_eco82353, w_eco82354, w_eco82355, w_eco82356, w_eco82357, w_eco82358, w_eco82359, w_eco82360, w_eco82361, w_eco82362, w_eco82363, w_eco82364, w_eco82365, w_eco82366, w_eco82367, w_eco82368, w_eco82369, w_eco82370, w_eco82371, w_eco82372, w_eco82373, w_eco82374, w_eco82375, w_eco82376, w_eco82377, w_eco82378, w_eco82379, w_eco82380, w_eco82381, w_eco82382, w_eco82383, w_eco82384, w_eco82385, w_eco82386, w_eco82387, w_eco82388, w_eco82389, w_eco82390, w_eco82391, w_eco82392, w_eco82393, w_eco82394, w_eco82395, w_eco82396, w_eco82397, w_eco82398, w_eco82399, w_eco82400, w_eco82401, w_eco82402, w_eco82403, w_eco82404, w_eco82405, w_eco82406, w_eco82407, w_eco82408, w_eco82409, w_eco82410, w_eco82411, w_eco82412, w_eco82413, w_eco82414, w_eco82415, w_eco82416, w_eco82417, w_eco82418, w_eco82419, w_eco82420, w_eco82421, w_eco82422, w_eco82423, w_eco82424, w_eco82425, w_eco82426, w_eco82427, w_eco82428, w_eco82429, w_eco82430, w_eco82431, w_eco82432, w_eco82433, w_eco82434, w_eco82435, w_eco82436, w_eco82437, w_eco82438, w_eco82439, w_eco82440, w_eco82441, w_eco82442, w_eco82443, w_eco82444, w_eco82445, w_eco82446, w_eco82447, w_eco82448, w_eco82449, w_eco82450, w_eco82451, w_eco82452, w_eco82453, w_eco82454, w_eco82455, w_eco82456, w_eco82457, w_eco82458, w_eco82459, w_eco82460, w_eco82461, w_eco82462, w_eco82463, w_eco82464, w_eco82465, w_eco82466, w_eco82467, w_eco82468, w_eco82469, w_eco82470, w_eco82471, w_eco82472, w_eco82473, w_eco82474, w_eco82475, w_eco82476, w_eco82477, w_eco82478, w_eco82479, w_eco82480, w_eco82481, w_eco82482, w_eco82483, w_eco82484, w_eco82485, w_eco82486, w_eco82487, w_eco82488, w_eco82489, w_eco82490, w_eco82491, w_eco82492, w_eco82493, w_eco82494, w_eco82495, w_eco82496, w_eco82497, w_eco82498, w_eco82499, w_eco82500, w_eco82501, w_eco82502, w_eco82503, w_eco82504, w_eco82505, w_eco82506, w_eco82507, w_eco82508, w_eco82509, w_eco82510, w_eco82511, w_eco82512, w_eco82513, w_eco82514, w_eco82515, w_eco82516, w_eco82517, w_eco82518, w_eco82519, w_eco82520, w_eco82521, w_eco82522, w_eco82523, w_eco82524, w_eco82525, w_eco82526, w_eco82527, w_eco82528, w_eco82529, w_eco82530, w_eco82531, w_eco82532, w_eco82533, w_eco82534, w_eco82535, w_eco82536, w_eco82537, w_eco82538, w_eco82539, w_eco82540, w_eco82541, w_eco82542, w_eco82543, w_eco82544, w_eco82545, w_eco82546, w_eco82547, w_eco82548, w_eco82549, w_eco82550, w_eco82551, w_eco82552, w_eco82553, w_eco82554, w_eco82555, w_eco82556, w_eco82557, w_eco82558, w_eco82559, w_eco82560, w_eco82561, w_eco82562, w_eco82563, w_eco82564, w_eco82565, w_eco82566, w_eco82567, w_eco82568, w_eco82569, w_eco82570, w_eco82571, w_eco82572, w_eco82573, w_eco82574, w_eco82575, w_eco82576, w_eco82577, w_eco82578, w_eco82579, w_eco82580, w_eco82581, w_eco82582, w_eco82583, w_eco82584, w_eco82585, w_eco82586, w_eco82587, w_eco82588, w_eco82589, w_eco82590, w_eco82591, w_eco82592, w_eco82593, w_eco82594, w_eco82595, w_eco82596, w_eco82597, w_eco82598, w_eco82599, w_eco82600, w_eco82601, w_eco82602, w_eco82603, w_eco82604, w_eco82605, w_eco82606, w_eco82607, w_eco82608, w_eco82609, w_eco82610, w_eco82611, w_eco82612, w_eco82613, w_eco82614, w_eco82615, w_eco82616, w_eco82617, w_eco82618, w_eco82619, w_eco82620, w_eco82621, w_eco82622, w_eco82623, w_eco82624, w_eco82625, w_eco82626, w_eco82627, w_eco82628, w_eco82629, w_eco82630, w_eco82631, w_eco82632, w_eco82633, w_eco82634, w_eco82635, w_eco82636, w_eco82637, w_eco82638, w_eco82639, w_eco82640, w_eco82641, w_eco82642, w_eco82643, w_eco82644, w_eco82645, w_eco82646, w_eco82647, w_eco82648, w_eco82649, w_eco82650, w_eco82651, w_eco82652, w_eco82653, w_eco82654, w_eco82655, w_eco82656, w_eco82657, w_eco82658, w_eco82659, w_eco82660, w_eco82661, w_eco82662, w_eco82663, w_eco82664, w_eco82665, w_eco82666, w_eco82667, w_eco82668, w_eco82669, w_eco82670, w_eco82671, w_eco82672, w_eco82673, w_eco82674, w_eco82675, w_eco82676, w_eco82677, w_eco82678, w_eco82679, w_eco82680, w_eco82681, w_eco82682, w_eco82683, w_eco82684, w_eco82685, w_eco82686, w_eco82687, w_eco82688, w_eco82689, w_eco82690, w_eco82691, w_eco82692, w_eco82693, w_eco82694, w_eco82695, w_eco82696, w_eco82697, w_eco82698, w_eco82699, w_eco82700, w_eco82701, w_eco82702, w_eco82703, w_eco82704, w_eco82705, w_eco82706, w_eco82707, w_eco82708, w_eco82709, w_eco82710, w_eco82711, w_eco82712, w_eco82713, w_eco82714, w_eco82715, w_eco82716, w_eco82717, w_eco82718, w_eco82719, w_eco82720, w_eco82721, w_eco82722, w_eco82723, w_eco82724, w_eco82725, w_eco82726, w_eco82727, w_eco82728, w_eco82729, w_eco82730, w_eco82731, w_eco82732, w_eco82733, w_eco82734, w_eco82735, w_eco82736, w_eco82737, w_eco82738, w_eco82739, w_eco82740, w_eco82741, w_eco82742, w_eco82743, w_eco82744, w_eco82745, w_eco82746, w_eco82747, w_eco82748, w_eco82749, w_eco82750, w_eco82751, w_eco82752, w_eco82753, w_eco82754, w_eco82755, w_eco82756, w_eco82757, w_eco82758, w_eco82759, w_eco82760, w_eco82761, w_eco82762, w_eco82763, w_eco82764, w_eco82765, w_eco82766, w_eco82767, w_eco82768, w_eco82769, w_eco82770, w_eco82771, w_eco82772, w_eco82773, w_eco82774, w_eco82775, w_eco82776, w_eco82777, w_eco82778, w_eco82779, w_eco82780, w_eco82781, w_eco82782, w_eco82783, w_eco82784, w_eco82785, w_eco82786, w_eco82787, w_eco82788, w_eco82789, w_eco82790, w_eco82791, w_eco82792, w_eco82793, w_eco82794, w_eco82795, w_eco82796, w_eco82797, w_eco82798, w_eco82799, w_eco82800, w_eco82801, w_eco82802, w_eco82803, w_eco82804, w_eco82805, w_eco82806, w_eco82807, w_eco82808, w_eco82809, w_eco82810, w_eco82811, w_eco82812, w_eco82813, w_eco82814, w_eco82815, w_eco82816, w_eco82817, w_eco82818, w_eco82819, w_eco82820, w_eco82821, w_eco82822, w_eco82823, w_eco82824, w_eco82825, w_eco82826, w_eco82827, w_eco82828, w_eco82829, w_eco82830, w_eco82831, w_eco82832, w_eco82833, w_eco82834, w_eco82835, w_eco82836, w_eco82837, w_eco82838, w_eco82839, w_eco82840, w_eco82841, w_eco82842, w_eco82843, w_eco82844, w_eco82845, w_eco82846, w_eco82847, w_eco82848, w_eco82849, w_eco82850, w_eco82851, w_eco82852, w_eco82853, w_eco82854, w_eco82855, w_eco82856, w_eco82857, w_eco82858, w_eco82859, w_eco82860, w_eco82861, w_eco82862, w_eco82863, w_eco82864, w_eco82865, w_eco82866, w_eco82867, w_eco82868, w_eco82869, w_eco82870, w_eco82871, w_eco82872, w_eco82873, w_eco82874, w_eco82875, w_eco82876, w_eco82877, w_eco82878, w_eco82879, w_eco82880, w_eco82881, w_eco82882, w_eco82883, w_eco82884, w_eco82885, w_eco82886, w_eco82887, w_eco82888, w_eco82889, w_eco82890, w_eco82891, w_eco82892, w_eco82893, w_eco82894, w_eco82895, w_eco82896, w_eco82897, w_eco82898, w_eco82899, w_eco82900, w_eco82901, w_eco82902, w_eco82903, w_eco82904, w_eco82905, w_eco82906, w_eco82907, w_eco82908, w_eco82909, w_eco82910, w_eco82911, w_eco82912, w_eco82913, w_eco82914, w_eco82915, w_eco82916, w_eco82917, w_eco82918, w_eco82919, w_eco82920, w_eco82921, w_eco82922, w_eco82923, w_eco82924, w_eco82925, w_eco82926, w_eco82927, w_eco82928, w_eco82929, w_eco82930, w_eco82931, w_eco82932, w_eco82933, w_eco82934, w_eco82935, w_eco82936, w_eco82937, w_eco82938, w_eco82939, w_eco82940, w_eco82941, w_eco82942, w_eco82943, w_eco82944, w_eco82945, w_eco82946, w_eco82947, w_eco82948, w_eco82949, w_eco82950, w_eco82951, w_eco82952, w_eco82953, w_eco82954, w_eco82955, w_eco82956, w_eco82957, w_eco82958, w_eco82959, w_eco82960, w_eco82961, w_eco82962, w_eco82963, w_eco82964, w_eco82965, w_eco82966, w_eco82967, w_eco82968, w_eco82969, w_eco82970, w_eco82971, w_eco82972, w_eco82973, w_eco82974, w_eco82975, w_eco82976, w_eco82977, w_eco82978, w_eco82979, w_eco82980, w_eco82981, w_eco82982, w_eco82983, w_eco82984, w_eco82985, w_eco82986, w_eco82987, w_eco82988, w_eco82989, w_eco82990, w_eco82991, w_eco82992, w_eco82993, w_eco82994, w_eco82995, w_eco82996, w_eco82997, w_eco82998, w_eco82999, w_eco83000, w_eco83001, w_eco83002, w_eco83003, w_eco83004, w_eco83005, w_eco83006, w_eco83007, w_eco83008, w_eco83009, w_eco83010, w_eco83011, w_eco83012, w_eco83013, w_eco83014, w_eco83015, w_eco83016, w_eco83017, w_eco83018, w_eco83019, w_eco83020, w_eco83021, w_eco83022, w_eco83023, w_eco83024, w_eco83025, w_eco83026, w_eco83027, w_eco83028, w_eco83029, w_eco83030, w_eco83031, w_eco83032, w_eco83033, w_eco83034, w_eco83035, w_eco83036, w_eco83037, w_eco83038, w_eco83039, w_eco83040, w_eco83041, w_eco83042, w_eco83043, w_eco83044, w_eco83045, w_eco83046, w_eco83047, w_eco83048, w_eco83049, w_eco83050, w_eco83051, w_eco83052, w_eco83053, w_eco83054, w_eco83055, w_eco83056, w_eco83057, w_eco83058, w_eco83059, w_eco83060, w_eco83061, w_eco83062, w_eco83063, w_eco83064, w_eco83065, w_eco83066, w_eco83067, w_eco83068, w_eco83069, w_eco83070, w_eco83071, w_eco83072, w_eco83073, w_eco83074, w_eco83075, w_eco83076, w_eco83077, w_eco83078, w_eco83079, w_eco83080, w_eco83081, w_eco83082, w_eco83083, w_eco83084, w_eco83085, w_eco83086, w_eco83087, w_eco83088, w_eco83089, w_eco83090, w_eco83091, w_eco83092, w_eco83093, w_eco83094, w_eco83095, w_eco83096, w_eco83097, w_eco83098, w_eco83099, w_eco83100, w_eco83101, w_eco83102, w_eco83103, w_eco83104, w_eco83105, w_eco83106, w_eco83107, w_eco83108, w_eco83109, w_eco83110, w_eco83111, w_eco83112, w_eco83113, w_eco83114, w_eco83115, w_eco83116, w_eco83117, w_eco83118, w_eco83119, w_eco83120, w_eco83121, w_eco83122, w_eco83123, w_eco83124, w_eco83125, w_eco83126, w_eco83127, w_eco83128, w_eco83129, w_eco83130, w_eco83131, w_eco83132, w_eco83133, w_eco83134, w_eco83135, w_eco83136, w_eco83137, w_eco83138, w_eco83139, w_eco83140, w_eco83141, w_eco83142, w_eco83143, w_eco83144, w_eco83145, w_eco83146, w_eco83147, w_eco83148, w_eco83149, w_eco83150, w_eco83151, w_eco83152, w_eco83153, w_eco83154, w_eco83155, w_eco83156, w_eco83157, w_eco83158, w_eco83159, w_eco83160, w_eco83161, w_eco83162, w_eco83163, w_eco83164, w_eco83165, w_eco83166, w_eco83167, w_eco83168, w_eco83169, w_eco83170, w_eco83171, w_eco83172, w_eco83173, w_eco83174, w_eco83175, w_eco83176, w_eco83177, w_eco83178, w_eco83179, w_eco83180, w_eco83181, w_eco83182, w_eco83183, w_eco83184, w_eco83185, w_eco83186, w_eco83187, w_eco83188, w_eco83189, w_eco83190, w_eco83191, w_eco83192, w_eco83193, w_eco83194, w_eco83195, w_eco83196, w_eco83197, w_eco83198, w_eco83199, w_eco83200, w_eco83201, w_eco83202, w_eco83203, w_eco83204, w_eco83205, w_eco83206, w_eco83207, w_eco83208, w_eco83209, w_eco83210, w_eco83211, w_eco83212, w_eco83213, w_eco83214, w_eco83215, w_eco83216, w_eco83217, w_eco83218, w_eco83219, w_eco83220, w_eco83221, w_eco83222, w_eco83223, w_eco83224, w_eco83225, w_eco83226, w_eco83227, w_eco83228, w_eco83229, w_eco83230, w_eco83231, w_eco83232, w_eco83233, w_eco83234, w_eco83235, w_eco83236, w_eco83237, w_eco83238, w_eco83239, w_eco83240, w_eco83241, w_eco83242, w_eco83243, w_eco83244, w_eco83245, w_eco83246, w_eco83247, w_eco83248, w_eco83249, w_eco83250, w_eco83251, w_eco83252, w_eco83253, w_eco83254, w_eco83255, w_eco83256, w_eco83257, w_eco83258, w_eco83259, w_eco83260, w_eco83261, w_eco83262, w_eco83263, w_eco83264, w_eco83265, w_eco83266, w_eco83267, w_eco83268, w_eco83269, w_eco83270, w_eco83271, w_eco83272, w_eco83273, w_eco83274, w_eco83275, w_eco83276, w_eco83277, w_eco83278, w_eco83279, w_eco83280, w_eco83281, w_eco83282, w_eco83283, w_eco83284, w_eco83285, w_eco83286, w_eco83287, w_eco83288, w_eco83289, w_eco83290, w_eco83291, w_eco83292, w_eco83293, w_eco83294, w_eco83295, w_eco83296, w_eco83297, w_eco83298, w_eco83299, w_eco83300, w_eco83301, w_eco83302, w_eco83303, w_eco83304, w_eco83305, w_eco83306, w_eco83307, w_eco83308, w_eco83309, w_eco83310, w_eco83311, w_eco83312, w_eco83313, w_eco83314, w_eco83315, w_eco83316, w_eco83317, w_eco83318, w_eco83319, w_eco83320, w_eco83321, w_eco83322, w_eco83323, w_eco83324, w_eco83325, w_eco83326, w_eco83327, w_eco83328, w_eco83329, w_eco83330, w_eco83331, w_eco83332, w_eco83333, w_eco83334, w_eco83335, w_eco83336, w_eco83337, w_eco83338, w_eco83339, w_eco83340, w_eco83341, w_eco83342, w_eco83343, w_eco83344, w_eco83345, w_eco83346, w_eco83347, w_eco83348, w_eco83349, w_eco83350, w_eco83351, w_eco83352, w_eco83353, w_eco83354, w_eco83355, w_eco83356, w_eco83357, w_eco83358, w_eco83359, w_eco83360, w_eco83361, w_eco83362, w_eco83363, w_eco83364, w_eco83365, w_eco83366, w_eco83367, w_eco83368, w_eco83369, w_eco83370, w_eco83371, w_eco83372, w_eco83373, w_eco83374, w_eco83375, w_eco83376, w_eco83377, w_eco83378, w_eco83379, w_eco83380, w_eco83381, w_eco83382, w_eco83383, w_eco83384, w_eco83385, w_eco83386, w_eco83387, w_eco83388, w_eco83389, w_eco83390, w_eco83391, w_eco83392, w_eco83393, w_eco83394, w_eco83395, w_eco83396, w_eco83397, w_eco83398, w_eco83399, w_eco83400, w_eco83401, w_eco83402, w_eco83403, w_eco83404, w_eco83405, w_eco83406, w_eco83407, w_eco83408, w_eco83409, w_eco83410, w_eco83411, w_eco83412, w_eco83413, w_eco83414, w_eco83415, w_eco83416, w_eco83417, w_eco83418, w_eco83419, w_eco83420, w_eco83421, w_eco83422, w_eco83423, w_eco83424, w_eco83425, w_eco83426, w_eco83427, w_eco83428, w_eco83429, w_eco83430, w_eco83431, w_eco83432, w_eco83433, w_eco83434, w_eco83435, w_eco83436, w_eco83437, w_eco83438, w_eco83439, w_eco83440, w_eco83441, w_eco83442, w_eco83443, w_eco83444, w_eco83445, w_eco83446, w_eco83447, w_eco83448, w_eco83449, w_eco83450, w_eco83451, w_eco83452, w_eco83453, w_eco83454, w_eco83455, w_eco83456, w_eco83457, w_eco83458, w_eco83459, w_eco83460, w_eco83461, w_eco83462, w_eco83463, w_eco83464, w_eco83465, w_eco83466, w_eco83467, w_eco83468, w_eco83469, w_eco83470, w_eco83471, w_eco83472, w_eco83473, w_eco83474, w_eco83475, w_eco83476, w_eco83477, w_eco83478, w_eco83479, w_eco83480, w_eco83481, w_eco83482, w_eco83483, w_eco83484, w_eco83485, w_eco83486, w_eco83487, w_eco83488, w_eco83489, w_eco83490, w_eco83491, w_eco83492, w_eco83493, w_eco83494, w_eco83495, w_eco83496, w_eco83497, w_eco83498, w_eco83499, w_eco83500, w_eco83501, w_eco83502, w_eco83503, w_eco83504, w_eco83505, w_eco83506, w_eco83507, w_eco83508, w_eco83509, w_eco83510, w_eco83511, w_eco83512, w_eco83513, w_eco83514, w_eco83515, w_eco83516, w_eco83517, w_eco83518, w_eco83519, w_eco83520, w_eco83521, w_eco83522, w_eco83523, w_eco83524, w_eco83525, w_eco83526, w_eco83527, w_eco83528, w_eco83529, w_eco83530, w_eco83531, w_eco83532, w_eco83533, w_eco83534, w_eco83535, w_eco83536, w_eco83537, w_eco83538, w_eco83539, w_eco83540, w_eco83541, w_eco83542, w_eco83543, w_eco83544, w_eco83545, w_eco83546, w_eco83547, w_eco83548, w_eco83549, w_eco83550, w_eco83551, w_eco83552, w_eco83553, w_eco83554, w_eco83555, w_eco83556, w_eco83557, w_eco83558, w_eco83559, w_eco83560, w_eco83561, w_eco83562, w_eco83563, w_eco83564, w_eco83565, w_eco83566, w_eco83567, w_eco83568, w_eco83569, w_eco83570, w_eco83571, w_eco83572, w_eco83573, w_eco83574, w_eco83575, w_eco83576, w_eco83577, w_eco83578, w_eco83579, w_eco83580, w_eco83581, w_eco83582, w_eco83583, w_eco83584, w_eco83585, w_eco83586, w_eco83587, w_eco83588, w_eco83589, w_eco83590, w_eco83591, w_eco83592, w_eco83593, w_eco83594, w_eco83595, w_eco83596, w_eco83597, w_eco83598, w_eco83599, w_eco83600, w_eco83601, w_eco83602, w_eco83603, w_eco83604, w_eco83605, w_eco83606, w_eco83607, w_eco83608, w_eco83609, w_eco83610, w_eco83611, w_eco83612, w_eco83613, w_eco83614, w_eco83615, w_eco83616, w_eco83617, w_eco83618, w_eco83619, w_eco83620, w_eco83621, w_eco83622, w_eco83623, w_eco83624, w_eco83625, w_eco83626, w_eco83627, w_eco83628, w_eco83629, w_eco83630, w_eco83631, w_eco83632, w_eco83633, w_eco83634, w_eco83635, w_eco83636, w_eco83637, w_eco83638, w_eco83639, w_eco83640, w_eco83641, w_eco83642, w_eco83643, w_eco83644, w_eco83645, w_eco83646, w_eco83647, w_eco83648, w_eco83649, w_eco83650, w_eco83651, w_eco83652, w_eco83653, w_eco83654, w_eco83655, w_eco83656, w_eco83657, w_eco83658, w_eco83659, w_eco83660, w_eco83661, w_eco83662, w_eco83663, w_eco83664, w_eco83665, w_eco83666, w_eco83667, w_eco83668, w_eco83669, w_eco83670, w_eco83671, w_eco83672, w_eco83673, w_eco83674, w_eco83675, w_eco83676, w_eco83677, w_eco83678, w_eco83679, w_eco83680, w_eco83681, w_eco83682, w_eco83683, w_eco83684, w_eco83685, w_eco83686, w_eco83687, w_eco83688, w_eco83689, w_eco83690, w_eco83691, w_eco83692, w_eco83693, w_eco83694, w_eco83695, w_eco83696, w_eco83697, w_eco83698, w_eco83699, w_eco83700, w_eco83701, w_eco83702, w_eco83703, w_eco83704, w_eco83705, w_eco83706, w_eco83707, w_eco83708, w_eco83709, w_eco83710, w_eco83711, w_eco83712, w_eco83713, w_eco83714, w_eco83715, w_eco83716, w_eco83717, w_eco83718, w_eco83719, w_eco83720, w_eco83721, w_eco83722, w_eco83723, w_eco83724, w_eco83725, w_eco83726, w_eco83727, w_eco83728, w_eco83729, w_eco83730, w_eco83731, w_eco83732, w_eco83733, w_eco83734, w_eco83735, w_eco83736, w_eco83737, w_eco83738, w_eco83739, w_eco83740, w_eco83741, w_eco83742, w_eco83743, w_eco83744, w_eco83745, w_eco83746, w_eco83747, w_eco83748, w_eco83749, w_eco83750, w_eco83751, w_eco83752, w_eco83753, w_eco83754, w_eco83755, w_eco83756, w_eco83757, w_eco83758, w_eco83759, w_eco83760, w_eco83761, w_eco83762, w_eco83763, w_eco83764, w_eco83765, w_eco83766, w_eco83767, w_eco83768, w_eco83769, w_eco83770, w_eco83771, w_eco83772, w_eco83773, w_eco83774, w_eco83775, w_eco83776, w_eco83777, w_eco83778, w_eco83779, w_eco83780, w_eco83781, w_eco83782, w_eco83783, w_eco83784, w_eco83785, w_eco83786, w_eco83787, w_eco83788, w_eco83789, w_eco83790, w_eco83791, w_eco83792, w_eco83793, w_eco83794, w_eco83795, w_eco83796, w_eco83797, w_eco83798, w_eco83799, w_eco83800, w_eco83801, w_eco83802, w_eco83803, w_eco83804, w_eco83805, w_eco83806, w_eco83807, w_eco83808, w_eco83809, w_eco83810, w_eco83811, w_eco83812, w_eco83813, w_eco83814, w_eco83815, w_eco83816, w_eco83817, w_eco83818, w_eco83819, w_eco83820, w_eco83821, w_eco83822, w_eco83823, w_eco83824, w_eco83825, w_eco83826, w_eco83827, w_eco83828, w_eco83829, w_eco83830, w_eco83831, w_eco83832, w_eco83833, w_eco83834, w_eco83835, w_eco83836, w_eco83837, w_eco83838, w_eco83839, w_eco83840, w_eco83841, w_eco83842, w_eco83843, w_eco83844, w_eco83845, w_eco83846, w_eco83847, w_eco83848, w_eco83849, w_eco83850, w_eco83851, w_eco83852, w_eco83853, w_eco83854, w_eco83855, w_eco83856, w_eco83857, w_eco83858, w_eco83859, w_eco83860, w_eco83861, w_eco83862, w_eco83863, w_eco83864, w_eco83865, w_eco83866, w_eco83867, w_eco83868, w_eco83869, w_eco83870, w_eco83871, w_eco83872, w_eco83873, w_eco83874, w_eco83875, w_eco83876, w_eco83877, w_eco83878, w_eco83879, w_eco83880, w_eco83881, w_eco83882, w_eco83883, w_eco83884, w_eco83885, w_eco83886, w_eco83887, w_eco83888, w_eco83889, w_eco83890, w_eco83891, w_eco83892, w_eco83893, w_eco83894, w_eco83895, w_eco83896, w_eco83897, w_eco83898, w_eco83899, w_eco83900, w_eco83901, w_eco83902, w_eco83903, w_eco83904, w_eco83905, w_eco83906, w_eco83907, w_eco83908, w_eco83909, w_eco83910, w_eco83911, w_eco83912, w_eco83913, w_eco83914, w_eco83915, w_eco83916, w_eco83917, w_eco83918, w_eco83919, w_eco83920, w_eco83921, w_eco83922, w_eco83923, w_eco83924, w_eco83925, w_eco83926, w_eco83927, w_eco83928, w_eco83929, w_eco83930, w_eco83931, w_eco83932, w_eco83933, w_eco83934, w_eco83935, w_eco83936, w_eco83937, w_eco83938, w_eco83939, w_eco83940, w_eco83941, w_eco83942, w_eco83943, w_eco83944, w_eco83945, w_eco83946, w_eco83947, w_eco83948, w_eco83949, w_eco83950, w_eco83951, w_eco83952, w_eco83953, w_eco83954, w_eco83955, w_eco83956, w_eco83957, w_eco83958, w_eco83959, w_eco83960, w_eco83961, w_eco83962, w_eco83963, w_eco83964, w_eco83965, w_eco83966, w_eco83967, w_eco83968, w_eco83969, w_eco83970, w_eco83971, w_eco83972, w_eco83973, w_eco83974, w_eco83975, w_eco83976, w_eco83977, w_eco83978, w_eco83979, w_eco83980, w_eco83981, w_eco83982, w_eco83983, w_eco83984, w_eco83985, w_eco83986, w_eco83987, w_eco83988, w_eco83989, w_eco83990, w_eco83991, w_eco83992, w_eco83993, w_eco83994, w_eco83995, w_eco83996, w_eco83997, w_eco83998, w_eco83999, w_eco84000, w_eco84001, w_eco84002, w_eco84003, w_eco84004, w_eco84005, w_eco84006, w_eco84007, w_eco84008, w_eco84009, w_eco84010, w_eco84011, w_eco84012, w_eco84013, w_eco84014, w_eco84015, w_eco84016, w_eco84017, w_eco84018, w_eco84019, w_eco84020, w_eco84021, w_eco84022, w_eco84023, w_eco84024, w_eco84025, w_eco84026, w_eco84027, w_eco84028, w_eco84029, w_eco84030, w_eco84031, w_eco84032, w_eco84033, w_eco84034, w_eco84035, w_eco84036, w_eco84037, w_eco84038, w_eco84039, w_eco84040, w_eco84041, w_eco84042, w_eco84043, w_eco84044, w_eco84045, w_eco84046, w_eco84047, w_eco84048, w_eco84049, w_eco84050, w_eco84051, w_eco84052, w_eco84053, w_eco84054, w_eco84055, w_eco84056, w_eco84057, w_eco84058, w_eco84059, w_eco84060, w_eco84061, w_eco84062, w_eco84063, w_eco84064, w_eco84065, w_eco84066, w_eco84067, w_eco84068, w_eco84069, w_eco84070, w_eco84071, w_eco84072, w_eco84073, w_eco84074, w_eco84075, w_eco84076, w_eco84077, w_eco84078, w_eco84079, w_eco84080, w_eco84081, w_eco84082, w_eco84083, w_eco84084, w_eco84085, w_eco84086, w_eco84087, w_eco84088, w_eco84089, w_eco84090, w_eco84091, w_eco84092, w_eco84093, w_eco84094, w_eco84095, w_eco84096, w_eco84097, w_eco84098, w_eco84099, w_eco84100, w_eco84101, w_eco84102, w_eco84103, w_eco84104, w_eco84105, w_eco84106, w_eco84107, w_eco84108, w_eco84109, w_eco84110, w_eco84111, w_eco84112, w_eco84113, w_eco84114, w_eco84115, w_eco84116, w_eco84117, w_eco84118, w_eco84119, w_eco84120, w_eco84121, w_eco84122, w_eco84123, w_eco84124, w_eco84125, w_eco84126, w_eco84127, w_eco84128, w_eco84129, w_eco84130, w_eco84131, w_eco84132, w_eco84133, w_eco84134, w_eco84135, w_eco84136, w_eco84137, w_eco84138, w_eco84139, w_eco84140, w_eco84141, w_eco84142, w_eco84143, w_eco84144, w_eco84145, w_eco84146, w_eco84147, w_eco84148, w_eco84149, w_eco84150, w_eco84151, w_eco84152, w_eco84153, w_eco84154, w_eco84155, w_eco84156, w_eco84157, w_eco84158, w_eco84159, w_eco84160, w_eco84161, w_eco84162, w_eco84163, w_eco84164, w_eco84165, w_eco84166, w_eco84167, w_eco84168, w_eco84169, w_eco84170, w_eco84171, w_eco84172, w_eco84173, w_eco84174, w_eco84175, w_eco84176, w_eco84177, w_eco84178, w_eco84179, w_eco84180, w_eco84181, w_eco84182, w_eco84183, w_eco84184, w_eco84185, w_eco84186, w_eco84187, w_eco84188, w_eco84189, w_eco84190, w_eco84191, w_eco84192, w_eco84193, w_eco84194, w_eco84195, w_eco84196, w_eco84197, w_eco84198, w_eco84199, w_eco84200, w_eco84201, w_eco84202, w_eco84203, w_eco84204, w_eco84205, w_eco84206, w_eco84207, w_eco84208, w_eco84209, w_eco84210, w_eco84211, w_eco84212, w_eco84213, w_eco84214, w_eco84215, w_eco84216, w_eco84217, w_eco84218, w_eco84219, w_eco84220, w_eco84221, w_eco84222, w_eco84223, w_eco84224, w_eco84225, w_eco84226, w_eco84227, w_eco84228, w_eco84229, w_eco84230, w_eco84231, w_eco84232, w_eco84233, w_eco84234, w_eco84235, w_eco84236, w_eco84237, w_eco84238, w_eco84239, w_eco84240, w_eco84241, w_eco84242, w_eco84243, w_eco84244, w_eco84245, w_eco84246, w_eco84247, w_eco84248, w_eco84249, w_eco84250, w_eco84251, w_eco84252, w_eco84253, w_eco84254, w_eco84255, w_eco84256, w_eco84257, w_eco84258, w_eco84259, w_eco84260, w_eco84261, w_eco84262, w_eco84263, w_eco84264, w_eco84265, w_eco84266, w_eco84267, w_eco84268, w_eco84269, w_eco84270, w_eco84271, w_eco84272, w_eco84273, w_eco84274, w_eco84275, w_eco84276, w_eco84277, w_eco84278, w_eco84279, w_eco84280, w_eco84281, w_eco84282, w_eco84283, w_eco84284, w_eco84285, w_eco84286, w_eco84287, w_eco84288, w_eco84289, w_eco84290, w_eco84291, w_eco84292, w_eco84293, w_eco84294, w_eco84295, w_eco84296, w_eco84297, w_eco84298, w_eco84299, w_eco84300, w_eco84301, w_eco84302, w_eco84303, w_eco84304, w_eco84305, w_eco84306, w_eco84307, w_eco84308, w_eco84309, w_eco84310, w_eco84311, w_eco84312, w_eco84313, w_eco84314, w_eco84315, w_eco84316, w_eco84317, w_eco84318, w_eco84319, w_eco84320, w_eco84321, w_eco84322, w_eco84323, w_eco84324, w_eco84325, w_eco84326, w_eco84327, w_eco84328, w_eco84329, w_eco84330, w_eco84331, w_eco84332, w_eco84333, w_eco84334, w_eco84335, w_eco84336, w_eco84337, w_eco84338, w_eco84339, w_eco84340, w_eco84341, w_eco84342, w_eco84343, w_eco84344, w_eco84345, w_eco84346, w_eco84347, w_eco84348, w_eco84349, w_eco84350, w_eco84351, w_eco84352, w_eco84353, w_eco84354, w_eco84355, w_eco84356, w_eco84357, w_eco84358, w_eco84359, w_eco84360, w_eco84361, w_eco84362, w_eco84363, w_eco84364, w_eco84365, w_eco84366, w_eco84367, w_eco84368, w_eco84369, w_eco84370, w_eco84371, w_eco84372, w_eco84373, w_eco84374, w_eco84375, w_eco84376, w_eco84377, w_eco84378, w_eco84379, w_eco84380, w_eco84381, w_eco84382, w_eco84383, w_eco84384, w_eco84385, w_eco84386, w_eco84387, w_eco84388, w_eco84389, w_eco84390, w_eco84391, w_eco84392, w_eco84393, w_eco84394, w_eco84395, w_eco84396, w_eco84397, w_eco84398, w_eco84399, w_eco84400, w_eco84401, w_eco84402, w_eco84403, w_eco84404, w_eco84405, w_eco84406, w_eco84407, w_eco84408, w_eco84409, w_eco84410, w_eco84411, w_eco84412, w_eco84413, w_eco84414, w_eco84415, w_eco84416, w_eco84417, w_eco84418, w_eco84419, w_eco84420, w_eco84421, w_eco84422, w_eco84423, w_eco84424, w_eco84425, w_eco84426, w_eco84427, w_eco84428, w_eco84429, w_eco84430, w_eco84431, w_eco84432, w_eco84433, w_eco84434, w_eco84435, w_eco84436, w_eco84437, w_eco84438, w_eco84439, w_eco84440, w_eco84441, w_eco84442, w_eco84443, w_eco84444, w_eco84445, w_eco84446, w_eco84447, w_eco84448, w_eco84449, w_eco84450, w_eco84451, w_eco84452, w_eco84453, w_eco84454, w_eco84455, w_eco84456, w_eco84457, w_eco84458, w_eco84459, w_eco84460, w_eco84461, w_eco84462, w_eco84463, w_eco84464, w_eco84465, w_eco84466, w_eco84467, w_eco84468, w_eco84469, w_eco84470, w_eco84471, w_eco84472, w_eco84473, w_eco84474, w_eco84475, w_eco84476, w_eco84477, w_eco84478, w_eco84479, w_eco84480, w_eco84481, w_eco84482, w_eco84483, w_eco84484, w_eco84485, w_eco84486, w_eco84487, w_eco84488, w_eco84489, w_eco84490, w_eco84491, w_eco84492, w_eco84493, w_eco84494, w_eco84495, w_eco84496, w_eco84497, w_eco84498, w_eco84499, w_eco84500, w_eco84501, w_eco84502, w_eco84503, w_eco84504, w_eco84505, w_eco84506, w_eco84507, w_eco84508, w_eco84509, w_eco84510, w_eco84511, w_eco84512, w_eco84513, w_eco84514, w_eco84515, w_eco84516, w_eco84517, w_eco84518, w_eco84519, w_eco84520, w_eco84521, w_eco84522, w_eco84523, w_eco84524, w_eco84525, w_eco84526, w_eco84527, w_eco84528, w_eco84529, w_eco84530, w_eco84531, w_eco84532, w_eco84533, w_eco84534, w_eco84535, w_eco84536, w_eco84537, w_eco84538, w_eco84539, w_eco84540, w_eco84541, w_eco84542, w_eco84543, w_eco84544, w_eco84545, w_eco84546, w_eco84547, w_eco84548, w_eco84549, w_eco84550, w_eco84551, w_eco84552, w_eco84553, w_eco84554, w_eco84555, w_eco84556, w_eco84557, w_eco84558, w_eco84559, w_eco84560, w_eco84561, w_eco84562, w_eco84563, w_eco84564, w_eco84565, w_eco84566, w_eco84567, w_eco84568, w_eco84569, w_eco84570, w_eco84571, w_eco84572, w_eco84573, w_eco84574, w_eco84575, w_eco84576, w_eco84577, w_eco84578, w_eco84579, w_eco84580, w_eco84581, w_eco84582, w_eco84583, w_eco84584, w_eco84585, w_eco84586, w_eco84587, w_eco84588, w_eco84589, w_eco84590, w_eco84591, w_eco84592, w_eco84593, w_eco84594, w_eco84595, w_eco84596, w_eco84597, w_eco84598, w_eco84599, w_eco84600, w_eco84601, w_eco84602, w_eco84603, w_eco84604, w_eco84605, w_eco84606, w_eco84607, w_eco84608, w_eco84609, w_eco84610, w_eco84611, w_eco84612, w_eco84613, w_eco84614, w_eco84615, w_eco84616, w_eco84617, w_eco84618, w_eco84619, w_eco84620, w_eco84621, w_eco84622, w_eco84623, w_eco84624, w_eco84625, w_eco84626, w_eco84627, w_eco84628, w_eco84629, w_eco84630, w_eco84631, w_eco84632, w_eco84633, w_eco84634, w_eco84635, w_eco84636, w_eco84637, w_eco84638, w_eco84639, w_eco84640, w_eco84641, w_eco84642, w_eco84643, w_eco84644, w_eco84645, w_eco84646, w_eco84647, w_eco84648, w_eco84649, w_eco84650, w_eco84651, w_eco84652, w_eco84653, w_eco84654, w_eco84655, w_eco84656, w_eco84657, w_eco84658, w_eco84659, w_eco84660, w_eco84661, w_eco84662, w_eco84663, w_eco84664, w_eco84665, w_eco84666, w_eco84667, w_eco84668, w_eco84669, w_eco84670, w_eco84671, w_eco84672, w_eco84673, w_eco84674, w_eco84675, w_eco84676, w_eco84677, w_eco84678, w_eco84679, w_eco84680, w_eco84681, w_eco84682, w_eco84683, w_eco84684, w_eco84685, w_eco84686, w_eco84687, w_eco84688, w_eco84689, w_eco84690, w_eco84691, w_eco84692, w_eco84693, w_eco84694, w_eco84695, w_eco84696, w_eco84697, w_eco84698, w_eco84699, w_eco84700, w_eco84701, w_eco84702, w_eco84703, w_eco84704, w_eco84705, w_eco84706, w_eco84707, w_eco84708, w_eco84709, w_eco84710, w_eco84711, w_eco84712, w_eco84713, w_eco84714, w_eco84715, w_eco84716, w_eco84717, w_eco84718, w_eco84719, w_eco84720, w_eco84721, w_eco84722, w_eco84723, w_eco84724, w_eco84725, w_eco84726, w_eco84727, w_eco84728, w_eco84729, w_eco84730, w_eco84731, w_eco84732, w_eco84733, w_eco84734, w_eco84735, w_eco84736, w_eco84737, w_eco84738, w_eco84739, w_eco84740, w_eco84741, w_eco84742, w_eco84743, w_eco84744, w_eco84745, w_eco84746, w_eco84747, w_eco84748, w_eco84749, w_eco84750, w_eco84751, w_eco84752, w_eco84753, w_eco84754, w_eco84755, w_eco84756, w_eco84757, w_eco84758, w_eco84759, w_eco84760, w_eco84761, w_eco84762, w_eco84763, w_eco84764, w_eco84765, w_eco84766, w_eco84767, w_eco84768, w_eco84769, w_eco84770, w_eco84771, w_eco84772, w_eco84773, w_eco84774, w_eco84775, w_eco84776, w_eco84777, w_eco84778, w_eco84779, w_eco84780, w_eco84781, w_eco84782, w_eco84783, w_eco84784, w_eco84785, w_eco84786, w_eco84787, w_eco84788, w_eco84789, w_eco84790, w_eco84791, w_eco84792, w_eco84793, w_eco84794, w_eco84795, w_eco84796, w_eco84797, w_eco84798, w_eco84799, w_eco84800, w_eco84801, w_eco84802, w_eco84803, w_eco84804, w_eco84805, w_eco84806, w_eco84807, w_eco84808, w_eco84809, w_eco84810, w_eco84811, w_eco84812, w_eco84813, w_eco84814, w_eco84815, w_eco84816, w_eco84817, w_eco84818, w_eco84819, w_eco84820, w_eco84821, w_eco84822, w_eco84823, w_eco84824, w_eco84825, w_eco84826, w_eco84827, w_eco84828, w_eco84829, w_eco84830, w_eco84831, w_eco84832, w_eco84833, w_eco84834, w_eco84835, w_eco84836, w_eco84837, w_eco84838, w_eco84839, w_eco84840, w_eco84841, w_eco84842, w_eco84843, w_eco84844, w_eco84845, w_eco84846, w_eco84847, w_eco84848, w_eco84849, w_eco84850, w_eco84851, w_eco84852, w_eco84853, w_eco84854, w_eco84855, w_eco84856, w_eco84857, w_eco84858, w_eco84859, w_eco84860, w_eco84861, w_eco84862, w_eco84863, w_eco84864, w_eco84865, w_eco84866, w_eco84867, w_eco84868, w_eco84869, w_eco84870, w_eco84871, w_eco84872, w_eco84873, w_eco84874, w_eco84875, w_eco84876, w_eco84877, w_eco84878, w_eco84879, w_eco84880, w_eco84881, w_eco84882, w_eco84883, w_eco84884, w_eco84885, w_eco84886, w_eco84887, w_eco84888, w_eco84889, w_eco84890, w_eco84891, w_eco84892, w_eco84893, w_eco84894, w_eco84895, w_eco84896, w_eco84897, w_eco84898, w_eco84899, w_eco84900, w_eco84901, w_eco84902, w_eco84903, w_eco84904, w_eco84905, w_eco84906, w_eco84907, w_eco84908, w_eco84909, w_eco84910, w_eco84911, w_eco84912, w_eco84913, w_eco84914, w_eco84915, w_eco84916, w_eco84917, w_eco84918, w_eco84919, w_eco84920, w_eco84921, w_eco84922, w_eco84923, w_eco84924, w_eco84925, w_eco84926, w_eco84927, w_eco84928, w_eco84929, w_eco84930, w_eco84931, w_eco84932, w_eco84933, w_eco84934, w_eco84935, w_eco84936, w_eco84937, w_eco84938, w_eco84939, w_eco84940, w_eco84941, w_eco84942, w_eco84943, w_eco84944, w_eco84945, w_eco84946, w_eco84947, w_eco84948, w_eco84949, w_eco84950, w_eco84951, w_eco84952, w_eco84953, w_eco84954, w_eco84955, w_eco84956, w_eco84957, w_eco84958, w_eco84959, w_eco84960, w_eco84961, w_eco84962, w_eco84963, w_eco84964, w_eco84965, w_eco84966, w_eco84967, w_eco84968, w_eco84969, w_eco84970, w_eco84971, w_eco84972, w_eco84973, w_eco84974, w_eco84975, w_eco84976, w_eco84977, w_eco84978, w_eco84979, w_eco84980, w_eco84981, w_eco84982, w_eco84983, w_eco84984, w_eco84985, w_eco84986, w_eco84987, w_eco84988, w_eco84989, w_eco84990, w_eco84991, w_eco84992, w_eco84993, w_eco84994, w_eco84995, w_eco84996, w_eco84997, w_eco84998, w_eco84999, w_eco85000, w_eco85001, w_eco85002, w_eco85003, w_eco85004, w_eco85005, w_eco85006, w_eco85007, w_eco85008, w_eco85009, w_eco85010, w_eco85011, w_eco85012, w_eco85013, w_eco85014, w_eco85015, w_eco85016, w_eco85017, w_eco85018, w_eco85019, w_eco85020, w_eco85021, w_eco85022, w_eco85023, w_eco85024, w_eco85025, w_eco85026, w_eco85027, w_eco85028, w_eco85029, w_eco85030, w_eco85031, w_eco85032, w_eco85033, w_eco85034, w_eco85035, w_eco85036, w_eco85037, w_eco85038, w_eco85039, w_eco85040, w_eco85041, w_eco85042, w_eco85043, w_eco85044, w_eco85045, w_eco85046, w_eco85047, w_eco85048, w_eco85049, w_eco85050, w_eco85051, w_eco85052, w_eco85053, w_eco85054, w_eco85055, w_eco85056, w_eco85057, w_eco85058, w_eco85059, w_eco85060, w_eco85061, w_eco85062, w_eco85063, w_eco85064, w_eco85065, w_eco85066, w_eco85067, w_eco85068, w_eco85069, w_eco85070, w_eco85071, w_eco85072, w_eco85073, w_eco85074, w_eco85075, w_eco85076, w_eco85077, w_eco85078, w_eco85079, w_eco85080, w_eco85081, w_eco85082, w_eco85083, w_eco85084, w_eco85085, w_eco85086, w_eco85087, w_eco85088, w_eco85089, w_eco85090, w_eco85091, w_eco85092, w_eco85093, w_eco85094, w_eco85095, w_eco85096, w_eco85097, w_eco85098, w_eco85099, w_eco85100, w_eco85101, w_eco85102, w_eco85103, w_eco85104, w_eco85105, w_eco85106, w_eco85107, w_eco85108, w_eco85109, w_eco85110, w_eco85111, w_eco85112, w_eco85113, w_eco85114, w_eco85115, w_eco85116, w_eco85117, w_eco85118, w_eco85119, w_eco85120, w_eco85121, w_eco85122, w_eco85123, w_eco85124, w_eco85125, w_eco85126, w_eco85127, w_eco85128, w_eco85129, w_eco85130, w_eco85131, w_eco85132, w_eco85133, w_eco85134, w_eco85135, w_eco85136, w_eco85137, w_eco85138, w_eco85139, w_eco85140, w_eco85141, w_eco85142, w_eco85143, w_eco85144, w_eco85145, w_eco85146, w_eco85147, w_eco85148, w_eco85149, w_eco85150, w_eco85151, w_eco85152, w_eco85153, w_eco85154, w_eco85155, w_eco85156, w_eco85157, w_eco85158, w_eco85159, w_eco85160, w_eco85161, w_eco85162, w_eco85163, w_eco85164, w_eco85165, w_eco85166, w_eco85167, w_eco85168, w_eco85169, w_eco85170, w_eco85171, w_eco85172, w_eco85173, w_eco85174, w_eco85175, w_eco85176, w_eco85177, w_eco85178, w_eco85179, w_eco85180, w_eco85181, w_eco85182, w_eco85183, w_eco85184, w_eco85185, w_eco85186, w_eco85187, w_eco85188, w_eco85189, w_eco85190, w_eco85191, w_eco85192, w_eco85193, w_eco85194, w_eco85195, w_eco85196, w_eco85197, w_eco85198, w_eco85199, w_eco85200, w_eco85201, w_eco85202, w_eco85203, w_eco85204, w_eco85205, w_eco85206, w_eco85207, w_eco85208, w_eco85209, w_eco85210, w_eco85211, w_eco85212, w_eco85213, w_eco85214, w_eco85215, w_eco85216, w_eco85217, w_eco85218, w_eco85219, w_eco85220, w_eco85221, w_eco85222, w_eco85223, w_eco85224, w_eco85225, w_eco85226, w_eco85227, w_eco85228, w_eco85229, w_eco85230, w_eco85231, w_eco85232, w_eco85233, w_eco85234, w_eco85235, w_eco85236, w_eco85237, w_eco85238, w_eco85239, w_eco85240, w_eco85241, w_eco85242, w_eco85243, w_eco85244, w_eco85245, w_eco85246, w_eco85247, w_eco85248, w_eco85249, w_eco85250, w_eco85251, w_eco85252, w_eco85253, w_eco85254, w_eco85255, w_eco85256, w_eco85257, w_eco85258, w_eco85259, w_eco85260, w_eco85261, w_eco85262, w_eco85263, w_eco85264, w_eco85265, w_eco85266, w_eco85267, w_eco85268, w_eco85269, w_eco85270, w_eco85271, w_eco85272, w_eco85273, w_eco85274, w_eco85275, w_eco85276, w_eco85277, w_eco85278, w_eco85279, w_eco85280, w_eco85281, w_eco85282, w_eco85283, w_eco85284, w_eco85285, w_eco85286, w_eco85287, w_eco85288, w_eco85289, w_eco85290, w_eco85291, w_eco85292, w_eco85293, w_eco85294, w_eco85295, w_eco85296, w_eco85297, w_eco85298, w_eco85299, w_eco85300, w_eco85301, w_eco85302, w_eco85303, w_eco85304, w_eco85305, w_eco85306, w_eco85307, w_eco85308, w_eco85309, w_eco85310, w_eco85311, w_eco85312, w_eco85313, w_eco85314, w_eco85315, w_eco85316, w_eco85317, w_eco85318, w_eco85319, w_eco85320, w_eco85321, w_eco85322, w_eco85323, w_eco85324, w_eco85325, w_eco85326, w_eco85327, w_eco85328, w_eco85329, w_eco85330, w_eco85331, w_eco85332, w_eco85333, w_eco85334, w_eco85335, w_eco85336, w_eco85337, w_eco85338, w_eco85339, w_eco85340, w_eco85341, w_eco85342, w_eco85343, w_eco85344, w_eco85345, w_eco85346, w_eco85347, w_eco85348, w_eco85349, w_eco85350, w_eco85351, w_eco85352, w_eco85353, w_eco85354, w_eco85355, w_eco85356, w_eco85357, w_eco85358, w_eco85359, w_eco85360, w_eco85361, w_eco85362, w_eco85363, w_eco85364, w_eco85365, w_eco85366, w_eco85367, w_eco85368, w_eco85369, w_eco85370, w_eco85371, w_eco85372, w_eco85373, w_eco85374, w_eco85375, w_eco85376, w_eco85377, w_eco85378, w_eco85379, w_eco85380, w_eco85381, w_eco85382, w_eco85383, w_eco85384, w_eco85385, w_eco85386, w_eco85387, w_eco85388, w_eco85389, w_eco85390, w_eco85391, w_eco85392, w_eco85393, w_eco85394, w_eco85395, w_eco85396, w_eco85397, w_eco85398, w_eco85399, w_eco85400, w_eco85401, w_eco85402, w_eco85403, w_eco85404, w_eco85405, w_eco85406, w_eco85407, w_eco85408, w_eco85409, w_eco85410, w_eco85411, w_eco85412, w_eco85413, w_eco85414, w_eco85415, w_eco85416, w_eco85417, w_eco85418, w_eco85419, w_eco85420, w_eco85421, w_eco85422, w_eco85423, w_eco85424, w_eco85425, w_eco85426, w_eco85427, w_eco85428, w_eco85429, w_eco85430, w_eco85431, w_eco85432, w_eco85433, w_eco85434, w_eco85435, w_eco85436, w_eco85437, w_eco85438, w_eco85439, w_eco85440, w_eco85441, w_eco85442, w_eco85443, w_eco85444, w_eco85445, w_eco85446, w_eco85447, w_eco85448, w_eco85449, w_eco85450, w_eco85451, w_eco85452, w_eco85453, w_eco85454, w_eco85455, w_eco85456, w_eco85457, w_eco85458, w_eco85459, w_eco85460, w_eco85461, w_eco85462, w_eco85463, w_eco85464, w_eco85465, w_eco85466, w_eco85467, w_eco85468, w_eco85469, w_eco85470, w_eco85471, w_eco85472, w_eco85473, w_eco85474, w_eco85475, w_eco85476, w_eco85477, w_eco85478, w_eco85479, w_eco85480, w_eco85481, w_eco85482, w_eco85483, w_eco85484, w_eco85485, w_eco85486, w_eco85487, w_eco85488, w_eco85489, w_eco85490, w_eco85491, w_eco85492, w_eco85493, w_eco85494, w_eco85495, w_eco85496, w_eco85497, w_eco85498, w_eco85499, w_eco85500, w_eco85501, w_eco85502, w_eco85503, w_eco85504, w_eco85505, w_eco85506, w_eco85507, w_eco85508, w_eco85509, w_eco85510, w_eco85511, w_eco85512, w_eco85513, w_eco85514, w_eco85515, w_eco85516, w_eco85517, w_eco85518, w_eco85519, w_eco85520, w_eco85521, w_eco85522, w_eco85523, w_eco85524, w_eco85525, w_eco85526, w_eco85527, w_eco85528, w_eco85529, w_eco85530, w_eco85531, w_eco85532, w_eco85533, w_eco85534, w_eco85535, w_eco85536, w_eco85537, w_eco85538, w_eco85539, w_eco85540, w_eco85541, w_eco85542, w_eco85543, w_eco85544, w_eco85545, w_eco85546, w_eco85547, w_eco85548, w_eco85549, w_eco85550, w_eco85551, w_eco85552, w_eco85553, w_eco85554, w_eco85555, w_eco85556, w_eco85557, w_eco85558, w_eco85559, w_eco85560, w_eco85561, w_eco85562, w_eco85563, w_eco85564, w_eco85565, w_eco85566, w_eco85567, w_eco85568, w_eco85569, w_eco85570, w_eco85571, w_eco85572, w_eco85573, w_eco85574, w_eco85575, w_eco85576, w_eco85577, w_eco85578, w_eco85579, w_eco85580, w_eco85581, w_eco85582, w_eco85583, w_eco85584, w_eco85585, w_eco85586, w_eco85587, w_eco85588, w_eco85589, w_eco85590, w_eco85591, w_eco85592, w_eco85593, w_eco85594, w_eco85595, w_eco85596, w_eco85597, w_eco85598, w_eco85599, w_eco85600, w_eco85601, w_eco85602, w_eco85603, w_eco85604, w_eco85605, w_eco85606, w_eco85607, w_eco85608, w_eco85609, w_eco85610, w_eco85611, w_eco85612, w_eco85613, w_eco85614, w_eco85615, w_eco85616, w_eco85617, w_eco85618, w_eco85619, w_eco85620, w_eco85621, w_eco85622, w_eco85623, w_eco85624, w_eco85625, w_eco85626, w_eco85627, w_eco85628, w_eco85629, w_eco85630, w_eco85631, w_eco85632, w_eco85633, w_eco85634, w_eco85635, w_eco85636, w_eco85637, w_eco85638, w_eco85639, w_eco85640, w_eco85641, w_eco85642, w_eco85643, w_eco85644, w_eco85645, w_eco85646, w_eco85647, w_eco85648, w_eco85649, w_eco85650, w_eco85651, w_eco85652, w_eco85653, w_eco85654, w_eco85655, w_eco85656, w_eco85657, w_eco85658, w_eco85659, w_eco85660, w_eco85661, w_eco85662, w_eco85663, w_eco85664, w_eco85665, w_eco85666, w_eco85667, w_eco85668, w_eco85669, w_eco85670, w_eco85671, w_eco85672, w_eco85673, w_eco85674, w_eco85675, w_eco85676, w_eco85677, w_eco85678, w_eco85679, w_eco85680, w_eco85681, w_eco85682, w_eco85683, w_eco85684, w_eco85685, w_eco85686, w_eco85687, w_eco85688, w_eco85689, w_eco85690, w_eco85691, w_eco85692, w_eco85693, w_eco85694, w_eco85695, w_eco85696, w_eco85697, w_eco85698, w_eco85699, w_eco85700, w_eco85701, w_eco85702, w_eco85703, w_eco85704, w_eco85705, w_eco85706, w_eco85707, w_eco85708, w_eco85709, w_eco85710, w_eco85711, w_eco85712, w_eco85713, w_eco85714, w_eco85715, w_eco85716, w_eco85717, w_eco85718, w_eco85719, w_eco85720, w_eco85721, w_eco85722, w_eco85723, w_eco85724, w_eco85725, w_eco85726, w_eco85727, w_eco85728, w_eco85729, w_eco85730, w_eco85731, w_eco85732, w_eco85733, w_eco85734, w_eco85735, w_eco85736, w_eco85737, w_eco85738, w_eco85739, w_eco85740, w_eco85741, w_eco85742, w_eco85743, w_eco85744, w_eco85745, w_eco85746, w_eco85747, w_eco85748, w_eco85749, w_eco85750, w_eco85751, w_eco85752, w_eco85753, w_eco85754, w_eco85755, w_eco85756, w_eco85757, w_eco85758, w_eco85759, w_eco85760, w_eco85761, w_eco85762, w_eco85763, w_eco85764, w_eco85765, w_eco85766, w_eco85767, w_eco85768, w_eco85769, w_eco85770, w_eco85771, w_eco85772, w_eco85773, w_eco85774, w_eco85775, w_eco85776, w_eco85777, w_eco85778, w_eco85779, w_eco85780, w_eco85781, w_eco85782, w_eco85783, w_eco85784, w_eco85785, w_eco85786, w_eco85787, w_eco85788, w_eco85789, w_eco85790, w_eco85791, w_eco85792, w_eco85793, w_eco85794, w_eco85795, w_eco85796, w_eco85797, w_eco85798, w_eco85799, w_eco85800, w_eco85801, w_eco85802, w_eco85803, w_eco85804, w_eco85805, w_eco85806, w_eco85807, w_eco85808, w_eco85809, w_eco85810, w_eco85811, w_eco85812, w_eco85813, w_eco85814, w_eco85815, w_eco85816, w_eco85817, w_eco85818, w_eco85819, w_eco85820, w_eco85821, w_eco85822, w_eco85823, w_eco85824, w_eco85825, w_eco85826, w_eco85827, w_eco85828, w_eco85829, w_eco85830, w_eco85831, w_eco85832, w_eco85833, w_eco85834, w_eco85835, w_eco85836, w_eco85837, w_eco85838, w_eco85839, w_eco85840, w_eco85841, w_eco85842, w_eco85843, w_eco85844, w_eco85845, w_eco85846, w_eco85847, w_eco85848, w_eco85849, w_eco85850, w_eco85851, w_eco85852, w_eco85853, w_eco85854, w_eco85855, w_eco85856, w_eco85857, w_eco85858, w_eco85859, w_eco85860, w_eco85861, w_eco85862, w_eco85863, w_eco85864, w_eco85865, w_eco85866, w_eco85867, w_eco85868, w_eco85869, w_eco85870, w_eco85871, w_eco85872, w_eco85873, w_eco85874, w_eco85875, w_eco85876, w_eco85877, w_eco85878, w_eco85879, w_eco85880, w_eco85881, w_eco85882, w_eco85883, w_eco85884, w_eco85885, w_eco85886, w_eco85887, w_eco85888, w_eco85889, w_eco85890, w_eco85891, w_eco85892, w_eco85893, w_eco85894, w_eco85895, w_eco85896, w_eco85897, w_eco85898, w_eco85899, w_eco85900, w_eco85901, w_eco85902, w_eco85903, w_eco85904, w_eco85905, w_eco85906, w_eco85907, w_eco85908, w_eco85909, w_eco85910, w_eco85911, w_eco85912, w_eco85913, w_eco85914, w_eco85915, w_eco85916, w_eco85917, w_eco85918, w_eco85919, w_eco85920, w_eco85921, w_eco85922, w_eco85923, w_eco85924, w_eco85925, w_eco85926, w_eco85927, w_eco85928, w_eco85929, w_eco85930, w_eco85931, w_eco85932, w_eco85933, w_eco85934, w_eco85935, w_eco85936, w_eco85937, w_eco85938, w_eco85939, w_eco85940, w_eco85941, w_eco85942, w_eco85943, w_eco85944, w_eco85945, w_eco85946, w_eco85947, w_eco85948, w_eco85949, w_eco85950, w_eco85951, w_eco85952, w_eco85953, w_eco85954, w_eco85955, w_eco85956, w_eco85957, w_eco85958, w_eco85959, w_eco85960, w_eco85961, w_eco85962, w_eco85963, w_eco85964, w_eco85965, w_eco85966, w_eco85967, w_eco85968, w_eco85969, w_eco85970, w_eco85971, w_eco85972, w_eco85973, w_eco85974, w_eco85975, w_eco85976, w_eco85977, w_eco85978, w_eco85979, w_eco85980, w_eco85981, w_eco85982, w_eco85983, w_eco85984, w_eco85985, w_eco85986, w_eco85987, w_eco85988, w_eco85989, w_eco85990, w_eco85991, w_eco85992, w_eco85993, w_eco85994, w_eco85995, w_eco85996, w_eco85997, w_eco85998, w_eco85999, w_eco86000, w_eco86001, w_eco86002, w_eco86003, w_eco86004, w_eco86005, w_eco86006, w_eco86007, w_eco86008, w_eco86009, w_eco86010, w_eco86011, w_eco86012, w_eco86013, w_eco86014, w_eco86015, w_eco86016, w_eco86017, w_eco86018, w_eco86019, w_eco86020, w_eco86021, w_eco86022, w_eco86023, w_eco86024, w_eco86025, w_eco86026, w_eco86027, w_eco86028, w_eco86029, w_eco86030, w_eco86031, w_eco86032, w_eco86033, w_eco86034, w_eco86035, w_eco86036, w_eco86037, w_eco86038, w_eco86039, w_eco86040, w_eco86041, w_eco86042, w_eco86043, w_eco86044, w_eco86045, w_eco86046, w_eco86047, w_eco86048, w_eco86049, w_eco86050, w_eco86051, w_eco86052, w_eco86053, w_eco86054, w_eco86055, w_eco86056, w_eco86057, w_eco86058, w_eco86059, w_eco86060, w_eco86061, w_eco86062, w_eco86063, w_eco86064, w_eco86065, w_eco86066, w_eco86067, w_eco86068, w_eco86069, w_eco86070, w_eco86071, w_eco86072, w_eco86073, w_eco86074, w_eco86075, w_eco86076, w_eco86077, w_eco86078, w_eco86079, w_eco86080, w_eco86081, w_eco86082, w_eco86083, w_eco86084, w_eco86085, w_eco86086, w_eco86087, w_eco86088, w_eco86089, w_eco86090, w_eco86091, w_eco86092, w_eco86093, w_eco86094, w_eco86095, w_eco86096, w_eco86097, w_eco86098, w_eco86099, w_eco86100, w_eco86101, w_eco86102, w_eco86103, w_eco86104, w_eco86105, w_eco86106, w_eco86107, w_eco86108, w_eco86109, w_eco86110, w_eco86111, w_eco86112, w_eco86113, w_eco86114, w_eco86115, w_eco86116, w_eco86117, w_eco86118, w_eco86119, w_eco86120, w_eco86121, w_eco86122, w_eco86123, w_eco86124, w_eco86125, w_eco86126, w_eco86127, w_eco86128, w_eco86129, w_eco86130, w_eco86131, w_eco86132, w_eco86133, w_eco86134, w_eco86135, w_eco86136, w_eco86137, w_eco86138, w_eco86139, w_eco86140, w_eco86141, w_eco86142, w_eco86143, w_eco86144, w_eco86145, w_eco86146, w_eco86147, w_eco86148, w_eco86149, w_eco86150, w_eco86151, w_eco86152, w_eco86153, w_eco86154, w_eco86155, w_eco86156, w_eco86157, w_eco86158, w_eco86159, w_eco86160, w_eco86161, w_eco86162, w_eco86163, w_eco86164, w_eco86165, w_eco86166, w_eco86167, w_eco86168, w_eco86169, w_eco86170, w_eco86171, w_eco86172, w_eco86173, w_eco86174, w_eco86175, w_eco86176, w_eco86177, w_eco86178, w_eco86179, w_eco86180, w_eco86181, w_eco86182, w_eco86183, w_eco86184, w_eco86185, w_eco86186, w_eco86187, w_eco86188, w_eco86189, w_eco86190, w_eco86191, w_eco86192, w_eco86193, w_eco86194, w_eco86195, w_eco86196, w_eco86197, w_eco86198, w_eco86199, w_eco86200, w_eco86201, w_eco86202, w_eco86203, w_eco86204, w_eco86205, w_eco86206, w_eco86207, w_eco86208, w_eco86209, w_eco86210, w_eco86211, w_eco86212, w_eco86213, w_eco86214, w_eco86215, w_eco86216, w_eco86217, w_eco86218, w_eco86219, w_eco86220, w_eco86221, w_eco86222, w_eco86223, w_eco86224, w_eco86225, w_eco86226, w_eco86227, w_eco86228, w_eco86229, w_eco86230, w_eco86231, w_eco86232, w_eco86233, w_eco86234, w_eco86235, w_eco86236, w_eco86237, w_eco86238, w_eco86239, w_eco86240, w_eco86241, w_eco86242, w_eco86243, w_eco86244, w_eco86245, w_eco86246, w_eco86247, w_eco86248, w_eco86249, w_eco86250, w_eco86251, w_eco86252, w_eco86253, w_eco86254, w_eco86255, w_eco86256, w_eco86257, w_eco86258, w_eco86259, w_eco86260, w_eco86261, w_eco86262, w_eco86263, w_eco86264, w_eco86265, w_eco86266, w_eco86267, w_eco86268, w_eco86269, w_eco86270, w_eco86271, w_eco86272, w_eco86273, w_eco86274, w_eco86275, w_eco86276, w_eco86277, w_eco86278, w_eco86279, w_eco86280, w_eco86281, w_eco86282, w_eco86283, w_eco86284, w_eco86285, w_eco86286, w_eco86287, w_eco86288, w_eco86289, w_eco86290, w_eco86291, w_eco86292, w_eco86293, w_eco86294, w_eco86295, w_eco86296, w_eco86297, w_eco86298, w_eco86299, w_eco86300, w_eco86301, w_eco86302, w_eco86303, w_eco86304, w_eco86305, w_eco86306, w_eco86307, w_eco86308, w_eco86309, w_eco86310, w_eco86311, w_eco86312, w_eco86313, w_eco86314, w_eco86315, w_eco86316, w_eco86317, w_eco86318, w_eco86319, w_eco86320, w_eco86321, w_eco86322, w_eco86323, w_eco86324, w_eco86325, w_eco86326, w_eco86327, w_eco86328, w_eco86329, w_eco86330, w_eco86331, w_eco86332, w_eco86333, w_eco86334, w_eco86335, w_eco86336, w_eco86337, w_eco86338, w_eco86339, w_eco86340, w_eco86341, w_eco86342, w_eco86343, w_eco86344, w_eco86345, w_eco86346, w_eco86347, w_eco86348, w_eco86349, w_eco86350, w_eco86351, w_eco86352, w_eco86353, w_eco86354, w_eco86355, w_eco86356, w_eco86357, w_eco86358, w_eco86359, w_eco86360, w_eco86361, w_eco86362, w_eco86363, w_eco86364, w_eco86365, w_eco86366, w_eco86367, w_eco86368, w_eco86369, w_eco86370, w_eco86371, w_eco86372, w_eco86373, w_eco86374, w_eco86375, w_eco86376, w_eco86377, w_eco86378, w_eco86379, w_eco86380, w_eco86381, w_eco86382, w_eco86383, w_eco86384, w_eco86385, w_eco86386, w_eco86387, w_eco86388, w_eco86389, w_eco86390, w_eco86391, w_eco86392, w_eco86393, w_eco86394, w_eco86395, w_eco86396, w_eco86397, w_eco86398, w_eco86399, w_eco86400, w_eco86401, w_eco86402, w_eco86403, w_eco86404, w_eco86405, w_eco86406, w_eco86407, w_eco86408, w_eco86409, w_eco86410, w_eco86411, w_eco86412, w_eco86413, w_eco86414, w_eco86415, w_eco86416, w_eco86417, w_eco86418, w_eco86419, w_eco86420, w_eco86421, w_eco86422, w_eco86423, w_eco86424, w_eco86425, w_eco86426, w_eco86427, w_eco86428, w_eco86429, w_eco86430, w_eco86431, w_eco86432, w_eco86433, w_eco86434, w_eco86435, w_eco86436, w_eco86437, w_eco86438, w_eco86439, w_eco86440, w_eco86441, w_eco86442, w_eco86443, w_eco86444, w_eco86445, w_eco86446, w_eco86447, w_eco86448, w_eco86449, w_eco86450, w_eco86451, w_eco86452, w_eco86453, w_eco86454, w_eco86455, w_eco86456, w_eco86457, w_eco86458, w_eco86459, w_eco86460, w_eco86461, w_eco86462, w_eco86463, w_eco86464, w_eco86465, w_eco86466, w_eco86467, w_eco86468, w_eco86469, w_eco86470, w_eco86471, w_eco86472, w_eco86473, w_eco86474, w_eco86475, w_eco86476, w_eco86477, w_eco86478, w_eco86479, w_eco86480, w_eco86481, w_eco86482, w_eco86483, w_eco86484, w_eco86485, w_eco86486, w_eco86487, w_eco86488, w_eco86489, w_eco86490, w_eco86491, w_eco86492, w_eco86493, w_eco86494, w_eco86495, w_eco86496, w_eco86497, w_eco86498, w_eco86499, w_eco86500, w_eco86501, w_eco86502, w_eco86503, w_eco86504, w_eco86505, w_eco86506, w_eco86507, w_eco86508, w_eco86509, w_eco86510, w_eco86511, w_eco86512, w_eco86513, w_eco86514, w_eco86515, w_eco86516, w_eco86517, w_eco86518, w_eco86519, w_eco86520, w_eco86521, w_eco86522, w_eco86523, w_eco86524, w_eco86525, w_eco86526, w_eco86527, w_eco86528, w_eco86529, w_eco86530, w_eco86531, w_eco86532, w_eco86533, w_eco86534, w_eco86535, w_eco86536, w_eco86537, w_eco86538, w_eco86539, w_eco86540, w_eco86541, w_eco86542, w_eco86543, w_eco86544, w_eco86545, w_eco86546, w_eco86547, w_eco86548, w_eco86549, w_eco86550, w_eco86551, w_eco86552, w_eco86553, w_eco86554, w_eco86555, w_eco86556, w_eco86557, w_eco86558, w_eco86559, w_eco86560, w_eco86561, w_eco86562, w_eco86563, w_eco86564, w_eco86565, w_eco86566, w_eco86567, w_eco86568, w_eco86569, w_eco86570, w_eco86571, w_eco86572, w_eco86573, w_eco86574, w_eco86575, w_eco86576, w_eco86577, w_eco86578, w_eco86579, w_eco86580, w_eco86581, w_eco86582, w_eco86583, w_eco86584, w_eco86585, w_eco86586, w_eco86587, w_eco86588, w_eco86589, w_eco86590, w_eco86591, w_eco86592, w_eco86593, w_eco86594, w_eco86595, w_eco86596, w_eco86597, w_eco86598, w_eco86599, w_eco86600, w_eco86601, w_eco86602, w_eco86603, w_eco86604, w_eco86605, w_eco86606, w_eco86607, w_eco86608, w_eco86609, w_eco86610, w_eco86611, w_eco86612, w_eco86613, w_eco86614, w_eco86615, w_eco86616, w_eco86617, w_eco86618, w_eco86619, w_eco86620, w_eco86621, w_eco86622, w_eco86623, w_eco86624, w_eco86625, w_eco86626, w_eco86627, w_eco86628, w_eco86629, w_eco86630, w_eco86631, w_eco86632, w_eco86633, w_eco86634, w_eco86635, w_eco86636, w_eco86637, w_eco86638, w_eco86639, w_eco86640, w_eco86641, w_eco86642, w_eco86643, w_eco86644, w_eco86645, w_eco86646, w_eco86647, w_eco86648, w_eco86649, w_eco86650, w_eco86651, w_eco86652, w_eco86653, w_eco86654, w_eco86655, w_eco86656, w_eco86657, w_eco86658, w_eco86659, w_eco86660, w_eco86661, w_eco86662, w_eco86663, w_eco86664, w_eco86665, w_eco86666, w_eco86667, w_eco86668, w_eco86669, w_eco86670, w_eco86671, w_eco86672, w_eco86673, w_eco86674, w_eco86675, w_eco86676, w_eco86677, w_eco86678, w_eco86679, w_eco86680, w_eco86681, w_eco86682, w_eco86683, w_eco86684, w_eco86685, w_eco86686, w_eco86687, w_eco86688, w_eco86689, w_eco86690, w_eco86691, w_eco86692, w_eco86693, w_eco86694, w_eco86695, w_eco86696, w_eco86697, w_eco86698, w_eco86699, w_eco86700, w_eco86701, w_eco86702, w_eco86703, w_eco86704, w_eco86705, w_eco86706, w_eco86707, w_eco86708, w_eco86709, w_eco86710, w_eco86711, w_eco86712, w_eco86713, w_eco86714, w_eco86715, w_eco86716, w_eco86717, w_eco86718, w_eco86719, w_eco86720, w_eco86721, w_eco86722, w_eco86723, w_eco86724, w_eco86725, w_eco86726, w_eco86727, w_eco86728, w_eco86729, w_eco86730, w_eco86731, w_eco86732, w_eco86733, w_eco86734, w_eco86735, w_eco86736, w_eco86737, w_eco86738, w_eco86739, w_eco86740, w_eco86741, w_eco86742, w_eco86743, w_eco86744, w_eco86745, w_eco86746, w_eco86747, w_eco86748, w_eco86749, w_eco86750, w_eco86751, w_eco86752, w_eco86753, w_eco86754, w_eco86755, w_eco86756, w_eco86757, w_eco86758, w_eco86759, w_eco86760, w_eco86761, w_eco86762, w_eco86763, w_eco86764, w_eco86765, w_eco86766, w_eco86767, w_eco86768, w_eco86769, w_eco86770, w_eco86771, w_eco86772, w_eco86773, w_eco86774, w_eco86775, w_eco86776, w_eco86777, w_eco86778, w_eco86779, w_eco86780, w_eco86781, w_eco86782, w_eco86783, w_eco86784, w_eco86785, w_eco86786, w_eco86787, w_eco86788, w_eco86789, w_eco86790, w_eco86791, w_eco86792, w_eco86793, w_eco86794, w_eco86795, w_eco86796, w_eco86797, w_eco86798, w_eco86799, w_eco86800, w_eco86801, w_eco86802, w_eco86803, w_eco86804, w_eco86805, w_eco86806, w_eco86807, w_eco86808, w_eco86809, w_eco86810, w_eco86811, w_eco86812, w_eco86813, w_eco86814, w_eco86815, w_eco86816, w_eco86817, w_eco86818, w_eco86819, w_eco86820, w_eco86821, w_eco86822, w_eco86823, w_eco86824, w_eco86825, w_eco86826, w_eco86827, w_eco86828, w_eco86829, w_eco86830, w_eco86831, w_eco86832, w_eco86833, w_eco86834, w_eco86835, w_eco86836, w_eco86837, w_eco86838, w_eco86839, w_eco86840, w_eco86841, w_eco86842, w_eco86843, w_eco86844, w_eco86845, w_eco86846, w_eco86847, w_eco86848, w_eco86849, w_eco86850, w_eco86851, w_eco86852, w_eco86853, w_eco86854, w_eco86855, w_eco86856, w_eco86857, w_eco86858, w_eco86859, w_eco86860, w_eco86861, w_eco86862, w_eco86863, w_eco86864, w_eco86865, w_eco86866, w_eco86867, w_eco86868, w_eco86869, w_eco86870, w_eco86871, w_eco86872, w_eco86873, w_eco86874, w_eco86875, w_eco86876, w_eco86877, w_eco86878, w_eco86879, w_eco86880, w_eco86881, w_eco86882, w_eco86883, w_eco86884, w_eco86885, w_eco86886, w_eco86887, w_eco86888, w_eco86889, w_eco86890, w_eco86891, w_eco86892, w_eco86893, w_eco86894, w_eco86895, w_eco86896, w_eco86897, w_eco86898, w_eco86899, w_eco86900, w_eco86901, w_eco86902, w_eco86903, w_eco86904, w_eco86905, w_eco86906, w_eco86907, w_eco86908, w_eco86909, w_eco86910, w_eco86911, w_eco86912, w_eco86913, w_eco86914, w_eco86915, w_eco86916, w_eco86917, w_eco86918, w_eco86919, w_eco86920, w_eco86921, w_eco86922, w_eco86923, w_eco86924, w_eco86925, w_eco86926, w_eco86927, w_eco86928, w_eco86929, w_eco86930, w_eco86931, w_eco86932, w_eco86933, w_eco86934, w_eco86935, w_eco86936, w_eco86937, w_eco86938, w_eco86939, w_eco86940, w_eco86941, w_eco86942, w_eco86943, w_eco86944, w_eco86945, w_eco86946, w_eco86947, w_eco86948, w_eco86949, w_eco86950, w_eco86951, w_eco86952, w_eco86953, w_eco86954, w_eco86955, w_eco86956, w_eco86957, w_eco86958, w_eco86959, w_eco86960, w_eco86961, w_eco86962, w_eco86963, w_eco86964, w_eco86965, w_eco86966, w_eco86967, w_eco86968, w_eco86969, w_eco86970, w_eco86971, w_eco86972, w_eco86973, w_eco86974, w_eco86975, w_eco86976, w_eco86977, w_eco86978, w_eco86979, w_eco86980, w_eco86981, w_eco86982, w_eco86983, w_eco86984, w_eco86985, w_eco86986, w_eco86987, w_eco86988, w_eco86989, w_eco86990, w_eco86991, w_eco86992, w_eco86993, w_eco86994, w_eco86995, w_eco86996, w_eco86997, w_eco86998, w_eco86999, w_eco87000, w_eco87001, w_eco87002, w_eco87003, w_eco87004, w_eco87005, w_eco87006, w_eco87007, w_eco87008, w_eco87009, w_eco87010, w_eco87011, w_eco87012, w_eco87013, w_eco87014, w_eco87015, w_eco87016, w_eco87017, w_eco87018, w_eco87019, w_eco87020, w_eco87021, w_eco87022, w_eco87023, w_eco87024, w_eco87025, w_eco87026, w_eco87027, w_eco87028, w_eco87029, w_eco87030, w_eco87031, w_eco87032, w_eco87033, w_eco87034, w_eco87035, w_eco87036, w_eco87037, w_eco87038, w_eco87039, w_eco87040, w_eco87041, w_eco87042, w_eco87043, w_eco87044, w_eco87045, w_eco87046, w_eco87047, w_eco87048, w_eco87049, w_eco87050, w_eco87051, w_eco87052, w_eco87053, w_eco87054, w_eco87055, w_eco87056, w_eco87057, w_eco87058, w_eco87059, w_eco87060, w_eco87061, w_eco87062, w_eco87063, w_eco87064, w_eco87065, w_eco87066, w_eco87067, w_eco87068, w_eco87069, w_eco87070, w_eco87071, w_eco87072, w_eco87073, w_eco87074, w_eco87075, w_eco87076, w_eco87077, w_eco87078, w_eco87079, w_eco87080, w_eco87081, w_eco87082, w_eco87083, w_eco87084, w_eco87085, w_eco87086, w_eco87087, w_eco87088, w_eco87089, w_eco87090, w_eco87091, w_eco87092, w_eco87093, w_eco87094, w_eco87095, w_eco87096, w_eco87097, w_eco87098, w_eco87099, w_eco87100, w_eco87101, w_eco87102, w_eco87103, w_eco87104, w_eco87105, w_eco87106, w_eco87107, w_eco87108, w_eco87109, w_eco87110, w_eco87111, w_eco87112, w_eco87113, w_eco87114, w_eco87115, w_eco87116, w_eco87117, w_eco87118, w_eco87119, w_eco87120, w_eco87121, w_eco87122, w_eco87123, w_eco87124, w_eco87125, w_eco87126, w_eco87127, w_eco87128, w_eco87129, w_eco87130, w_eco87131, w_eco87132, w_eco87133, w_eco87134, w_eco87135, w_eco87136, w_eco87137, w_eco87138, w_eco87139, w_eco87140, w_eco87141, w_eco87142, w_eco87143, w_eco87144, w_eco87145, w_eco87146, w_eco87147, w_eco87148, w_eco87149, w_eco87150, w_eco87151, w_eco87152, w_eco87153, w_eco87154, w_eco87155, w_eco87156, w_eco87157, w_eco87158, w_eco87159, w_eco87160, w_eco87161, w_eco87162, w_eco87163, w_eco87164, w_eco87165, w_eco87166, w_eco87167, w_eco87168, w_eco87169, w_eco87170, w_eco87171, w_eco87172, w_eco87173, w_eco87174, w_eco87175, w_eco87176, w_eco87177, w_eco87178, w_eco87179, w_eco87180, w_eco87181, w_eco87182, w_eco87183, w_eco87184, w_eco87185, w_eco87186, w_eco87187, w_eco87188, w_eco87189, w_eco87190, w_eco87191, w_eco87192, w_eco87193, w_eco87194, w_eco87195, w_eco87196, w_eco87197, w_eco87198, w_eco87199, w_eco87200, w_eco87201, w_eco87202, w_eco87203, w_eco87204, w_eco87205, w_eco87206, w_eco87207, w_eco87208, w_eco87209, w_eco87210, w_eco87211, w_eco87212, w_eco87213, w_eco87214, w_eco87215, w_eco87216, w_eco87217, w_eco87218, w_eco87219, w_eco87220, w_eco87221, w_eco87222, w_eco87223, w_eco87224, w_eco87225, w_eco87226, w_eco87227, w_eco87228, w_eco87229, w_eco87230, w_eco87231, w_eco87232, w_eco87233, w_eco87234, w_eco87235, w_eco87236, w_eco87237, w_eco87238, w_eco87239, w_eco87240, w_eco87241, w_eco87242, w_eco87243, w_eco87244, w_eco87245, w_eco87246, w_eco87247, w_eco87248, w_eco87249, w_eco87250, w_eco87251, w_eco87252, w_eco87253, w_eco87254, w_eco87255, w_eco87256, w_eco87257, w_eco87258, w_eco87259, w_eco87260, w_eco87261, w_eco87262, w_eco87263, w_eco87264, w_eco87265, w_eco87266, w_eco87267, w_eco87268, w_eco87269, w_eco87270, w_eco87271, w_eco87272, w_eco87273, w_eco87274, w_eco87275, w_eco87276, w_eco87277, w_eco87278, w_eco87279, w_eco87280, w_eco87281, w_eco87282, w_eco87283, w_eco87284, w_eco87285, w_eco87286, w_eco87287, w_eco87288, w_eco87289, w_eco87290, w_eco87291, w_eco87292, w_eco87293, w_eco87294, w_eco87295, w_eco87296, w_eco87297, w_eco87298, w_eco87299, w_eco87300, w_eco87301, w_eco87302, w_eco87303, w_eco87304, w_eco87305, w_eco87306, w_eco87307, w_eco87308, w_eco87309, w_eco87310, w_eco87311, w_eco87312, w_eco87313, w_eco87314, w_eco87315, w_eco87316, w_eco87317, w_eco87318, w_eco87319, w_eco87320, w_eco87321, w_eco87322, w_eco87323, w_eco87324, w_eco87325, w_eco87326, w_eco87327, w_eco87328, w_eco87329, w_eco87330, w_eco87331, w_eco87332, w_eco87333, w_eco87334, w_eco87335, w_eco87336, w_eco87337, w_eco87338, w_eco87339, w_eco87340, w_eco87341, w_eco87342, w_eco87343, w_eco87344, w_eco87345, w_eco87346, w_eco87347, w_eco87348, w_eco87349, w_eco87350, w_eco87351, w_eco87352, w_eco87353, w_eco87354, w_eco87355, w_eco87356, w_eco87357, w_eco87358, w_eco87359, w_eco87360, w_eco87361, w_eco87362, w_eco87363, w_eco87364, w_eco87365, w_eco87366, w_eco87367, w_eco87368, w_eco87369, w_eco87370, w_eco87371, w_eco87372, w_eco87373, w_eco87374, w_eco87375, w_eco87376, w_eco87377, w_eco87378, w_eco87379, w_eco87380, w_eco87381, w_eco87382, w_eco87383, w_eco87384, w_eco87385, w_eco87386, w_eco87387, w_eco87388, w_eco87389, w_eco87390, w_eco87391, w_eco87392, w_eco87393, w_eco87394, w_eco87395, w_eco87396, w_eco87397, w_eco87398, w_eco87399, w_eco87400, w_eco87401, w_eco87402, w_eco87403, w_eco87404, w_eco87405, w_eco87406, w_eco87407, w_eco87408, w_eco87409, w_eco87410, w_eco87411, w_eco87412, w_eco87413, w_eco87414, w_eco87415, w_eco87416, w_eco87417, w_eco87418, w_eco87419, w_eco87420, w_eco87421, w_eco87422, w_eco87423, w_eco87424, w_eco87425, w_eco87426, w_eco87427, w_eco87428, w_eco87429, w_eco87430, w_eco87431, w_eco87432, w_eco87433, w_eco87434, w_eco87435, w_eco87436, w_eco87437, w_eco87438, w_eco87439, w_eco87440, w_eco87441, w_eco87442, w_eco87443, w_eco87444, w_eco87445, w_eco87446, w_eco87447, w_eco87448, w_eco87449, w_eco87450, w_eco87451, w_eco87452, w_eco87453, w_eco87454, w_eco87455, w_eco87456, w_eco87457, w_eco87458, w_eco87459, w_eco87460, w_eco87461, w_eco87462, w_eco87463, w_eco87464, w_eco87465, w_eco87466, w_eco87467, w_eco87468, w_eco87469, w_eco87470, w_eco87471, w_eco87472, w_eco87473, w_eco87474, w_eco87475, w_eco87476, w_eco87477, w_eco87478, w_eco87479, w_eco87480, w_eco87481, w_eco87482, w_eco87483, w_eco87484, w_eco87485, w_eco87486, w_eco87487, w_eco87488, w_eco87489, w_eco87490, w_eco87491, w_eco87492, w_eco87493, w_eco87494, w_eco87495, w_eco87496, w_eco87497, w_eco87498, w_eco87499, w_eco87500, w_eco87501, w_eco87502, w_eco87503, w_eco87504, w_eco87505, w_eco87506, w_eco87507, w_eco87508, w_eco87509, w_eco87510, w_eco87511, w_eco87512, w_eco87513, w_eco87514, w_eco87515, w_eco87516, w_eco87517, w_eco87518, w_eco87519, w_eco87520, w_eco87521, w_eco87522, w_eco87523, w_eco87524, w_eco87525, w_eco87526, w_eco87527, w_eco87528, w_eco87529, w_eco87530, w_eco87531, w_eco87532, w_eco87533, w_eco87534, w_eco87535, w_eco87536, w_eco87537, w_eco87538, w_eco87539, w_eco87540, w_eco87541, w_eco87542, w_eco87543, w_eco87544, w_eco87545, w_eco87546, w_eco87547, w_eco87548, w_eco87549, w_eco87550, w_eco87551, w_eco87552, w_eco87553, w_eco87554, w_eco87555, w_eco87556, w_eco87557, w_eco87558, w_eco87559, w_eco87560, w_eco87561, w_eco87562, w_eco87563, w_eco87564, w_eco87565, w_eco87566, w_eco87567, w_eco87568, w_eco87569, w_eco87570, w_eco87571, w_eco87572, w_eco87573, w_eco87574, w_eco87575, w_eco87576, w_eco87577, w_eco87578, w_eco87579, w_eco87580, w_eco87581, w_eco87582, w_eco87583, w_eco87584, w_eco87585, w_eco87586, w_eco87587, w_eco87588, w_eco87589, w_eco87590, w_eco87591, w_eco87592, w_eco87593, w_eco87594, w_eco87595, w_eco87596, w_eco87597, w_eco87598, w_eco87599, w_eco87600, w_eco87601, w_eco87602, w_eco87603, w_eco87604, w_eco87605, w_eco87606, w_eco87607, w_eco87608, w_eco87609, w_eco87610, w_eco87611, w_eco87612, w_eco87613, w_eco87614, w_eco87615, w_eco87616, w_eco87617, w_eco87618, w_eco87619, w_eco87620, w_eco87621, w_eco87622, w_eco87623, w_eco87624, w_eco87625, w_eco87626, w_eco87627, w_eco87628, w_eco87629, w_eco87630, w_eco87631, w_eco87632, w_eco87633, w_eco87634, w_eco87635, w_eco87636, w_eco87637, w_eco87638, w_eco87639, w_eco87640, w_eco87641, w_eco87642, w_eco87643, w_eco87644, w_eco87645, w_eco87646, w_eco87647, w_eco87648, w_eco87649, w_eco87650, w_eco87651, w_eco87652, w_eco87653, w_eco87654, w_eco87655, w_eco87656, w_eco87657, w_eco87658, w_eco87659, w_eco87660, w_eco87661, w_eco87662, w_eco87663, w_eco87664, w_eco87665, w_eco87666, w_eco87667, w_eco87668, w_eco87669, w_eco87670, w_eco87671, w_eco87672, w_eco87673, w_eco87674, w_eco87675, w_eco87676, w_eco87677, w_eco87678, w_eco87679, w_eco87680, w_eco87681, w_eco87682, w_eco87683, w_eco87684, w_eco87685, w_eco87686, w_eco87687, w_eco87688, w_eco87689, w_eco87690, w_eco87691, w_eco87692, w_eco87693, w_eco87694, w_eco87695, w_eco87696, w_eco87697, w_eco87698, w_eco87699, w_eco87700, w_eco87701, w_eco87702, w_eco87703, w_eco87704, w_eco87705, w_eco87706, w_eco87707, w_eco87708, w_eco87709, w_eco87710, w_eco87711, w_eco87712, w_eco87713, w_eco87714, w_eco87715, w_eco87716, w_eco87717, w_eco87718, w_eco87719, w_eco87720, w_eco87721, w_eco87722, w_eco87723, w_eco87724, w_eco87725, w_eco87726, w_eco87727, w_eco87728, w_eco87729, w_eco87730, w_eco87731, w_eco87732, w_eco87733, w_eco87734, w_eco87735, w_eco87736, w_eco87737, w_eco87738, w_eco87739, w_eco87740, w_eco87741, w_eco87742, w_eco87743, w_eco87744, w_eco87745, w_eco87746, w_eco87747, w_eco87748, w_eco87749, w_eco87750, w_eco87751, w_eco87752, w_eco87753, w_eco87754, w_eco87755, w_eco87756, w_eco87757, w_eco87758, w_eco87759, w_eco87760, w_eco87761, w_eco87762, w_eco87763, w_eco87764, w_eco87765, w_eco87766, w_eco87767, w_eco87768, w_eco87769, w_eco87770, w_eco87771, w_eco87772, w_eco87773, w_eco87774, w_eco87775, w_eco87776, w_eco87777, w_eco87778, w_eco87779, w_eco87780, w_eco87781, w_eco87782, w_eco87783, w_eco87784, w_eco87785, w_eco87786, w_eco87787, w_eco87788, w_eco87789, w_eco87790, w_eco87791, w_eco87792, w_eco87793, w_eco87794, w_eco87795, w_eco87796, w_eco87797, w_eco87798, w_eco87799, w_eco87800, w_eco87801, w_eco87802, w_eco87803, w_eco87804, w_eco87805, w_eco87806, w_eco87807, w_eco87808, w_eco87809, w_eco87810, w_eco87811, w_eco87812, w_eco87813, w_eco87814, w_eco87815, w_eco87816, w_eco87817, w_eco87818, w_eco87819, w_eco87820, w_eco87821, w_eco87822, w_eco87823, w_eco87824, w_eco87825, w_eco87826, w_eco87827, w_eco87828, w_eco87829, w_eco87830, w_eco87831, w_eco87832, w_eco87833, w_eco87834, w_eco87835, w_eco87836, w_eco87837, w_eco87838, w_eco87839, w_eco87840, w_eco87841, w_eco87842, w_eco87843, w_eco87844, w_eco87845, w_eco87846, w_eco87847, w_eco87848, w_eco87849, w_eco87850, w_eco87851, w_eco87852, w_eco87853, w_eco87854, w_eco87855, w_eco87856, w_eco87857, w_eco87858, w_eco87859, w_eco87860, w_eco87861, w_eco87862, w_eco87863, w_eco87864, w_eco87865, w_eco87866, w_eco87867, w_eco87868, w_eco87869, w_eco87870, w_eco87871, w_eco87872, w_eco87873, w_eco87874, w_eco87875, w_eco87876, w_eco87877, w_eco87878, w_eco87879, w_eco87880, w_eco87881, w_eco87882, w_eco87883, w_eco87884, w_eco87885, w_eco87886, w_eco87887, w_eco87888, w_eco87889, w_eco87890, w_eco87891, w_eco87892, w_eco87893, w_eco87894, w_eco87895, w_eco87896, w_eco87897, w_eco87898, w_eco87899, w_eco87900, w_eco87901, w_eco87902, w_eco87903, w_eco87904, w_eco87905, w_eco87906, w_eco87907, w_eco87908, w_eco87909, w_eco87910, w_eco87911, w_eco87912, w_eco87913, w_eco87914, w_eco87915, w_eco87916, w_eco87917, w_eco87918, w_eco87919, w_eco87920, w_eco87921, w_eco87922, w_eco87923, w_eco87924, w_eco87925, w_eco87926, w_eco87927, w_eco87928, w_eco87929, w_eco87930, w_eco87931, w_eco87932, w_eco87933, w_eco87934, w_eco87935, w_eco87936, w_eco87937, w_eco87938, w_eco87939, w_eco87940, w_eco87941, w_eco87942, w_eco87943, w_eco87944, w_eco87945, w_eco87946, w_eco87947, w_eco87948, w_eco87949, w_eco87950, w_eco87951, w_eco87952, w_eco87953, w_eco87954, w_eco87955, w_eco87956, w_eco87957, w_eco87958, w_eco87959, w_eco87960, w_eco87961, w_eco87962, w_eco87963, w_eco87964, w_eco87965, w_eco87966, w_eco87967, w_eco87968, w_eco87969, w_eco87970, w_eco87971, w_eco87972, w_eco87973, w_eco87974, w_eco87975, w_eco87976, w_eco87977, w_eco87978, w_eco87979, w_eco87980, w_eco87981, w_eco87982, w_eco87983, w_eco87984, w_eco87985, w_eco87986, w_eco87987, w_eco87988, w_eco87989, w_eco87990, w_eco87991, w_eco87992, w_eco87993, w_eco87994, w_eco87995, w_eco87996, w_eco87997, w_eco87998, w_eco87999, w_eco88000, w_eco88001, w_eco88002, w_eco88003, w_eco88004, w_eco88005, w_eco88006, w_eco88007, w_eco88008, w_eco88009, w_eco88010, w_eco88011, w_eco88012, w_eco88013, w_eco88014, w_eco88015, w_eco88016, w_eco88017, w_eco88018, w_eco88019, w_eco88020, w_eco88021, w_eco88022, w_eco88023, w_eco88024, w_eco88025, w_eco88026, w_eco88027, w_eco88028, w_eco88029, w_eco88030, w_eco88031, w_eco88032, w_eco88033, w_eco88034, w_eco88035, w_eco88036, w_eco88037, w_eco88038, w_eco88039, w_eco88040, w_eco88041, w_eco88042, w_eco88043, w_eco88044, w_eco88045, w_eco88046, w_eco88047, w_eco88048, w_eco88049, w_eco88050, w_eco88051, w_eco88052, w_eco88053, w_eco88054, w_eco88055, w_eco88056, w_eco88057, w_eco88058, w_eco88059, w_eco88060, w_eco88061, w_eco88062, w_eco88063, w_eco88064, w_eco88065, w_eco88066, w_eco88067, w_eco88068, w_eco88069, w_eco88070, w_eco88071, w_eco88072, w_eco88073, w_eco88074, w_eco88075, w_eco88076, w_eco88077, w_eco88078, w_eco88079, w_eco88080, w_eco88081, w_eco88082, w_eco88083, w_eco88084, w_eco88085, w_eco88086, w_eco88087, w_eco88088, w_eco88089, w_eco88090, w_eco88091, w_eco88092, w_eco88093, w_eco88094, w_eco88095, w_eco88096, w_eco88097, w_eco88098, w_eco88099, w_eco88100, w_eco88101, w_eco88102, w_eco88103, w_eco88104, w_eco88105, w_eco88106, w_eco88107, w_eco88108, w_eco88109, w_eco88110, w_eco88111, w_eco88112, w_eco88113, w_eco88114, w_eco88115, w_eco88116, w_eco88117, w_eco88118, w_eco88119, w_eco88120, w_eco88121, w_eco88122, w_eco88123, w_eco88124, w_eco88125, w_eco88126, w_eco88127, w_eco88128, w_eco88129, w_eco88130, w_eco88131, w_eco88132, w_eco88133, w_eco88134, w_eco88135, w_eco88136, w_eco88137, w_eco88138, w_eco88139, w_eco88140, w_eco88141, w_eco88142, w_eco88143, w_eco88144, w_eco88145, w_eco88146, w_eco88147, w_eco88148, w_eco88149, w_eco88150, w_eco88151, w_eco88152, w_eco88153, w_eco88154, w_eco88155, w_eco88156, w_eco88157, w_eco88158, w_eco88159, w_eco88160, w_eco88161, w_eco88162, w_eco88163, w_eco88164, w_eco88165, w_eco88166, w_eco88167, w_eco88168, w_eco88169, w_eco88170, w_eco88171, w_eco88172, w_eco88173, w_eco88174, w_eco88175, w_eco88176, w_eco88177, w_eco88178, w_eco88179, w_eco88180, w_eco88181, w_eco88182, w_eco88183, w_eco88184, w_eco88185, w_eco88186, w_eco88187, w_eco88188, w_eco88189, w_eco88190, w_eco88191, w_eco88192, w_eco88193, w_eco88194, w_eco88195, w_eco88196, w_eco88197, w_eco88198, w_eco88199, w_eco88200, w_eco88201, w_eco88202, w_eco88203, w_eco88204, w_eco88205, w_eco88206, w_eco88207, w_eco88208, w_eco88209, w_eco88210, w_eco88211, w_eco88212, w_eco88213, w_eco88214, w_eco88215, w_eco88216, w_eco88217, w_eco88218, w_eco88219, w_eco88220, w_eco88221, w_eco88222, w_eco88223, w_eco88224, w_eco88225, w_eco88226, w_eco88227, w_eco88228, w_eco88229, w_eco88230, w_eco88231, w_eco88232, w_eco88233, w_eco88234, w_eco88235, w_eco88236, w_eco88237, w_eco88238, w_eco88239, w_eco88240, w_eco88241, w_eco88242, w_eco88243, w_eco88244, w_eco88245, w_eco88246, w_eco88247, w_eco88248, w_eco88249, w_eco88250, w_eco88251, w_eco88252, w_eco88253, w_eco88254, w_eco88255, w_eco88256, w_eco88257, w_eco88258, w_eco88259, w_eco88260, w_eco88261, w_eco88262, w_eco88263, w_eco88264, w_eco88265, w_eco88266, w_eco88267, w_eco88268, w_eco88269, w_eco88270, w_eco88271, w_eco88272, w_eco88273, w_eco88274, w_eco88275, w_eco88276, w_eco88277, w_eco88278, w_eco88279, w_eco88280, w_eco88281, w_eco88282, w_eco88283, w_eco88284, w_eco88285, w_eco88286, w_eco88287, w_eco88288, w_eco88289, w_eco88290, w_eco88291, w_eco88292, w_eco88293, w_eco88294, w_eco88295, w_eco88296, w_eco88297, w_eco88298, w_eco88299, w_eco88300, w_eco88301, w_eco88302, w_eco88303, w_eco88304, w_eco88305, w_eco88306, w_eco88307, w_eco88308, w_eco88309, w_eco88310, w_eco88311, w_eco88312, w_eco88313, w_eco88314, w_eco88315, w_eco88316, w_eco88317, w_eco88318, w_eco88319, w_eco88320, w_eco88321, w_eco88322, w_eco88323, w_eco88324, w_eco88325, w_eco88326, w_eco88327, w_eco88328, w_eco88329, w_eco88330, w_eco88331, w_eco88332, w_eco88333, w_eco88334, w_eco88335, w_eco88336, w_eco88337, w_eco88338, w_eco88339, w_eco88340, w_eco88341, w_eco88342, w_eco88343, w_eco88344, w_eco88345, w_eco88346, w_eco88347, w_eco88348, w_eco88349, w_eco88350, w_eco88351, w_eco88352, w_eco88353, w_eco88354, w_eco88355, w_eco88356, w_eco88357, w_eco88358, w_eco88359, w_eco88360, w_eco88361, w_eco88362, w_eco88363, w_eco88364, w_eco88365, w_eco88366, w_eco88367, w_eco88368, w_eco88369, w_eco88370, w_eco88371, w_eco88372, w_eco88373, w_eco88374, w_eco88375, w_eco88376, w_eco88377, w_eco88378, w_eco88379, w_eco88380, w_eco88381, w_eco88382, w_eco88383, w_eco88384, w_eco88385, w_eco88386, w_eco88387, w_eco88388, w_eco88389, w_eco88390, w_eco88391, w_eco88392, w_eco88393, w_eco88394, w_eco88395, w_eco88396, w_eco88397, w_eco88398, w_eco88399, w_eco88400, w_eco88401, w_eco88402, w_eco88403, w_eco88404, w_eco88405, w_eco88406, w_eco88407, w_eco88408, w_eco88409, w_eco88410, w_eco88411, w_eco88412, w_eco88413, w_eco88414, w_eco88415, w_eco88416, w_eco88417, w_eco88418, w_eco88419, w_eco88420, w_eco88421, w_eco88422, w_eco88423, w_eco88424, w_eco88425, w_eco88426, w_eco88427, w_eco88428, w_eco88429, w_eco88430, w_eco88431, w_eco88432, w_eco88433, w_eco88434, w_eco88435, w_eco88436, w_eco88437, w_eco88438, w_eco88439, w_eco88440, w_eco88441, w_eco88442, w_eco88443, w_eco88444, w_eco88445, w_eco88446, w_eco88447, w_eco88448, w_eco88449, w_eco88450, w_eco88451, w_eco88452, w_eco88453, w_eco88454, w_eco88455, w_eco88456, w_eco88457, w_eco88458, w_eco88459, w_eco88460, w_eco88461, w_eco88462, w_eco88463, w_eco88464, w_eco88465, w_eco88466, w_eco88467, w_eco88468, w_eco88469, w_eco88470, w_eco88471, w_eco88472, w_eco88473, w_eco88474, w_eco88475, w_eco88476, w_eco88477, w_eco88478, w_eco88479, w_eco88480, w_eco88481, w_eco88482, w_eco88483, w_eco88484, w_eco88485, w_eco88486, w_eco88487, w_eco88488, w_eco88489, w_eco88490, w_eco88491, w_eco88492, w_eco88493, w_eco88494, w_eco88495, w_eco88496, w_eco88497, w_eco88498, w_eco88499, w_eco88500, w_eco88501, w_eco88502, w_eco88503, w_eco88504, w_eco88505, w_eco88506, w_eco88507, w_eco88508, w_eco88509, w_eco88510, w_eco88511, w_eco88512, w_eco88513, w_eco88514, w_eco88515, w_eco88516, w_eco88517, w_eco88518, w_eco88519, w_eco88520, w_eco88521, w_eco88522, w_eco88523, w_eco88524, w_eco88525, w_eco88526, w_eco88527, w_eco88528, w_eco88529, w_eco88530, w_eco88531, w_eco88532, w_eco88533, w_eco88534, w_eco88535, w_eco88536, w_eco88537, w_eco88538, w_eco88539, w_eco88540, w_eco88541, w_eco88542, w_eco88543, w_eco88544, w_eco88545, w_eco88546, w_eco88547, w_eco88548, w_eco88549, w_eco88550, w_eco88551, w_eco88552, w_eco88553, w_eco88554, w_eco88555, w_eco88556, w_eco88557, w_eco88558, w_eco88559, w_eco88560, w_eco88561, w_eco88562, w_eco88563, w_eco88564, w_eco88565, w_eco88566, w_eco88567, w_eco88568, w_eco88569, w_eco88570, w_eco88571, w_eco88572, w_eco88573, w_eco88574, w_eco88575, w_eco88576, w_eco88577, w_eco88578, w_eco88579, w_eco88580, w_eco88581, w_eco88582, w_eco88583, w_eco88584, w_eco88585, w_eco88586, w_eco88587, w_eco88588, w_eco88589, w_eco88590, w_eco88591, w_eco88592, w_eco88593, w_eco88594, w_eco88595, w_eco88596, w_eco88597, w_eco88598, w_eco88599, w_eco88600, w_eco88601, w_eco88602, w_eco88603, w_eco88604, w_eco88605, w_eco88606, w_eco88607, w_eco88608, w_eco88609, w_eco88610, w_eco88611, w_eco88612, w_eco88613, w_eco88614, w_eco88615, w_eco88616, w_eco88617, w_eco88618, w_eco88619, w_eco88620, w_eco88621, w_eco88622, w_eco88623, w_eco88624, w_eco88625, w_eco88626, w_eco88627, w_eco88628, w_eco88629, w_eco88630, w_eco88631, w_eco88632, w_eco88633, w_eco88634, w_eco88635, w_eco88636, w_eco88637, w_eco88638, w_eco88639, w_eco88640, w_eco88641, w_eco88642, w_eco88643, w_eco88644, w_eco88645, w_eco88646, w_eco88647, w_eco88648, w_eco88649, w_eco88650, w_eco88651, w_eco88652, w_eco88653, w_eco88654, w_eco88655, w_eco88656, w_eco88657, w_eco88658, w_eco88659, w_eco88660, w_eco88661, w_eco88662, w_eco88663, w_eco88664, w_eco88665, w_eco88666, w_eco88667, w_eco88668, w_eco88669, w_eco88670, w_eco88671, w_eco88672, w_eco88673, w_eco88674, w_eco88675, w_eco88676, w_eco88677, w_eco88678, w_eco88679, w_eco88680, w_eco88681, w_eco88682, w_eco88683, w_eco88684, w_eco88685, w_eco88686, w_eco88687, w_eco88688, w_eco88689, w_eco88690, w_eco88691, w_eco88692, w_eco88693, w_eco88694, w_eco88695, w_eco88696, w_eco88697, w_eco88698, w_eco88699, w_eco88700, w_eco88701, w_eco88702, w_eco88703, w_eco88704, w_eco88705, w_eco88706, w_eco88707, w_eco88708, w_eco88709, w_eco88710, w_eco88711, w_eco88712, w_eco88713, w_eco88714, w_eco88715, w_eco88716, w_eco88717, w_eco88718, w_eco88719, w_eco88720, w_eco88721, w_eco88722, w_eco88723, w_eco88724, w_eco88725, w_eco88726, w_eco88727, w_eco88728, w_eco88729, w_eco88730, w_eco88731, w_eco88732, w_eco88733, w_eco88734, w_eco88735, w_eco88736, w_eco88737, w_eco88738, w_eco88739, w_eco88740, w_eco88741, w_eco88742, w_eco88743, w_eco88744, w_eco88745, w_eco88746, w_eco88747, w_eco88748, w_eco88749, w_eco88750, w_eco88751, w_eco88752, w_eco88753, w_eco88754, w_eco88755, w_eco88756, w_eco88757, w_eco88758, w_eco88759, w_eco88760, w_eco88761, w_eco88762, w_eco88763, w_eco88764, w_eco88765, w_eco88766, w_eco88767, w_eco88768, w_eco88769, w_eco88770, w_eco88771, w_eco88772, w_eco88773, w_eco88774, w_eco88775, w_eco88776, w_eco88777, w_eco88778, w_eco88779, w_eco88780, w_eco88781, w_eco88782, w_eco88783, w_eco88784, w_eco88785, w_eco88786, w_eco88787, w_eco88788, w_eco88789, w_eco88790, w_eco88791, w_eco88792, w_eco88793, w_eco88794, w_eco88795, w_eco88796, w_eco88797, w_eco88798, w_eco88799, w_eco88800, w_eco88801, w_eco88802, w_eco88803, w_eco88804, w_eco88805, w_eco88806, w_eco88807, w_eco88808, w_eco88809, w_eco88810, w_eco88811, w_eco88812, w_eco88813, w_eco88814, w_eco88815, w_eco88816, w_eco88817, w_eco88818, w_eco88819, w_eco88820, w_eco88821, w_eco88822, w_eco88823, w_eco88824, w_eco88825, w_eco88826, w_eco88827, w_eco88828, w_eco88829, w_eco88830, w_eco88831, w_eco88832, w_eco88833, w_eco88834, w_eco88835, w_eco88836, w_eco88837, w_eco88838, w_eco88839, w_eco88840, w_eco88841, w_eco88842, w_eco88843, w_eco88844, w_eco88845, w_eco88846, w_eco88847, w_eco88848, w_eco88849, w_eco88850, w_eco88851, w_eco88852, w_eco88853, w_eco88854, w_eco88855, w_eco88856, w_eco88857, w_eco88858, w_eco88859, w_eco88860, w_eco88861, w_eco88862, w_eco88863, w_eco88864, w_eco88865, w_eco88866, w_eco88867, w_eco88868, w_eco88869, w_eco88870, w_eco88871, w_eco88872, w_eco88873, w_eco88874, w_eco88875, w_eco88876, w_eco88877, w_eco88878, w_eco88879, w_eco88880, w_eco88881, w_eco88882, w_eco88883, w_eco88884, w_eco88885, w_eco88886, w_eco88887, w_eco88888, w_eco88889, w_eco88890, w_eco88891, w_eco88892, w_eco88893, w_eco88894, w_eco88895, w_eco88896, w_eco88897, w_eco88898, w_eco88899, w_eco88900, w_eco88901, w_eco88902, w_eco88903, w_eco88904, w_eco88905, w_eco88906, w_eco88907, w_eco88908, w_eco88909, w_eco88910, w_eco88911, w_eco88912, w_eco88913, w_eco88914, w_eco88915, w_eco88916, w_eco88917, w_eco88918, w_eco88919, w_eco88920, w_eco88921, w_eco88922, w_eco88923, w_eco88924, w_eco88925, w_eco88926, w_eco88927, w_eco88928, w_eco88929, w_eco88930, w_eco88931, w_eco88932, w_eco88933, w_eco88934, w_eco88935, w_eco88936, w_eco88937, w_eco88938, w_eco88939, w_eco88940, w_eco88941, w_eco88942, w_eco88943, w_eco88944, w_eco88945, w_eco88946, w_eco88947, w_eco88948, w_eco88949, w_eco88950, w_eco88951, w_eco88952, w_eco88953, w_eco88954, w_eco88955, w_eco88956, w_eco88957, w_eco88958, w_eco88959, w_eco88960, w_eco88961, w_eco88962, w_eco88963, w_eco88964, w_eco88965, w_eco88966, w_eco88967, w_eco88968, w_eco88969, w_eco88970, w_eco88971, w_eco88972, w_eco88973, w_eco88974, w_eco88975, w_eco88976, w_eco88977, w_eco88978, w_eco88979, w_eco88980, w_eco88981, w_eco88982, w_eco88983, w_eco88984, w_eco88985, w_eco88986, w_eco88987, w_eco88988, w_eco88989, w_eco88990, w_eco88991, w_eco88992, w_eco88993, w_eco88994, w_eco88995, w_eco88996, w_eco88997, w_eco88998, w_eco88999, w_eco89000, w_eco89001, w_eco89002, w_eco89003, w_eco89004, w_eco89005, w_eco89006, w_eco89007, w_eco89008, w_eco89009, w_eco89010, w_eco89011, w_eco89012, w_eco89013, w_eco89014, w_eco89015, w_eco89016, w_eco89017, w_eco89018, w_eco89019, w_eco89020, w_eco89021, w_eco89022, w_eco89023, w_eco89024, w_eco89025, w_eco89026, w_eco89027, w_eco89028, w_eco89029, w_eco89030, w_eco89031, w_eco89032, w_eco89033, w_eco89034, w_eco89035, w_eco89036, w_eco89037, w_eco89038, w_eco89039, w_eco89040, w_eco89041, w_eco89042, w_eco89043, w_eco89044, w_eco89045, w_eco89046, w_eco89047, w_eco89048, w_eco89049, w_eco89050, w_eco89051, w_eco89052, w_eco89053, w_eco89054, w_eco89055, w_eco89056, w_eco89057, w_eco89058, w_eco89059, w_eco89060, w_eco89061, w_eco89062, w_eco89063, w_eco89064, w_eco89065, w_eco89066, w_eco89067, w_eco89068, w_eco89069, w_eco89070, w_eco89071, w_eco89072, w_eco89073, w_eco89074, w_eco89075, w_eco89076, w_eco89077, w_eco89078, w_eco89079, w_eco89080, w_eco89081, w_eco89082, w_eco89083, w_eco89084, w_eco89085, w_eco89086, w_eco89087, w_eco89088, w_eco89089, w_eco89090, w_eco89091, w_eco89092, w_eco89093, w_eco89094, w_eco89095, w_eco89096, w_eco89097, w_eco89098, w_eco89099, w_eco89100, w_eco89101, w_eco89102, w_eco89103, w_eco89104, w_eco89105, w_eco89106, w_eco89107, w_eco89108, w_eco89109, w_eco89110, w_eco89111, w_eco89112, w_eco89113, w_eco89114, w_eco89115, w_eco89116, w_eco89117, w_eco89118, w_eco89119, w_eco89120, w_eco89121, w_eco89122, w_eco89123, w_eco89124, w_eco89125, w_eco89126, w_eco89127, w_eco89128, w_eco89129, w_eco89130, w_eco89131, w_eco89132, w_eco89133, w_eco89134, w_eco89135, w_eco89136, w_eco89137, w_eco89138, w_eco89139, w_eco89140, w_eco89141, w_eco89142, w_eco89143, w_eco89144, w_eco89145, w_eco89146, w_eco89147, w_eco89148, w_eco89149, w_eco89150, w_eco89151, w_eco89152, w_eco89153, w_eco89154, w_eco89155, w_eco89156, w_eco89157, w_eco89158, w_eco89159, w_eco89160, w_eco89161, w_eco89162, w_eco89163, w_eco89164, w_eco89165, w_eco89166, w_eco89167, w_eco89168, w_eco89169, w_eco89170, w_eco89171, w_eco89172, w_eco89173, w_eco89174, w_eco89175, w_eco89176, w_eco89177, w_eco89178, w_eco89179, w_eco89180, w_eco89181, w_eco89182, w_eco89183, w_eco89184, w_eco89185, w_eco89186, w_eco89187, w_eco89188, w_eco89189, w_eco89190, w_eco89191, w_eco89192, w_eco89193, w_eco89194, w_eco89195, w_eco89196, w_eco89197, w_eco89198, w_eco89199, w_eco89200, w_eco89201, w_eco89202, w_eco89203, w_eco89204, w_eco89205, w_eco89206, w_eco89207, w_eco89208, w_eco89209, w_eco89210, w_eco89211, w_eco89212, w_eco89213, w_eco89214, w_eco89215, w_eco89216, w_eco89217, w_eco89218, w_eco89219, w_eco89220, w_eco89221, w_eco89222, w_eco89223, w_eco89224, w_eco89225, w_eco89226, w_eco89227, w_eco89228, w_eco89229, w_eco89230, w_eco89231, w_eco89232, w_eco89233, w_eco89234, w_eco89235, w_eco89236, w_eco89237, w_eco89238, w_eco89239, w_eco89240, w_eco89241, w_eco89242, w_eco89243, w_eco89244, w_eco89245, w_eco89246, w_eco89247, w_eco89248, w_eco89249, w_eco89250, w_eco89251, w_eco89252, w_eco89253, w_eco89254, w_eco89255, w_eco89256, w_eco89257, w_eco89258, w_eco89259, w_eco89260, w_eco89261, w_eco89262, w_eco89263, w_eco89264, w_eco89265, w_eco89266, w_eco89267, w_eco89268, w_eco89269, w_eco89270, w_eco89271, w_eco89272, w_eco89273, w_eco89274, w_eco89275, w_eco89276, w_eco89277, w_eco89278, w_eco89279, w_eco89280, w_eco89281, w_eco89282, w_eco89283, w_eco89284, w_eco89285, w_eco89286, w_eco89287, w_eco89288, w_eco89289, w_eco89290, w_eco89291, w_eco89292, w_eco89293, w_eco89294, w_eco89295, w_eco89296, w_eco89297, w_eco89298, w_eco89299, w_eco89300, w_eco89301, w_eco89302, w_eco89303, w_eco89304, w_eco89305, w_eco89306, w_eco89307, w_eco89308, w_eco89309, w_eco89310, w_eco89311, w_eco89312, w_eco89313, w_eco89314, w_eco89315, w_eco89316, w_eco89317, w_eco89318, w_eco89319, w_eco89320, w_eco89321, w_eco89322, w_eco89323, w_eco89324, w_eco89325, w_eco89326, w_eco89327, w_eco89328, w_eco89329, w_eco89330, w_eco89331, w_eco89332, w_eco89333, w_eco89334, w_eco89335, w_eco89336, w_eco89337, w_eco89338, w_eco89339, w_eco89340, w_eco89341, w_eco89342, w_eco89343, w_eco89344, w_eco89345, w_eco89346, w_eco89347, w_eco89348, w_eco89349, w_eco89350, w_eco89351, w_eco89352, w_eco89353, w_eco89354, w_eco89355, w_eco89356, w_eco89357, w_eco89358, w_eco89359, w_eco89360, w_eco89361, w_eco89362, w_eco89363, w_eco89364, w_eco89365, w_eco89366, w_eco89367, w_eco89368, w_eco89369, w_eco89370, w_eco89371, w_eco89372, w_eco89373, w_eco89374, w_eco89375, w_eco89376, w_eco89377, w_eco89378, w_eco89379, w_eco89380, w_eco89381, w_eco89382, w_eco89383, w_eco89384, w_eco89385, w_eco89386, w_eco89387, w_eco89388, w_eco89389, w_eco89390, w_eco89391, w_eco89392, w_eco89393, w_eco89394, w_eco89395, w_eco89396, w_eco89397, w_eco89398, w_eco89399, w_eco89400, w_eco89401, w_eco89402, w_eco89403, w_eco89404, w_eco89405, w_eco89406, w_eco89407, w_eco89408, w_eco89409, w_eco89410, w_eco89411, w_eco89412, w_eco89413, w_eco89414, w_eco89415, w_eco89416, w_eco89417, w_eco89418, w_eco89419, w_eco89420, w_eco89421, w_eco89422, w_eco89423, w_eco89424, w_eco89425, w_eco89426, w_eco89427, w_eco89428, w_eco89429, w_eco89430, w_eco89431, w_eco89432, w_eco89433, w_eco89434, w_eco89435, w_eco89436, w_eco89437, w_eco89438, w_eco89439, w_eco89440, w_eco89441, w_eco89442, w_eco89443, w_eco89444, w_eco89445, w_eco89446, w_eco89447, w_eco89448, w_eco89449, w_eco89450, w_eco89451, w_eco89452, w_eco89453, w_eco89454, w_eco89455, w_eco89456, w_eco89457, w_eco89458, w_eco89459, w_eco89460, w_eco89461, w_eco89462, w_eco89463, w_eco89464, w_eco89465, w_eco89466, w_eco89467, w_eco89468, w_eco89469, w_eco89470, w_eco89471, w_eco89472, w_eco89473, w_eco89474, w_eco89475, w_eco89476, w_eco89477, w_eco89478, w_eco89479, w_eco89480, w_eco89481, w_eco89482, w_eco89483, w_eco89484, w_eco89485, w_eco89486, w_eco89487, w_eco89488, w_eco89489, w_eco89490, w_eco89491, w_eco89492, w_eco89493, w_eco89494, w_eco89495, w_eco89496, w_eco89497, w_eco89498, w_eco89499, w_eco89500, w_eco89501, w_eco89502, w_eco89503, w_eco89504, w_eco89505, w_eco89506, w_eco89507, w_eco89508, w_eco89509, w_eco89510, w_eco89511, w_eco89512, w_eco89513, w_eco89514, w_eco89515, w_eco89516, w_eco89517, w_eco89518, w_eco89519, w_eco89520, w_eco89521, w_eco89522, w_eco89523, w_eco89524, w_eco89525, w_eco89526, w_eco89527, w_eco89528, w_eco89529, w_eco89530, w_eco89531, w_eco89532, w_eco89533, w_eco89534, w_eco89535, w_eco89536, w_eco89537, w_eco89538, w_eco89539, w_eco89540, w_eco89541, w_eco89542, w_eco89543, w_eco89544, w_eco89545, w_eco89546, w_eco89547, w_eco89548, w_eco89549, w_eco89550, w_eco89551, w_eco89552, w_eco89553, w_eco89554, w_eco89555, w_eco89556, w_eco89557, w_eco89558, w_eco89559, w_eco89560, w_eco89561, w_eco89562, w_eco89563, w_eco89564, w_eco89565, w_eco89566, w_eco89567, w_eco89568, w_eco89569, w_eco89570, w_eco89571, w_eco89572, w_eco89573, w_eco89574, w_eco89575, w_eco89576, w_eco89577, w_eco89578, w_eco89579, w_eco89580, w_eco89581, w_eco89582, w_eco89583, w_eco89584, w_eco89585, w_eco89586, w_eco89587, w_eco89588, w_eco89589, w_eco89590, w_eco89591, w_eco89592, w_eco89593, w_eco89594, w_eco89595, w_eco89596, w_eco89597, w_eco89598, w_eco89599, w_eco89600, w_eco89601, w_eco89602, w_eco89603, w_eco89604, w_eco89605, w_eco89606, w_eco89607, w_eco89608, w_eco89609, w_eco89610, w_eco89611, w_eco89612, w_eco89613, w_eco89614, w_eco89615, w_eco89616, w_eco89617, w_eco89618, w_eco89619, w_eco89620, w_eco89621, w_eco89622, w_eco89623, w_eco89624, w_eco89625, w_eco89626, w_eco89627, w_eco89628, w_eco89629, w_eco89630, w_eco89631, w_eco89632, w_eco89633, w_eco89634, w_eco89635, w_eco89636, w_eco89637, w_eco89638, w_eco89639, w_eco89640, w_eco89641, w_eco89642, w_eco89643, w_eco89644, w_eco89645, w_eco89646, w_eco89647, w_eco89648, w_eco89649, w_eco89650, w_eco89651, w_eco89652, w_eco89653, w_eco89654, w_eco89655, w_eco89656, w_eco89657, w_eco89658, w_eco89659, w_eco89660, w_eco89661, w_eco89662, w_eco89663, w_eco89664, w_eco89665, w_eco89666, w_eco89667, w_eco89668, w_eco89669, w_eco89670, w_eco89671, w_eco89672, w_eco89673, w_eco89674, w_eco89675, w_eco89676, w_eco89677, w_eco89678, w_eco89679, w_eco89680, w_eco89681, w_eco89682, w_eco89683, w_eco89684, w_eco89685, w_eco89686, w_eco89687, w_eco89688, w_eco89689, w_eco89690, w_eco89691, w_eco89692, w_eco89693, w_eco89694, w_eco89695, w_eco89696, w_eco89697, w_eco89698, w_eco89699, w_eco89700, w_eco89701, w_eco89702, w_eco89703, w_eco89704, w_eco89705, w_eco89706, w_eco89707, w_eco89708, w_eco89709, w_eco89710, w_eco89711, w_eco89712, w_eco89713, w_eco89714, w_eco89715, w_eco89716, w_eco89717, w_eco89718, w_eco89719, w_eco89720, w_eco89721, w_eco89722, w_eco89723, w_eco89724, w_eco89725, w_eco89726, w_eco89727, w_eco89728, w_eco89729, w_eco89730, w_eco89731, w_eco89732, w_eco89733, w_eco89734, w_eco89735, w_eco89736, w_eco89737, w_eco89738, w_eco89739, w_eco89740, w_eco89741, w_eco89742, w_eco89743, w_eco89744, w_eco89745, w_eco89746, w_eco89747, w_eco89748, w_eco89749, w_eco89750, w_eco89751, w_eco89752, w_eco89753, w_eco89754, w_eco89755, w_eco89756, w_eco89757, w_eco89758, w_eco89759, w_eco89760, w_eco89761, w_eco89762, w_eco89763, w_eco89764, w_eco89765, w_eco89766, w_eco89767, w_eco89768, w_eco89769, w_eco89770, w_eco89771, w_eco89772, w_eco89773, w_eco89774, w_eco89775, w_eco89776, w_eco89777, w_eco89778, w_eco89779, w_eco89780, w_eco89781, w_eco89782, w_eco89783, w_eco89784, w_eco89785, w_eco89786, w_eco89787, w_eco89788, w_eco89789, w_eco89790, w_eco89791, w_eco89792, w_eco89793, w_eco89794, w_eco89795, w_eco89796, w_eco89797, w_eco89798, w_eco89799, w_eco89800, w_eco89801, w_eco89802, w_eco89803, w_eco89804, w_eco89805, w_eco89806, w_eco89807, w_eco89808, w_eco89809, w_eco89810, w_eco89811, w_eco89812, w_eco89813, w_eco89814, w_eco89815, w_eco89816, w_eco89817, w_eco89818, w_eco89819, w_eco89820, w_eco89821, w_eco89822, w_eco89823, w_eco89824, w_eco89825, w_eco89826, w_eco89827, w_eco89828, w_eco89829, w_eco89830, w_eco89831, w_eco89832, w_eco89833, w_eco89834, w_eco89835, w_eco89836, w_eco89837, w_eco89838, w_eco89839, w_eco89840, w_eco89841, w_eco89842, w_eco89843, w_eco89844, w_eco89845, w_eco89846, w_eco89847, w_eco89848, w_eco89849, w_eco89850, w_eco89851, w_eco89852, w_eco89853, w_eco89854, w_eco89855, w_eco89856, w_eco89857, w_eco89858, w_eco89859, w_eco89860, w_eco89861, w_eco89862, w_eco89863, w_eco89864, w_eco89865, w_eco89866, w_eco89867, w_eco89868, w_eco89869, w_eco89870, w_eco89871, w_eco89872, w_eco89873, w_eco89874, w_eco89875, w_eco89876, w_eco89877, w_eco89878, w_eco89879, w_eco89880, w_eco89881, w_eco89882, w_eco89883, w_eco89884, w_eco89885, w_eco89886, w_eco89887, w_eco89888, w_eco89889, w_eco89890, w_eco89891, w_eco89892, w_eco89893, w_eco89894, w_eco89895, w_eco89896, w_eco89897, w_eco89898, w_eco89899, w_eco89900, w_eco89901, w_eco89902, w_eco89903, w_eco89904, w_eco89905, w_eco89906, w_eco89907, w_eco89908, w_eco89909, w_eco89910, w_eco89911, w_eco89912, w_eco89913, w_eco89914, w_eco89915, w_eco89916, w_eco89917, w_eco89918, w_eco89919, w_eco89920, w_eco89921, w_eco89922, w_eco89923, w_eco89924, w_eco89925, w_eco89926, w_eco89927, w_eco89928, w_eco89929, w_eco89930, w_eco89931, w_eco89932, w_eco89933, w_eco89934, w_eco89935, w_eco89936, w_eco89937, w_eco89938, w_eco89939, w_eco89940, w_eco89941, w_eco89942, w_eco89943, w_eco89944, w_eco89945, w_eco89946, w_eco89947, w_eco89948, w_eco89949, w_eco89950, w_eco89951, w_eco89952, w_eco89953, w_eco89954, w_eco89955, w_eco89956, w_eco89957, w_eco89958, w_eco89959, w_eco89960, w_eco89961, w_eco89962, w_eco89963, w_eco89964, w_eco89965, w_eco89966, w_eco89967, w_eco89968, w_eco89969, w_eco89970, w_eco89971, w_eco89972, w_eco89973, w_eco89974, w_eco89975, w_eco89976, w_eco89977, w_eco89978, w_eco89979, w_eco89980, w_eco89981, w_eco89982, w_eco89983, w_eco89984, w_eco89985, w_eco89986, w_eco89987, w_eco89988, w_eco89989, w_eco89990, w_eco89991, w_eco89992, w_eco89993, w_eco89994, w_eco89995, w_eco89996, w_eco89997, w_eco89998, w_eco89999, w_eco90000, w_eco90001, w_eco90002, w_eco90003, w_eco90004, w_eco90005, w_eco90006, w_eco90007, w_eco90008, w_eco90009, w_eco90010, w_eco90011, w_eco90012, w_eco90013, w_eco90014, w_eco90015, w_eco90016, w_eco90017, w_eco90018, w_eco90019, w_eco90020, w_eco90021, w_eco90022, w_eco90023, w_eco90024, w_eco90025, w_eco90026, w_eco90027, w_eco90028, w_eco90029, w_eco90030, w_eco90031, w_eco90032, w_eco90033, w_eco90034, w_eco90035, w_eco90036, w_eco90037, w_eco90038, w_eco90039, w_eco90040, w_eco90041, w_eco90042, w_eco90043, w_eco90044, w_eco90045, w_eco90046, w_eco90047, w_eco90048, w_eco90049, w_eco90050, w_eco90051, w_eco90052, w_eco90053, w_eco90054, w_eco90055, w_eco90056, w_eco90057, w_eco90058, w_eco90059, w_eco90060, w_eco90061, w_eco90062, w_eco90063, w_eco90064, w_eco90065, w_eco90066, w_eco90067, w_eco90068, w_eco90069, w_eco90070, w_eco90071, w_eco90072, w_eco90073, w_eco90074, w_eco90075, w_eco90076, w_eco90077, w_eco90078, w_eco90079, w_eco90080, w_eco90081, w_eco90082, w_eco90083, w_eco90084, w_eco90085, w_eco90086, w_eco90087, w_eco90088, w_eco90089, w_eco90090, w_eco90091, w_eco90092, w_eco90093, w_eco90094, w_eco90095, w_eco90096, w_eco90097, w_eco90098, w_eco90099, w_eco90100, w_eco90101, w_eco90102, w_eco90103, w_eco90104, w_eco90105, w_eco90106, w_eco90107, w_eco90108, w_eco90109, w_eco90110, w_eco90111, w_eco90112, w_eco90113, w_eco90114, w_eco90115, w_eco90116, w_eco90117, w_eco90118, w_eco90119, w_eco90120, w_eco90121, w_eco90122, w_eco90123, w_eco90124, w_eco90125, w_eco90126, w_eco90127, w_eco90128, w_eco90129, w_eco90130, w_eco90131, w_eco90132, w_eco90133, w_eco90134, w_eco90135, w_eco90136, w_eco90137, w_eco90138, w_eco90139, w_eco90140, w_eco90141, w_eco90142, w_eco90143, w_eco90144, w_eco90145, w_eco90146, w_eco90147, w_eco90148, w_eco90149, w_eco90150, w_eco90151, w_eco90152, w_eco90153, w_eco90154, w_eco90155, w_eco90156, w_eco90157, w_eco90158, w_eco90159, w_eco90160, w_eco90161, w_eco90162, w_eco90163, w_eco90164, w_eco90165, w_eco90166, w_eco90167, w_eco90168, w_eco90169, w_eco90170, w_eco90171, w_eco90172, w_eco90173, w_eco90174, w_eco90175, w_eco90176, w_eco90177, w_eco90178, w_eco90179, w_eco90180, w_eco90181, w_eco90182, w_eco90183, w_eco90184, w_eco90185, w_eco90186, w_eco90187, w_eco90188, w_eco90189, w_eco90190, w_eco90191, w_eco90192, w_eco90193, w_eco90194, w_eco90195, w_eco90196, w_eco90197, w_eco90198, w_eco90199, w_eco90200, w_eco90201, w_eco90202, w_eco90203, w_eco90204, w_eco90205, w_eco90206, w_eco90207, w_eco90208, w_eco90209, w_eco90210, w_eco90211, w_eco90212, w_eco90213, w_eco90214, w_eco90215, w_eco90216, w_eco90217, w_eco90218, w_eco90219, w_eco90220, w_eco90221, w_eco90222, w_eco90223, w_eco90224, w_eco90225, w_eco90226, w_eco90227, w_eco90228, w_eco90229, w_eco90230, w_eco90231, w_eco90232, w_eco90233, w_eco90234, w_eco90235, w_eco90236, w_eco90237, w_eco90238, w_eco90239, w_eco90240, w_eco90241, w_eco90242, w_eco90243, w_eco90244, w_eco90245, w_eco90246, w_eco90247, w_eco90248, w_eco90249, w_eco90250, w_eco90251, w_eco90252, w_eco90253, w_eco90254, w_eco90255, w_eco90256, w_eco90257, w_eco90258, w_eco90259, w_eco90260, w_eco90261, w_eco90262, w_eco90263, w_eco90264, w_eco90265, w_eco90266, w_eco90267, w_eco90268, w_eco90269, w_eco90270, w_eco90271, w_eco90272, w_eco90273, w_eco90274, w_eco90275, w_eco90276, w_eco90277, w_eco90278, w_eco90279, w_eco90280, w_eco90281, w_eco90282, w_eco90283, w_eco90284, w_eco90285, w_eco90286, w_eco90287, w_eco90288, w_eco90289, w_eco90290, w_eco90291, w_eco90292, w_eco90293, w_eco90294, w_eco90295, w_eco90296, w_eco90297, w_eco90298, w_eco90299, w_eco90300, w_eco90301, w_eco90302, w_eco90303, w_eco90304, w_eco90305, w_eco90306, w_eco90307, w_eco90308, w_eco90309, w_eco90310, w_eco90311, w_eco90312, w_eco90313, w_eco90314, w_eco90315, w_eco90316, w_eco90317, w_eco90318, w_eco90319, w_eco90320, w_eco90321, w_eco90322, w_eco90323, w_eco90324, w_eco90325, w_eco90326, w_eco90327, w_eco90328, w_eco90329, w_eco90330, w_eco90331, w_eco90332, w_eco90333, w_eco90334, w_eco90335, w_eco90336, w_eco90337, w_eco90338, w_eco90339, w_eco90340, w_eco90341, w_eco90342, w_eco90343, w_eco90344, w_eco90345, w_eco90346, w_eco90347, w_eco90348, w_eco90349, w_eco90350, w_eco90351, w_eco90352, w_eco90353, w_eco90354, w_eco90355, w_eco90356, w_eco90357, w_eco90358, w_eco90359, w_eco90360, w_eco90361, w_eco90362, w_eco90363, w_eco90364, w_eco90365, w_eco90366, w_eco90367, w_eco90368, w_eco90369, w_eco90370, w_eco90371, w_eco90372, w_eco90373, w_eco90374, w_eco90375, w_eco90376, w_eco90377, w_eco90378, w_eco90379, w_eco90380, w_eco90381, w_eco90382, w_eco90383, w_eco90384, w_eco90385, w_eco90386, w_eco90387, w_eco90388, w_eco90389, w_eco90390, w_eco90391, w_eco90392, w_eco90393, w_eco90394, w_eco90395, w_eco90396, w_eco90397, w_eco90398, w_eco90399, w_eco90400, w_eco90401, w_eco90402, w_eco90403, w_eco90404, w_eco90405, w_eco90406, w_eco90407, w_eco90408, w_eco90409, w_eco90410, w_eco90411, w_eco90412, w_eco90413, w_eco90414, w_eco90415, w_eco90416, w_eco90417, w_eco90418, w_eco90419, w_eco90420, w_eco90421, w_eco90422, w_eco90423, w_eco90424, w_eco90425, w_eco90426, w_eco90427, w_eco90428, w_eco90429, w_eco90430, w_eco90431, w_eco90432, w_eco90433, w_eco90434, w_eco90435, w_eco90436, w_eco90437, w_eco90438, w_eco90439, w_eco90440, w_eco90441, w_eco90442, w_eco90443, w_eco90444, w_eco90445, w_eco90446, w_eco90447, w_eco90448, w_eco90449, w_eco90450, w_eco90451, w_eco90452, w_eco90453, w_eco90454, w_eco90455, w_eco90456, w_eco90457, w_eco90458, w_eco90459, w_eco90460, w_eco90461, w_eco90462, w_eco90463, w_eco90464, w_eco90465, w_eco90466, w_eco90467, w_eco90468, w_eco90469, w_eco90470, w_eco90471, w_eco90472, w_eco90473, w_eco90474, w_eco90475, w_eco90476, w_eco90477, w_eco90478, w_eco90479, w_eco90480, w_eco90481, w_eco90482, w_eco90483, w_eco90484, w_eco90485, w_eco90486, w_eco90487, w_eco90488, w_eco90489, w_eco90490, w_eco90491, w_eco90492, w_eco90493, w_eco90494, w_eco90495, w_eco90496, w_eco90497, w_eco90498, w_eco90499, w_eco90500, w_eco90501, w_eco90502, w_eco90503, w_eco90504, w_eco90505, w_eco90506, w_eco90507, w_eco90508, w_eco90509, w_eco90510, w_eco90511, w_eco90512, w_eco90513, w_eco90514, w_eco90515, w_eco90516, w_eco90517, w_eco90518, w_eco90519, w_eco90520, w_eco90521, w_eco90522, w_eco90523, w_eco90524, w_eco90525, w_eco90526, w_eco90527, w_eco90528, w_eco90529, w_eco90530, w_eco90531, w_eco90532, w_eco90533, w_eco90534, w_eco90535, w_eco90536, w_eco90537, w_eco90538, w_eco90539, w_eco90540, w_eco90541, w_eco90542, w_eco90543, w_eco90544, w_eco90545, w_eco90546, w_eco90547, w_eco90548, w_eco90549, w_eco90550, w_eco90551, w_eco90552, w_eco90553, w_eco90554, w_eco90555, w_eco90556, w_eco90557, w_eco90558, w_eco90559, w_eco90560, w_eco90561, w_eco90562, w_eco90563, w_eco90564, w_eco90565, w_eco90566, w_eco90567, w_eco90568, w_eco90569, w_eco90570, w_eco90571, w_eco90572, w_eco90573, w_eco90574, w_eco90575, w_eco90576, w_eco90577, w_eco90578, w_eco90579, w_eco90580, w_eco90581, w_eco90582, w_eco90583, w_eco90584, w_eco90585, w_eco90586, w_eco90587, w_eco90588, w_eco90589, w_eco90590, w_eco90591, w_eco90592, w_eco90593, w_eco90594, w_eco90595, w_eco90596, w_eco90597, w_eco90598, w_eco90599, w_eco90600, w_eco90601, w_eco90602, w_eco90603, w_eco90604, w_eco90605, w_eco90606, w_eco90607, w_eco90608, w_eco90609, w_eco90610, w_eco90611, w_eco90612, w_eco90613, w_eco90614, w_eco90615, w_eco90616, w_eco90617, w_eco90618, w_eco90619, w_eco90620, w_eco90621, w_eco90622, w_eco90623, w_eco90624, w_eco90625, w_eco90626, w_eco90627, w_eco90628, w_eco90629, w_eco90630, w_eco90631, w_eco90632, w_eco90633, w_eco90634, w_eco90635, w_eco90636, w_eco90637, w_eco90638, w_eco90639, w_eco90640, w_eco90641, w_eco90642, w_eco90643, w_eco90644, w_eco90645, w_eco90646, w_eco90647, w_eco90648, w_eco90649, w_eco90650, w_eco90651, w_eco90652, w_eco90653, w_eco90654, w_eco90655, w_eco90656, w_eco90657, w_eco90658, w_eco90659, w_eco90660, w_eco90661, w_eco90662, w_eco90663, w_eco90664, w_eco90665, w_eco90666, w_eco90667, w_eco90668, w_eco90669, w_eco90670, w_eco90671, w_eco90672, w_eco90673, w_eco90674, w_eco90675, w_eco90676, w_eco90677, w_eco90678, w_eco90679, w_eco90680, w_eco90681, w_eco90682, w_eco90683, w_eco90684, w_eco90685, w_eco90686, w_eco90687, w_eco90688, w_eco90689, w_eco90690, w_eco90691, w_eco90692, w_eco90693, w_eco90694, w_eco90695, w_eco90696, w_eco90697, w_eco90698, w_eco90699, w_eco90700, w_eco90701, w_eco90702, w_eco90703, w_eco90704, w_eco90705, w_eco90706, w_eco90707, w_eco90708, w_eco90709, w_eco90710, w_eco90711, w_eco90712, w_eco90713, w_eco90714, w_eco90715, w_eco90716, w_eco90717, w_eco90718, w_eco90719, w_eco90720, w_eco90721, w_eco90722, w_eco90723, w_eco90724, w_eco90725, w_eco90726, w_eco90727, w_eco90728, w_eco90729, w_eco90730, w_eco90731, w_eco90732, w_eco90733, w_eco90734, w_eco90735, w_eco90736, w_eco90737, w_eco90738, w_eco90739, w_eco90740, w_eco90741, w_eco90742, w_eco90743, w_eco90744, w_eco90745, w_eco90746, w_eco90747, w_eco90748, w_eco90749, w_eco90750, w_eco90751, w_eco90752, w_eco90753, w_eco90754, w_eco90755, w_eco90756, w_eco90757, w_eco90758, w_eco90759, w_eco90760, w_eco90761, w_eco90762, w_eco90763, w_eco90764, w_eco90765, w_eco90766, w_eco90767, w_eco90768, w_eco90769, w_eco90770, w_eco90771, w_eco90772, w_eco90773, w_eco90774, w_eco90775, w_eco90776, w_eco90777, w_eco90778, w_eco90779, w_eco90780, w_eco90781, w_eco90782, w_eco90783, w_eco90784, w_eco90785, w_eco90786, w_eco90787, w_eco90788, w_eco90789, w_eco90790, w_eco90791, w_eco90792, w_eco90793, w_eco90794, w_eco90795, w_eco90796, w_eco90797, w_eco90798, w_eco90799, w_eco90800, w_eco90801, w_eco90802, w_eco90803, w_eco90804, w_eco90805, w_eco90806, w_eco90807, w_eco90808, w_eco90809, w_eco90810, w_eco90811, w_eco90812, w_eco90813, w_eco90814, w_eco90815, w_eco90816, w_eco90817, w_eco90818, w_eco90819, w_eco90820, w_eco90821, w_eco90822, w_eco90823, w_eco90824, w_eco90825, w_eco90826, w_eco90827, w_eco90828, w_eco90829, w_eco90830, w_eco90831, w_eco90832, w_eco90833, w_eco90834, w_eco90835, w_eco90836, w_eco90837, w_eco90838, w_eco90839, w_eco90840, w_eco90841, w_eco90842, w_eco90843, w_eco90844, w_eco90845, w_eco90846, w_eco90847, w_eco90848, w_eco90849, w_eco90850, w_eco90851, w_eco90852, w_eco90853, w_eco90854, w_eco90855, w_eco90856, w_eco90857, w_eco90858, w_eco90859, w_eco90860, w_eco90861, w_eco90862, w_eco90863, w_eco90864, w_eco90865, w_eco90866, w_eco90867, w_eco90868, w_eco90869, w_eco90870, w_eco90871, w_eco90872, w_eco90873, w_eco90874, w_eco90875, w_eco90876, w_eco90877, w_eco90878, w_eco90879, w_eco90880, w_eco90881, w_eco90882, w_eco90883, w_eco90884, w_eco90885, w_eco90886, w_eco90887, w_eco90888, w_eco90889, w_eco90890, w_eco90891, w_eco90892, w_eco90893, w_eco90894, w_eco90895, w_eco90896, w_eco90897, w_eco90898, w_eco90899, w_eco90900, w_eco90901, w_eco90902, w_eco90903, w_eco90904, w_eco90905, w_eco90906, w_eco90907, w_eco90908, w_eco90909, w_eco90910, w_eco90911, w_eco90912, w_eco90913, w_eco90914, w_eco90915, w_eco90916, w_eco90917, w_eco90918, w_eco90919, w_eco90920, w_eco90921, w_eco90922, w_eco90923, w_eco90924, w_eco90925, w_eco90926, w_eco90927, w_eco90928, w_eco90929, w_eco90930, w_eco90931, w_eco90932, w_eco90933, w_eco90934, w_eco90935, w_eco90936, w_eco90937, w_eco90938, w_eco90939, w_eco90940, w_eco90941, w_eco90942, w_eco90943, w_eco90944, w_eco90945, w_eco90946, w_eco90947, w_eco90948, w_eco90949, w_eco90950, w_eco90951, w_eco90952, w_eco90953, w_eco90954, w_eco90955, w_eco90956, w_eco90957, w_eco90958, w_eco90959, w_eco90960, w_eco90961, w_eco90962, w_eco90963, w_eco90964, w_eco90965, w_eco90966, w_eco90967, w_eco90968, w_eco90969, w_eco90970, w_eco90971, w_eco90972, w_eco90973, w_eco90974, w_eco90975, w_eco90976, w_eco90977, w_eco90978, w_eco90979, w_eco90980, w_eco90981, w_eco90982, w_eco90983, w_eco90984, w_eco90985, w_eco90986, w_eco90987, w_eco90988, w_eco90989, w_eco90990, w_eco90991, w_eco90992, w_eco90993, w_eco90994, w_eco90995, w_eco90996, w_eco90997, w_eco90998, w_eco90999, w_eco91000, w_eco91001, w_eco91002, w_eco91003, w_eco91004, w_eco91005, w_eco91006, w_eco91007, w_eco91008, w_eco91009, w_eco91010, w_eco91011, w_eco91012, w_eco91013, w_eco91014, w_eco91015, w_eco91016, w_eco91017, w_eco91018, w_eco91019, w_eco91020, w_eco91021, w_eco91022, w_eco91023, w_eco91024, w_eco91025, w_eco91026, w_eco91027, w_eco91028, w_eco91029, w_eco91030, w_eco91031, w_eco91032, w_eco91033, w_eco91034, w_eco91035, w_eco91036, w_eco91037, w_eco91038, w_eco91039, w_eco91040, w_eco91041, w_eco91042, w_eco91043, w_eco91044, w_eco91045, w_eco91046, w_eco91047, w_eco91048, w_eco91049, w_eco91050, w_eco91051, w_eco91052, w_eco91053, w_eco91054, w_eco91055, w_eco91056, w_eco91057, w_eco91058, w_eco91059, w_eco91060, w_eco91061, w_eco91062, w_eco91063, w_eco91064, w_eco91065, w_eco91066, w_eco91067, w_eco91068, w_eco91069, w_eco91070, w_eco91071, w_eco91072, w_eco91073, w_eco91074, w_eco91075, w_eco91076, w_eco91077, w_eco91078, w_eco91079, w_eco91080, w_eco91081, w_eco91082, w_eco91083, w_eco91084, w_eco91085, w_eco91086, w_eco91087, w_eco91088, w_eco91089, w_eco91090, w_eco91091, w_eco91092, w_eco91093, w_eco91094, w_eco91095, w_eco91096, w_eco91097, w_eco91098, w_eco91099, w_eco91100, w_eco91101, w_eco91102, w_eco91103, w_eco91104, w_eco91105, w_eco91106, w_eco91107, w_eco91108, w_eco91109, w_eco91110, w_eco91111, w_eco91112, w_eco91113, w_eco91114, w_eco91115, w_eco91116, w_eco91117, w_eco91118, w_eco91119, w_eco91120, w_eco91121, w_eco91122, w_eco91123, w_eco91124, w_eco91125, w_eco91126, w_eco91127, w_eco91128, w_eco91129, w_eco91130, w_eco91131, w_eco91132, w_eco91133, w_eco91134, w_eco91135, w_eco91136, w_eco91137, w_eco91138, w_eco91139, w_eco91140, w_eco91141, w_eco91142, w_eco91143, w_eco91144, w_eco91145, w_eco91146, w_eco91147, w_eco91148, w_eco91149, w_eco91150, w_eco91151, w_eco91152, w_eco91153, w_eco91154, w_eco91155, w_eco91156, w_eco91157, w_eco91158, w_eco91159, w_eco91160, w_eco91161, w_eco91162, w_eco91163, w_eco91164, w_eco91165, w_eco91166, w_eco91167, w_eco91168, w_eco91169, w_eco91170, w_eco91171, w_eco91172, w_eco91173, w_eco91174, w_eco91175, w_eco91176, w_eco91177, w_eco91178, w_eco91179, w_eco91180, w_eco91181, w_eco91182, w_eco91183, w_eco91184, w_eco91185, w_eco91186, w_eco91187, w_eco91188, w_eco91189, w_eco91190, w_eco91191, w_eco91192, w_eco91193, w_eco91194, w_eco91195, w_eco91196, w_eco91197, w_eco91198, w_eco91199, w_eco91200, w_eco91201, w_eco91202, w_eco91203, w_eco91204, w_eco91205, w_eco91206, w_eco91207, w_eco91208, w_eco91209, w_eco91210, w_eco91211, w_eco91212, w_eco91213, w_eco91214, w_eco91215, w_eco91216, w_eco91217, w_eco91218, w_eco91219, w_eco91220, w_eco91221, w_eco91222, w_eco91223, w_eco91224, w_eco91225, w_eco91226, w_eco91227, w_eco91228, w_eco91229, w_eco91230, w_eco91231, w_eco91232, w_eco91233, w_eco91234, w_eco91235, w_eco91236, w_eco91237, w_eco91238, w_eco91239, w_eco91240, w_eco91241, w_eco91242, w_eco91243, w_eco91244, w_eco91245, w_eco91246, w_eco91247, w_eco91248, w_eco91249, w_eco91250, w_eco91251, w_eco91252, w_eco91253, w_eco91254, w_eco91255, w_eco91256, w_eco91257, w_eco91258, w_eco91259, w_eco91260, w_eco91261, w_eco91262, w_eco91263, w_eco91264, w_eco91265, w_eco91266, w_eco91267, w_eco91268, w_eco91269, w_eco91270, w_eco91271, w_eco91272, w_eco91273, w_eco91274, w_eco91275, w_eco91276, w_eco91277, w_eco91278, w_eco91279, w_eco91280, w_eco91281, w_eco91282, w_eco91283, w_eco91284, w_eco91285, w_eco91286, w_eco91287, w_eco91288, w_eco91289, w_eco91290, w_eco91291, w_eco91292, w_eco91293, w_eco91294, w_eco91295, w_eco91296, w_eco91297, w_eco91298, w_eco91299, w_eco91300, w_eco91301, w_eco91302, w_eco91303, w_eco91304, w_eco91305, w_eco91306, w_eco91307, w_eco91308, w_eco91309, w_eco91310, w_eco91311, w_eco91312, w_eco91313, w_eco91314, w_eco91315, w_eco91316, w_eco91317, w_eco91318, w_eco91319, w_eco91320, w_eco91321, w_eco91322, w_eco91323, w_eco91324, w_eco91325, w_eco91326, w_eco91327, w_eco91328, w_eco91329, w_eco91330, w_eco91331, w_eco91332, w_eco91333, w_eco91334, w_eco91335, w_eco91336, w_eco91337, w_eco91338, w_eco91339, w_eco91340, w_eco91341, w_eco91342, w_eco91343, w_eco91344, w_eco91345, w_eco91346, w_eco91347, w_eco91348, w_eco91349, w_eco91350, w_eco91351, w_eco91352, w_eco91353, w_eco91354, w_eco91355, w_eco91356, w_eco91357, w_eco91358, w_eco91359, w_eco91360, w_eco91361, w_eco91362, w_eco91363, w_eco91364, w_eco91365, w_eco91366, w_eco91367, w_eco91368, w_eco91369, w_eco91370, w_eco91371, w_eco91372, w_eco91373, w_eco91374, w_eco91375, w_eco91376, w_eco91377, w_eco91378, w_eco91379, w_eco91380, w_eco91381, w_eco91382, w_eco91383, w_eco91384, w_eco91385, w_eco91386, w_eco91387, w_eco91388, w_eco91389, w_eco91390, w_eco91391, w_eco91392, w_eco91393, w_eco91394, w_eco91395, w_eco91396, w_eco91397, w_eco91398, w_eco91399, w_eco91400, w_eco91401, w_eco91402, w_eco91403, w_eco91404, w_eco91405, w_eco91406, w_eco91407, w_eco91408, w_eco91409, w_eco91410, w_eco91411, w_eco91412, w_eco91413, w_eco91414, w_eco91415, w_eco91416, w_eco91417, w_eco91418, w_eco91419, w_eco91420, w_eco91421, w_eco91422, w_eco91423, w_eco91424, w_eco91425, w_eco91426, w_eco91427, w_eco91428, w_eco91429, w_eco91430, w_eco91431, w_eco91432, w_eco91433, w_eco91434, w_eco91435, w_eco91436, w_eco91437, w_eco91438, w_eco91439, w_eco91440, w_eco91441, w_eco91442, w_eco91443, w_eco91444, w_eco91445, w_eco91446, w_eco91447, w_eco91448, w_eco91449, w_eco91450, w_eco91451, w_eco91452, w_eco91453, w_eco91454, w_eco91455, w_eco91456, w_eco91457, w_eco91458, w_eco91459, w_eco91460, w_eco91461, w_eco91462, w_eco91463, w_eco91464, w_eco91465, w_eco91466, w_eco91467, w_eco91468, w_eco91469, w_eco91470, w_eco91471, w_eco91472, w_eco91473, w_eco91474, w_eco91475, w_eco91476, w_eco91477, w_eco91478, w_eco91479, w_eco91480, w_eco91481, w_eco91482, w_eco91483, w_eco91484, w_eco91485, w_eco91486, w_eco91487, w_eco91488, w_eco91489, w_eco91490, w_eco91491, w_eco91492, w_eco91493, w_eco91494, w_eco91495, w_eco91496, w_eco91497, w_eco91498, w_eco91499, w_eco91500, w_eco91501, w_eco91502, w_eco91503, w_eco91504, w_eco91505, w_eco91506, w_eco91507, w_eco91508, w_eco91509, w_eco91510, w_eco91511, w_eco91512, w_eco91513, w_eco91514, w_eco91515, w_eco91516, w_eco91517, w_eco91518, w_eco91519, w_eco91520, w_eco91521, w_eco91522, w_eco91523, w_eco91524, w_eco91525, w_eco91526, w_eco91527, w_eco91528, w_eco91529, w_eco91530, w_eco91531, w_eco91532, w_eco91533, w_eco91534, w_eco91535, w_eco91536, w_eco91537, w_eco91538, w_eco91539, w_eco91540, w_eco91541, w_eco91542, w_eco91543, w_eco91544, w_eco91545, w_eco91546, w_eco91547, w_eco91548, w_eco91549, w_eco91550, w_eco91551, w_eco91552, w_eco91553, w_eco91554, w_eco91555, w_eco91556, w_eco91557, w_eco91558, w_eco91559, w_eco91560, w_eco91561, w_eco91562, w_eco91563, w_eco91564, w_eco91565, w_eco91566, w_eco91567, w_eco91568, w_eco91569, w_eco91570, w_eco91571, w_eco91572, w_eco91573, w_eco91574, w_eco91575, w_eco91576, w_eco91577, w_eco91578, w_eco91579, w_eco91580, w_eco91581, w_eco91582, w_eco91583, w_eco91584, w_eco91585, w_eco91586, w_eco91587, w_eco91588, w_eco91589, w_eco91590, w_eco91591, w_eco91592, w_eco91593, w_eco91594, w_eco91595, w_eco91596, w_eco91597, w_eco91598, w_eco91599, w_eco91600, w_eco91601, w_eco91602, w_eco91603, w_eco91604, w_eco91605, w_eco91606, w_eco91607, w_eco91608, w_eco91609, w_eco91610, w_eco91611, w_eco91612, w_eco91613, w_eco91614, w_eco91615, w_eco91616, w_eco91617, w_eco91618, w_eco91619, w_eco91620, w_eco91621, w_eco91622, w_eco91623, w_eco91624, w_eco91625, w_eco91626, w_eco91627, w_eco91628, w_eco91629, w_eco91630, w_eco91631, w_eco91632, w_eco91633, w_eco91634, w_eco91635, w_eco91636, w_eco91637, w_eco91638, w_eco91639, w_eco91640, w_eco91641, w_eco91642, w_eco91643, w_eco91644, w_eco91645, w_eco91646, w_eco91647, w_eco91648, w_eco91649, w_eco91650, w_eco91651, w_eco91652, w_eco91653, w_eco91654, w_eco91655, w_eco91656, w_eco91657, w_eco91658, w_eco91659, w_eco91660, w_eco91661, w_eco91662, w_eco91663, w_eco91664, w_eco91665, w_eco91666, w_eco91667, w_eco91668, w_eco91669, w_eco91670, w_eco91671, w_eco91672, w_eco91673, w_eco91674, w_eco91675, w_eco91676, w_eco91677, w_eco91678, w_eco91679, w_eco91680, w_eco91681, w_eco91682, w_eco91683, w_eco91684, w_eco91685, w_eco91686, w_eco91687, w_eco91688, w_eco91689, w_eco91690, w_eco91691, w_eco91692, w_eco91693, w_eco91694, w_eco91695, w_eco91696, w_eco91697, w_eco91698, w_eco91699, w_eco91700, w_eco91701, w_eco91702, w_eco91703, w_eco91704, w_eco91705, w_eco91706, w_eco91707, w_eco91708, w_eco91709, w_eco91710, w_eco91711, w_eco91712, w_eco91713, w_eco91714, w_eco91715, w_eco91716, w_eco91717, w_eco91718, w_eco91719, w_eco91720, w_eco91721, w_eco91722, w_eco91723, w_eco91724, w_eco91725, w_eco91726, w_eco91727, w_eco91728, w_eco91729, w_eco91730, w_eco91731, w_eco91732, w_eco91733, w_eco91734, w_eco91735, w_eco91736, w_eco91737, w_eco91738, w_eco91739, w_eco91740, w_eco91741, w_eco91742, w_eco91743, w_eco91744, w_eco91745, w_eco91746, w_eco91747, w_eco91748, w_eco91749, w_eco91750, w_eco91751, w_eco91752, w_eco91753, w_eco91754, w_eco91755, w_eco91756, w_eco91757, w_eco91758, w_eco91759, w_eco91760, w_eco91761, w_eco91762, w_eco91763, w_eco91764, w_eco91765, w_eco91766, w_eco91767, w_eco91768, w_eco91769, w_eco91770, w_eco91771, w_eco91772, w_eco91773, w_eco91774, w_eco91775, w_eco91776, w_eco91777, w_eco91778, w_eco91779, w_eco91780, w_eco91781, w_eco91782, w_eco91783, w_eco91784, w_eco91785, w_eco91786, w_eco91787, w_eco91788, w_eco91789, w_eco91790, w_eco91791, w_eco91792, w_eco91793, w_eco91794, w_eco91795, w_eco91796, w_eco91797, w_eco91798, w_eco91799, w_eco91800, w_eco91801, w_eco91802, w_eco91803, w_eco91804, w_eco91805, w_eco91806, w_eco91807, w_eco91808, w_eco91809, w_eco91810, w_eco91811, w_eco91812, w_eco91813, w_eco91814, w_eco91815, w_eco91816, w_eco91817, w_eco91818, w_eco91819, w_eco91820, w_eco91821, w_eco91822, w_eco91823, w_eco91824, w_eco91825, w_eco91826, w_eco91827, w_eco91828, w_eco91829, w_eco91830, w_eco91831, w_eco91832, w_eco91833, w_eco91834, w_eco91835, w_eco91836, w_eco91837, w_eco91838, w_eco91839, w_eco91840, w_eco91841, w_eco91842, w_eco91843, w_eco91844, w_eco91845, w_eco91846, w_eco91847, w_eco91848, w_eco91849, w_eco91850, w_eco91851, w_eco91852, w_eco91853, w_eco91854, w_eco91855, w_eco91856, w_eco91857, w_eco91858, w_eco91859, w_eco91860, w_eco91861, w_eco91862, w_eco91863, w_eco91864, w_eco91865, w_eco91866, w_eco91867, w_eco91868, w_eco91869, w_eco91870, w_eco91871, w_eco91872, w_eco91873, w_eco91874, w_eco91875, w_eco91876, w_eco91877, w_eco91878, w_eco91879, w_eco91880, w_eco91881, w_eco91882, w_eco91883, w_eco91884, w_eco91885, w_eco91886, w_eco91887, w_eco91888, w_eco91889, w_eco91890, w_eco91891, w_eco91892, w_eco91893, w_eco91894, w_eco91895, w_eco91896, w_eco91897, w_eco91898, w_eco91899, w_eco91900, w_eco91901, w_eco91902, w_eco91903, w_eco91904, w_eco91905, w_eco91906, w_eco91907, w_eco91908, w_eco91909, w_eco91910, w_eco91911, w_eco91912, w_eco91913, w_eco91914, w_eco91915, w_eco91916, w_eco91917, w_eco91918, w_eco91919, w_eco91920, w_eco91921, w_eco91922, w_eco91923, w_eco91924, w_eco91925, w_eco91926, w_eco91927, w_eco91928, w_eco91929, w_eco91930, w_eco91931, w_eco91932, w_eco91933, w_eco91934, w_eco91935, w_eco91936, w_eco91937, w_eco91938, w_eco91939, w_eco91940, w_eco91941, w_eco91942, w_eco91943, w_eco91944, w_eco91945, w_eco91946, w_eco91947, w_eco91948, w_eco91949, w_eco91950, w_eco91951, w_eco91952, w_eco91953, w_eco91954, w_eco91955, w_eco91956, w_eco91957, w_eco91958, w_eco91959, w_eco91960, w_eco91961, w_eco91962, w_eco91963, w_eco91964, w_eco91965, w_eco91966, w_eco91967, w_eco91968, w_eco91969, w_eco91970, w_eco91971, w_eco91972, w_eco91973, w_eco91974, w_eco91975, w_eco91976, w_eco91977, w_eco91978, w_eco91979, w_eco91980, w_eco91981, w_eco91982, w_eco91983, w_eco91984, w_eco91985, w_eco91986, w_eco91987, w_eco91988, w_eco91989, w_eco91990, w_eco91991, w_eco91992, w_eco91993, w_eco91994, w_eco91995, w_eco91996, w_eco91997, w_eco91998, w_eco91999, w_eco92000, w_eco92001, w_eco92002, w_eco92003, w_eco92004, w_eco92005, w_eco92006, w_eco92007, w_eco92008, w_eco92009, w_eco92010, w_eco92011, w_eco92012, w_eco92013, w_eco92014, w_eco92015, w_eco92016, w_eco92017, w_eco92018, w_eco92019, w_eco92020, w_eco92021, w_eco92022, w_eco92023, w_eco92024, w_eco92025, w_eco92026, w_eco92027, w_eco92028, w_eco92029, w_eco92030, w_eco92031, w_eco92032, w_eco92033, w_eco92034, w_eco92035, w_eco92036, w_eco92037, w_eco92038, w_eco92039, w_eco92040, w_eco92041, w_eco92042, w_eco92043, w_eco92044, w_eco92045, w_eco92046, w_eco92047, w_eco92048, w_eco92049, w_eco92050, w_eco92051, w_eco92052, w_eco92053, w_eco92054, w_eco92055, w_eco92056, w_eco92057, w_eco92058, w_eco92059, w_eco92060, w_eco92061, w_eco92062, w_eco92063, w_eco92064, w_eco92065, w_eco92066, w_eco92067, w_eco92068, w_eco92069, w_eco92070, w_eco92071, w_eco92072, w_eco92073, w_eco92074, w_eco92075, w_eco92076, w_eco92077, w_eco92078, w_eco92079, w_eco92080, w_eco92081, w_eco92082, w_eco92083, w_eco92084, w_eco92085, w_eco92086, w_eco92087, w_eco92088, w_eco92089, w_eco92090, w_eco92091, w_eco92092, w_eco92093, w_eco92094, w_eco92095, w_eco92096, w_eco92097, w_eco92098, w_eco92099, w_eco92100, w_eco92101, w_eco92102, w_eco92103, w_eco92104, w_eco92105, w_eco92106, w_eco92107, w_eco92108, w_eco92109, w_eco92110, w_eco92111, w_eco92112, w_eco92113, w_eco92114, w_eco92115, w_eco92116, w_eco92117, w_eco92118, w_eco92119, w_eco92120, w_eco92121, w_eco92122, w_eco92123, w_eco92124, w_eco92125, w_eco92126, w_eco92127, w_eco92128, w_eco92129, w_eco92130, w_eco92131, w_eco92132, w_eco92133, w_eco92134, w_eco92135, w_eco92136, w_eco92137, w_eco92138, w_eco92139, w_eco92140, w_eco92141, w_eco92142, w_eco92143, w_eco92144, w_eco92145, w_eco92146, w_eco92147, w_eco92148, w_eco92149, w_eco92150, w_eco92151, w_eco92152, w_eco92153, w_eco92154, w_eco92155, w_eco92156, w_eco92157, w_eco92158, w_eco92159, w_eco92160, w_eco92161, w_eco92162, w_eco92163, w_eco92164, w_eco92165, w_eco92166, w_eco92167, w_eco92168, w_eco92169, w_eco92170, w_eco92171, w_eco92172, w_eco92173, w_eco92174, w_eco92175, w_eco92176, w_eco92177, w_eco92178, w_eco92179, w_eco92180, w_eco92181, w_eco92182, w_eco92183, w_eco92184, w_eco92185, w_eco92186, w_eco92187, w_eco92188, w_eco92189, w_eco92190, w_eco92191, w_eco92192, w_eco92193, w_eco92194, w_eco92195, w_eco92196, w_eco92197, w_eco92198, w_eco92199, w_eco92200, w_eco92201, w_eco92202, w_eco92203, w_eco92204, w_eco92205, w_eco92206, w_eco92207, w_eco92208, w_eco92209, w_eco92210, w_eco92211, w_eco92212, w_eco92213, w_eco92214, w_eco92215, w_eco92216, w_eco92217, w_eco92218, w_eco92219, w_eco92220, w_eco92221, w_eco92222, w_eco92223, w_eco92224, w_eco92225, w_eco92226, w_eco92227, w_eco92228, w_eco92229, w_eco92230, w_eco92231, w_eco92232, w_eco92233, w_eco92234, w_eco92235, w_eco92236, w_eco92237, w_eco92238, w_eco92239, w_eco92240, w_eco92241, w_eco92242, w_eco92243, w_eco92244, w_eco92245, w_eco92246, w_eco92247, w_eco92248, w_eco92249, w_eco92250, w_eco92251, w_eco92252, w_eco92253, w_eco92254, w_eco92255, w_eco92256, w_eco92257, w_eco92258, w_eco92259, w_eco92260, w_eco92261, w_eco92262, w_eco92263, w_eco92264, w_eco92265, w_eco92266, w_eco92267, w_eco92268, w_eco92269, w_eco92270, w_eco92271, w_eco92272, w_eco92273, w_eco92274, w_eco92275, w_eco92276, w_eco92277, w_eco92278, w_eco92279, w_eco92280, w_eco92281, w_eco92282, w_eco92283, w_eco92284, w_eco92285, w_eco92286, w_eco92287, w_eco92288, w_eco92289, w_eco92290, w_eco92291, w_eco92292, w_eco92293, w_eco92294, w_eco92295, w_eco92296, w_eco92297, w_eco92298, w_eco92299, w_eco92300, w_eco92301, w_eco92302, w_eco92303, w_eco92304, w_eco92305, w_eco92306, w_eco92307, w_eco92308, w_eco92309, w_eco92310, w_eco92311, w_eco92312, w_eco92313, w_eco92314, w_eco92315, w_eco92316, w_eco92317, w_eco92318, w_eco92319, w_eco92320, w_eco92321, w_eco92322, w_eco92323, w_eco92324, w_eco92325, w_eco92326, w_eco92327, w_eco92328, w_eco92329, w_eco92330, w_eco92331, w_eco92332, w_eco92333, w_eco92334, w_eco92335, w_eco92336, w_eco92337, w_eco92338, w_eco92339, w_eco92340, w_eco92341, w_eco92342, w_eco92343, w_eco92344, w_eco92345, w_eco92346, w_eco92347, w_eco92348, w_eco92349, w_eco92350, w_eco92351, w_eco92352, w_eco92353, w_eco92354, w_eco92355, w_eco92356, w_eco92357, w_eco92358, w_eco92359, w_eco92360, w_eco92361, w_eco92362, w_eco92363, w_eco92364, w_eco92365, w_eco92366, w_eco92367, w_eco92368, w_eco92369, w_eco92370, w_eco92371, w_eco92372, w_eco92373, w_eco92374, w_eco92375, w_eco92376, w_eco92377, w_eco92378, w_eco92379, w_eco92380, w_eco92381, w_eco92382, w_eco92383, w_eco92384, w_eco92385, w_eco92386, w_eco92387, w_eco92388, w_eco92389, w_eco92390, w_eco92391, w_eco92392, w_eco92393, w_eco92394, w_eco92395, w_eco92396, w_eco92397, w_eco92398, w_eco92399, w_eco92400, w_eco92401, w_eco92402, w_eco92403, w_eco92404, w_eco92405, w_eco92406, w_eco92407, w_eco92408, w_eco92409, w_eco92410, w_eco92411, w_eco92412, w_eco92413, w_eco92414, w_eco92415, w_eco92416, w_eco92417, w_eco92418, w_eco92419, w_eco92420, w_eco92421, w_eco92422, w_eco92423, w_eco92424, w_eco92425, w_eco92426, w_eco92427, w_eco92428, w_eco92429, w_eco92430, w_eco92431, w_eco92432, w_eco92433, w_eco92434, w_eco92435, w_eco92436, w_eco92437, w_eco92438, w_eco92439, w_eco92440, w_eco92441, w_eco92442, w_eco92443, w_eco92444, w_eco92445, w_eco92446, w_eco92447, w_eco92448, w_eco92449, w_eco92450, w_eco92451, w_eco92452, w_eco92453, w_eco92454, w_eco92455, w_eco92456, w_eco92457, w_eco92458, w_eco92459, w_eco92460, w_eco92461, w_eco92462, w_eco92463, w_eco92464, w_eco92465, w_eco92466, w_eco92467, w_eco92468, w_eco92469, w_eco92470, w_eco92471, w_eco92472, w_eco92473, w_eco92474, w_eco92475, w_eco92476, w_eco92477, w_eco92478, w_eco92479, w_eco92480, w_eco92481, w_eco92482, w_eco92483, w_eco92484, w_eco92485, w_eco92486, w_eco92487, w_eco92488, w_eco92489, w_eco92490, w_eco92491, w_eco92492, w_eco92493, w_eco92494, w_eco92495, w_eco92496, w_eco92497, w_eco92498, w_eco92499, w_eco92500, w_eco92501, w_eco92502, w_eco92503, w_eco92504, w_eco92505, w_eco92506, w_eco92507, w_eco92508, w_eco92509, w_eco92510, w_eco92511, w_eco92512, w_eco92513, w_eco92514, w_eco92515, w_eco92516, w_eco92517, w_eco92518, w_eco92519, w_eco92520, w_eco92521, w_eco92522, w_eco92523, w_eco92524, w_eco92525, w_eco92526, w_eco92527, w_eco92528, w_eco92529, w_eco92530, w_eco92531, w_eco92532, w_eco92533, w_eco92534, w_eco92535, w_eco92536, w_eco92537, w_eco92538, w_eco92539, w_eco92540, w_eco92541, w_eco92542, w_eco92543, w_eco92544, w_eco92545, w_eco92546, w_eco92547, w_eco92548, w_eco92549, w_eco92550, w_eco92551, w_eco92552, w_eco92553, w_eco92554, w_eco92555, w_eco92556, w_eco92557, w_eco92558, w_eco92559, w_eco92560, w_eco92561, w_eco92562, w_eco92563, w_eco92564, w_eco92565, w_eco92566, w_eco92567, w_eco92568, w_eco92569, w_eco92570, w_eco92571, w_eco92572, w_eco92573, w_eco92574, w_eco92575, w_eco92576, w_eco92577, w_eco92578, w_eco92579, w_eco92580, w_eco92581, w_eco92582, w_eco92583, w_eco92584, w_eco92585, w_eco92586, w_eco92587, w_eco92588, w_eco92589, w_eco92590, w_eco92591, w_eco92592, w_eco92593, w_eco92594, w_eco92595, w_eco92596, w_eco92597, w_eco92598, w_eco92599, w_eco92600, w_eco92601, w_eco92602, w_eco92603, w_eco92604, w_eco92605, w_eco92606, w_eco92607, w_eco92608, w_eco92609, w_eco92610, w_eco92611, w_eco92612, w_eco92613, w_eco92614, w_eco92615, w_eco92616, w_eco92617, w_eco92618, w_eco92619, w_eco92620, w_eco92621, w_eco92622, w_eco92623, w_eco92624, w_eco92625, w_eco92626, w_eco92627, w_eco92628, w_eco92629, w_eco92630, w_eco92631, w_eco92632, w_eco92633, w_eco92634, w_eco92635, w_eco92636, w_eco92637, w_eco92638, w_eco92639, w_eco92640, w_eco92641, w_eco92642, w_eco92643, w_eco92644, w_eco92645, w_eco92646, w_eco92647, w_eco92648, w_eco92649, w_eco92650, w_eco92651, w_eco92652, w_eco92653, w_eco92654, w_eco92655, w_eco92656, w_eco92657, w_eco92658, w_eco92659, w_eco92660, w_eco92661, w_eco92662, w_eco92663, w_eco92664, w_eco92665, w_eco92666, w_eco92667, w_eco92668, w_eco92669, w_eco92670, w_eco92671, w_eco92672, w_eco92673, w_eco92674, w_eco92675, w_eco92676, w_eco92677, w_eco92678, w_eco92679, w_eco92680, w_eco92681, w_eco92682, w_eco92683, w_eco92684, w_eco92685, w_eco92686, w_eco92687, w_eco92688, w_eco92689, w_eco92690, w_eco92691, w_eco92692, w_eco92693, w_eco92694, w_eco92695, w_eco92696, w_eco92697, w_eco92698, w_eco92699, w_eco92700, w_eco92701, w_eco92702, w_eco92703, w_eco92704, w_eco92705, w_eco92706, w_eco92707, w_eco92708, w_eco92709, w_eco92710, w_eco92711, w_eco92712, w_eco92713, w_eco92714, w_eco92715, w_eco92716, w_eco92717, w_eco92718, w_eco92719, w_eco92720, w_eco92721, w_eco92722, w_eco92723, w_eco92724, w_eco92725, w_eco92726, w_eco92727, w_eco92728, w_eco92729, w_eco92730, w_eco92731, w_eco92732, w_eco92733, w_eco92734, w_eco92735, w_eco92736, w_eco92737, w_eco92738, w_eco92739, w_eco92740, w_eco92741, w_eco92742, w_eco92743, w_eco92744, w_eco92745, w_eco92746, w_eco92747, w_eco92748, w_eco92749, w_eco92750, w_eco92751, w_eco92752, w_eco92753, w_eco92754, w_eco92755, w_eco92756, w_eco92757, w_eco92758, w_eco92759, w_eco92760, w_eco92761, w_eco92762, w_eco92763, w_eco92764, w_eco92765, w_eco92766, w_eco92767, w_eco92768, w_eco92769, w_eco92770, w_eco92771, w_eco92772, w_eco92773, w_eco92774, w_eco92775, w_eco92776, w_eco92777, w_eco92778, w_eco92779, w_eco92780, w_eco92781, w_eco92782, w_eco92783, w_eco92784, w_eco92785, w_eco92786, w_eco92787, w_eco92788, w_eco92789, w_eco92790, w_eco92791, w_eco92792, w_eco92793, w_eco92794, w_eco92795, w_eco92796, w_eco92797, w_eco92798, w_eco92799, w_eco92800, w_eco92801, w_eco92802, w_eco92803, w_eco92804, w_eco92805, w_eco92806, w_eco92807, w_eco92808, w_eco92809, w_eco92810, w_eco92811, w_eco92812, w_eco92813, w_eco92814, w_eco92815, w_eco92816, w_eco92817, w_eco92818, w_eco92819, w_eco92820, w_eco92821, w_eco92822, w_eco92823, w_eco92824, w_eco92825, w_eco92826, w_eco92827, w_eco92828, w_eco92829, w_eco92830, w_eco92831, w_eco92832, w_eco92833, w_eco92834, w_eco92835, w_eco92836, w_eco92837, w_eco92838, w_eco92839, w_eco92840, w_eco92841, w_eco92842, w_eco92843, w_eco92844, w_eco92845, w_eco92846, w_eco92847, w_eco92848, w_eco92849, w_eco92850, w_eco92851, w_eco92852, w_eco92853, w_eco92854, w_eco92855, w_eco92856, w_eco92857, w_eco92858, w_eco92859, w_eco92860, w_eco92861, w_eco92862, w_eco92863, w_eco92864, w_eco92865, w_eco92866, w_eco92867, w_eco92868, w_eco92869, w_eco92870, w_eco92871, w_eco92872, w_eco92873, w_eco92874, w_eco92875, w_eco92876, w_eco92877, w_eco92878, w_eco92879, w_eco92880, w_eco92881, w_eco92882, w_eco92883, w_eco92884, w_eco92885, w_eco92886, w_eco92887, w_eco92888, w_eco92889, w_eco92890, w_eco92891, w_eco92892, w_eco92893, w_eco92894, w_eco92895, w_eco92896, w_eco92897, w_eco92898, w_eco92899, w_eco92900, w_eco92901, w_eco92902, w_eco92903, w_eco92904, w_eco92905, w_eco92906, w_eco92907, w_eco92908, w_eco92909, w_eco92910, w_eco92911, w_eco92912, w_eco92913, w_eco92914, w_eco92915, w_eco92916, w_eco92917, w_eco92918, w_eco92919, w_eco92920, w_eco92921, w_eco92922, w_eco92923, w_eco92924, w_eco92925, w_eco92926, w_eco92927, w_eco92928, w_eco92929, w_eco92930, w_eco92931, w_eco92932, w_eco92933, w_eco92934, w_eco92935, w_eco92936, w_eco92937, w_eco92938, w_eco92939, w_eco92940, w_eco92941, w_eco92942, w_eco92943, w_eco92944, w_eco92945, w_eco92946, w_eco92947, w_eco92948, w_eco92949, w_eco92950, w_eco92951, w_eco92952, w_eco92953, w_eco92954, w_eco92955, w_eco92956, w_eco92957, w_eco92958, w_eco92959, w_eco92960, w_eco92961, w_eco92962, w_eco92963, w_eco92964, w_eco92965, w_eco92966, w_eco92967, w_eco92968, w_eco92969, w_eco92970, w_eco92971, w_eco92972, w_eco92973, w_eco92974, w_eco92975, w_eco92976, w_eco92977, w_eco92978, w_eco92979, w_eco92980, w_eco92981, w_eco92982, w_eco92983, w_eco92984, w_eco92985, w_eco92986, w_eco92987, w_eco92988, w_eco92989, w_eco92990, w_eco92991, w_eco92992, w_eco92993, w_eco92994, w_eco92995, w_eco92996, w_eco92997, w_eco92998, w_eco92999, w_eco93000, w_eco93001, w_eco93002, w_eco93003, w_eco93004, w_eco93005, w_eco93006, w_eco93007, w_eco93008, w_eco93009, w_eco93010, w_eco93011, w_eco93012, w_eco93013, w_eco93014, w_eco93015, w_eco93016, w_eco93017, w_eco93018, w_eco93019, w_eco93020, w_eco93021, w_eco93022, w_eco93023, w_eco93024, w_eco93025, w_eco93026, w_eco93027, w_eco93028, w_eco93029, w_eco93030, w_eco93031, w_eco93032, w_eco93033, w_eco93034, w_eco93035, w_eco93036, w_eco93037, w_eco93038, w_eco93039, w_eco93040, w_eco93041, w_eco93042, w_eco93043, w_eco93044, w_eco93045, w_eco93046, w_eco93047, w_eco93048, w_eco93049, w_eco93050, w_eco93051, w_eco93052, w_eco93053, w_eco93054, w_eco93055, w_eco93056, w_eco93057, w_eco93058, w_eco93059, w_eco93060, w_eco93061, w_eco93062, w_eco93063, w_eco93064, w_eco93065, w_eco93066, w_eco93067, w_eco93068, w_eco93069, w_eco93070, w_eco93071, w_eco93072, w_eco93073, w_eco93074, w_eco93075, w_eco93076, w_eco93077, w_eco93078, w_eco93079, w_eco93080, w_eco93081, w_eco93082, w_eco93083, w_eco93084, w_eco93085, w_eco93086, w_eco93087, w_eco93088, w_eco93089, w_eco93090, w_eco93091, w_eco93092, w_eco93093, w_eco93094, w_eco93095, w_eco93096, w_eco93097, w_eco93098, w_eco93099, w_eco93100, w_eco93101, w_eco93102, w_eco93103, w_eco93104, w_eco93105, w_eco93106, w_eco93107, w_eco93108, w_eco93109, w_eco93110, w_eco93111, w_eco93112, w_eco93113, w_eco93114, w_eco93115, w_eco93116, w_eco93117, w_eco93118, w_eco93119, w_eco93120, w_eco93121, w_eco93122, w_eco93123, w_eco93124, w_eco93125, w_eco93126, w_eco93127, w_eco93128, w_eco93129, w_eco93130, w_eco93131, w_eco93132, w_eco93133, w_eco93134, w_eco93135, w_eco93136, w_eco93137, w_eco93138, w_eco93139, w_eco93140, w_eco93141, w_eco93142, w_eco93143, w_eco93144, w_eco93145, w_eco93146, w_eco93147, w_eco93148, w_eco93149, w_eco93150, w_eco93151, w_eco93152, w_eco93153, w_eco93154, w_eco93155, w_eco93156, w_eco93157, w_eco93158, w_eco93159, w_eco93160, w_eco93161, w_eco93162, w_eco93163, w_eco93164, w_eco93165, w_eco93166, w_eco93167, w_eco93168, w_eco93169, w_eco93170, w_eco93171, w_eco93172, w_eco93173, w_eco93174, w_eco93175, w_eco93176, w_eco93177, w_eco93178, w_eco93179, w_eco93180, w_eco93181, w_eco93182, w_eco93183, w_eco93184, w_eco93185, w_eco93186, w_eco93187, w_eco93188, w_eco93189, w_eco93190, w_eco93191, w_eco93192, w_eco93193, w_eco93194, w_eco93195, w_eco93196, w_eco93197, w_eco93198, w_eco93199, w_eco93200, w_eco93201, w_eco93202, w_eco93203, w_eco93204, w_eco93205, w_eco93206, w_eco93207, w_eco93208, w_eco93209, w_eco93210, w_eco93211, w_eco93212, w_eco93213, w_eco93214, w_eco93215, w_eco93216, w_eco93217, w_eco93218, w_eco93219, w_eco93220, w_eco93221, w_eco93222, w_eco93223, w_eco93224, w_eco93225, w_eco93226, w_eco93227, w_eco93228, w_eco93229, w_eco93230, w_eco93231, w_eco93232, w_eco93233, w_eco93234, w_eco93235, w_eco93236, w_eco93237, w_eco93238, w_eco93239, w_eco93240, w_eco93241, w_eco93242, w_eco93243, w_eco93244, w_eco93245, w_eco93246, w_eco93247, w_eco93248, w_eco93249, w_eco93250, w_eco93251, w_eco93252, w_eco93253, w_eco93254, w_eco93255, w_eco93256, w_eco93257, w_eco93258, w_eco93259, w_eco93260, w_eco93261, w_eco93262, w_eco93263, w_eco93264, w_eco93265, w_eco93266, w_eco93267, w_eco93268, w_eco93269, w_eco93270, w_eco93271, w_eco93272, w_eco93273, w_eco93274, w_eco93275, w_eco93276, w_eco93277, w_eco93278, w_eco93279, w_eco93280, w_eco93281, w_eco93282, w_eco93283, w_eco93284, w_eco93285, w_eco93286, w_eco93287, w_eco93288, w_eco93289, w_eco93290, w_eco93291, w_eco93292, w_eco93293, w_eco93294, w_eco93295, w_eco93296, w_eco93297, w_eco93298, w_eco93299, w_eco93300, w_eco93301, w_eco93302, w_eco93303, w_eco93304, w_eco93305, w_eco93306, w_eco93307, w_eco93308, w_eco93309, w_eco93310, w_eco93311, w_eco93312, w_eco93313, w_eco93314, w_eco93315, w_eco93316, w_eco93317, w_eco93318, w_eco93319, w_eco93320, w_eco93321, w_eco93322, w_eco93323, w_eco93324, w_eco93325, w_eco93326, w_eco93327, w_eco93328, w_eco93329, w_eco93330, w_eco93331, w_eco93332, w_eco93333, w_eco93334, w_eco93335, w_eco93336, w_eco93337, w_eco93338, w_eco93339, w_eco93340, w_eco93341, w_eco93342, w_eco93343, w_eco93344, w_eco93345, w_eco93346, w_eco93347, w_eco93348, w_eco93349, w_eco93350, w_eco93351, w_eco93352, w_eco93353, w_eco93354, w_eco93355, w_eco93356, w_eco93357, w_eco93358, w_eco93359, w_eco93360, w_eco93361, w_eco93362, w_eco93363, w_eco93364, w_eco93365, w_eco93366, w_eco93367, w_eco93368, w_eco93369, w_eco93370, w_eco93371, w_eco93372, w_eco93373, w_eco93374, w_eco93375, w_eco93376, w_eco93377, w_eco93378, w_eco93379, w_eco93380, w_eco93381, w_eco93382, w_eco93383, w_eco93384, w_eco93385, w_eco93386, w_eco93387, w_eco93388, w_eco93389, w_eco93390, w_eco93391, w_eco93392, w_eco93393, w_eco93394, w_eco93395, w_eco93396, w_eco93397, w_eco93398, w_eco93399, w_eco93400, w_eco93401, w_eco93402, w_eco93403, w_eco93404, w_eco93405, w_eco93406, w_eco93407, w_eco93408, w_eco93409, w_eco93410, w_eco93411, w_eco93412, w_eco93413, w_eco93414, w_eco93415, w_eco93416, w_eco93417, w_eco93418, w_eco93419, w_eco93420, w_eco93421, w_eco93422, w_eco93423, w_eco93424, w_eco93425, w_eco93426, w_eco93427, w_eco93428, w_eco93429, w_eco93430, w_eco93431, w_eco93432, w_eco93433, w_eco93434, w_eco93435, w_eco93436, w_eco93437, w_eco93438, w_eco93439, w_eco93440, w_eco93441, w_eco93442, w_eco93443, w_eco93444, w_eco93445, w_eco93446, w_eco93447, w_eco93448, w_eco93449, w_eco93450, w_eco93451, w_eco93452, w_eco93453, w_eco93454, w_eco93455, w_eco93456, w_eco93457, w_eco93458, w_eco93459, w_eco93460, w_eco93461, w_eco93462, w_eco93463, w_eco93464, w_eco93465, w_eco93466, w_eco93467, w_eco93468, w_eco93469, w_eco93470, w_eco93471, w_eco93472, w_eco93473, w_eco93474, w_eco93475, w_eco93476, w_eco93477, w_eco93478, w_eco93479, w_eco93480, w_eco93481, w_eco93482, w_eco93483, w_eco93484, w_eco93485, w_eco93486, w_eco93487, w_eco93488, w_eco93489, w_eco93490, w_eco93491, w_eco93492, w_eco93493, w_eco93494, w_eco93495, w_eco93496, w_eco93497, w_eco93498, w_eco93499, w_eco93500, w_eco93501, w_eco93502, w_eco93503, w_eco93504, w_eco93505, w_eco93506, w_eco93507, w_eco93508, w_eco93509, w_eco93510, w_eco93511, w_eco93512, w_eco93513, w_eco93514, w_eco93515, w_eco93516, w_eco93517, w_eco93518, w_eco93519, w_eco93520, w_eco93521, w_eco93522, w_eco93523, w_eco93524, w_eco93525, w_eco93526, w_eco93527, w_eco93528, w_eco93529, w_eco93530, w_eco93531, w_eco93532, w_eco93533, w_eco93534, w_eco93535, w_eco93536, w_eco93537, w_eco93538, w_eco93539, w_eco93540, w_eco93541, w_eco93542, w_eco93543, w_eco93544, w_eco93545, w_eco93546, w_eco93547, w_eco93548, w_eco93549, w_eco93550, w_eco93551, w_eco93552, w_eco93553, w_eco93554, w_eco93555, w_eco93556, w_eco93557, w_eco93558, w_eco93559, w_eco93560, w_eco93561, w_eco93562, w_eco93563, w_eco93564, w_eco93565, w_eco93566, w_eco93567, w_eco93568, w_eco93569, w_eco93570, w_eco93571, w_eco93572, w_eco93573, w_eco93574, w_eco93575, w_eco93576, w_eco93577, w_eco93578, w_eco93579, w_eco93580, w_eco93581, w_eco93582, w_eco93583, w_eco93584, w_eco93585, w_eco93586, w_eco93587, w_eco93588, w_eco93589, w_eco93590, w_eco93591, w_eco93592, w_eco93593, w_eco93594, w_eco93595, w_eco93596, w_eco93597, w_eco93598, w_eco93599, w_eco93600, w_eco93601, w_eco93602, w_eco93603, w_eco93604, w_eco93605, w_eco93606, w_eco93607, w_eco93608, w_eco93609, w_eco93610, w_eco93611, w_eco93612, w_eco93613, w_eco93614, w_eco93615, w_eco93616, w_eco93617, w_eco93618, w_eco93619, w_eco93620, w_eco93621, w_eco93622, w_eco93623, w_eco93624, w_eco93625, w_eco93626, w_eco93627, w_eco93628, w_eco93629, w_eco93630, w_eco93631, w_eco93632, w_eco93633, w_eco93634, w_eco93635, w_eco93636, w_eco93637, w_eco93638, w_eco93639, w_eco93640, w_eco93641, w_eco93642, w_eco93643, w_eco93644, w_eco93645, w_eco93646, w_eco93647, w_eco93648, w_eco93649, w_eco93650, w_eco93651, w_eco93652, w_eco93653, w_eco93654, w_eco93655, w_eco93656, w_eco93657, w_eco93658, w_eco93659, w_eco93660, w_eco93661, w_eco93662, w_eco93663, w_eco93664, w_eco93665, w_eco93666, w_eco93667, w_eco93668, w_eco93669, w_eco93670, w_eco93671, w_eco93672, w_eco93673, w_eco93674, w_eco93675, w_eco93676, w_eco93677, w_eco93678, w_eco93679, w_eco93680, w_eco93681, w_eco93682, w_eco93683, w_eco93684, w_eco93685, w_eco93686, w_eco93687, w_eco93688, w_eco93689, w_eco93690, w_eco93691, w_eco93692, w_eco93693, w_eco93694, w_eco93695, w_eco93696, w_eco93697, w_eco93698, w_eco93699, w_eco93700, w_eco93701, w_eco93702, w_eco93703, w_eco93704, w_eco93705, w_eco93706, w_eco93707, w_eco93708, w_eco93709, w_eco93710, w_eco93711, w_eco93712, w_eco93713, w_eco93714, w_eco93715, w_eco93716, w_eco93717, w_eco93718, w_eco93719, w_eco93720, w_eco93721, w_eco93722, w_eco93723, w_eco93724, w_eco93725, w_eco93726, w_eco93727, w_eco93728, w_eco93729, w_eco93730, w_eco93731, w_eco93732, w_eco93733, w_eco93734, w_eco93735, w_eco93736, w_eco93737, w_eco93738, w_eco93739, w_eco93740, w_eco93741, w_eco93742, w_eco93743, w_eco93744, w_eco93745, w_eco93746, w_eco93747, w_eco93748, w_eco93749, w_eco93750, w_eco93751, w_eco93752, w_eco93753, w_eco93754, w_eco93755, w_eco93756, w_eco93757, w_eco93758, w_eco93759, w_eco93760, w_eco93761, w_eco93762, w_eco93763, w_eco93764, w_eco93765, w_eco93766, w_eco93767, w_eco93768, w_eco93769, w_eco93770, w_eco93771, w_eco93772, w_eco93773, w_eco93774, w_eco93775, w_eco93776, w_eco93777, w_eco93778, w_eco93779, w_eco93780, w_eco93781, w_eco93782, w_eco93783, w_eco93784, w_eco93785, w_eco93786, w_eco93787, w_eco93788, w_eco93789, w_eco93790, w_eco93791, w_eco93792, w_eco93793, w_eco93794, w_eco93795, w_eco93796, w_eco93797, w_eco93798, w_eco93799, w_eco93800, w_eco93801, w_eco93802, w_eco93803, w_eco93804, w_eco93805, w_eco93806, w_eco93807, w_eco93808, w_eco93809, w_eco93810, w_eco93811, w_eco93812, w_eco93813, w_eco93814, w_eco93815, w_eco93816, w_eco93817, w_eco93818, w_eco93819, w_eco93820, w_eco93821, w_eco93822, w_eco93823, w_eco93824, w_eco93825, w_eco93826, w_eco93827, w_eco93828, w_eco93829, w_eco93830, w_eco93831, w_eco93832, w_eco93833, w_eco93834, w_eco93835, w_eco93836, w_eco93837, w_eco93838, w_eco93839, w_eco93840, w_eco93841, w_eco93842, w_eco93843, w_eco93844, w_eco93845, w_eco93846, w_eco93847, w_eco93848, w_eco93849, w_eco93850, w_eco93851, w_eco93852, w_eco93853, w_eco93854, w_eco93855, w_eco93856, w_eco93857, w_eco93858, w_eco93859, w_eco93860, w_eco93861, w_eco93862, w_eco93863, w_eco93864, w_eco93865, w_eco93866, w_eco93867, w_eco93868, w_eco93869, w_eco93870, w_eco93871, w_eco93872, w_eco93873, w_eco93874, w_eco93875, w_eco93876, w_eco93877, w_eco93878, w_eco93879, w_eco93880, w_eco93881, w_eco93882, w_eco93883, w_eco93884, w_eco93885, w_eco93886, w_eco93887, w_eco93888, w_eco93889, w_eco93890, w_eco93891, w_eco93892, w_eco93893, w_eco93894, w_eco93895, w_eco93896, w_eco93897, w_eco93898, w_eco93899, w_eco93900, w_eco93901, w_eco93902, w_eco93903, w_eco93904, w_eco93905, w_eco93906, w_eco93907, w_eco93908, w_eco93909, w_eco93910, w_eco93911, w_eco93912, w_eco93913, w_eco93914, w_eco93915, w_eco93916, w_eco93917, w_eco93918, w_eco93919, w_eco93920, w_eco93921, w_eco93922, w_eco93923, w_eco93924, w_eco93925, w_eco93926, w_eco93927, w_eco93928, w_eco93929, w_eco93930, w_eco93931, w_eco93932, w_eco93933, w_eco93934, w_eco93935, w_eco93936, w_eco93937, w_eco93938, w_eco93939, w_eco93940, w_eco93941, w_eco93942, w_eco93943, w_eco93944, w_eco93945, w_eco93946, w_eco93947, w_eco93948, w_eco93949, w_eco93950, w_eco93951, w_eco93952, w_eco93953, w_eco93954, w_eco93955, w_eco93956, w_eco93957, w_eco93958, w_eco93959, w_eco93960, w_eco93961, w_eco93962, w_eco93963, w_eco93964, w_eco93965, w_eco93966, w_eco93967, w_eco93968, w_eco93969, w_eco93970, w_eco93971, w_eco93972, w_eco93973, w_eco93974, w_eco93975, w_eco93976, w_eco93977, w_eco93978, w_eco93979, w_eco93980, w_eco93981, w_eco93982, w_eco93983, w_eco93984, w_eco93985, w_eco93986, w_eco93987, w_eco93988, w_eco93989, w_eco93990, w_eco93991, w_eco93992, w_eco93993, w_eco93994, w_eco93995, w_eco93996, w_eco93997, w_eco93998, w_eco93999, w_eco94000, w_eco94001, w_eco94002, w_eco94003, w_eco94004, w_eco94005, w_eco94006, w_eco94007, w_eco94008, w_eco94009, w_eco94010, w_eco94011, w_eco94012, w_eco94013, w_eco94014, w_eco94015, w_eco94016, w_eco94017, w_eco94018, w_eco94019, w_eco94020, w_eco94021, w_eco94022, w_eco94023, w_eco94024, w_eco94025, w_eco94026, w_eco94027, w_eco94028, w_eco94029, w_eco94030, w_eco94031, w_eco94032, w_eco94033, w_eco94034, w_eco94035, w_eco94036, w_eco94037, w_eco94038, w_eco94039, w_eco94040, w_eco94041, w_eco94042, w_eco94043, w_eco94044, w_eco94045, w_eco94046, w_eco94047, w_eco94048, w_eco94049, w_eco94050, w_eco94051, w_eco94052, w_eco94053, w_eco94054, w_eco94055, w_eco94056, w_eco94057, w_eco94058, w_eco94059, w_eco94060, w_eco94061, w_eco94062, w_eco94063, w_eco94064, w_eco94065, w_eco94066, w_eco94067, w_eco94068, w_eco94069, w_eco94070, w_eco94071, w_eco94072, w_eco94073, w_eco94074, w_eco94075, w_eco94076, w_eco94077, w_eco94078, w_eco94079, w_eco94080, w_eco94081, w_eco94082, w_eco94083, w_eco94084, w_eco94085, w_eco94086, w_eco94087, w_eco94088, w_eco94089, w_eco94090, w_eco94091, w_eco94092, w_eco94093, w_eco94094, w_eco94095, w_eco94096, w_eco94097, w_eco94098, w_eco94099, w_eco94100, w_eco94101, w_eco94102, w_eco94103, w_eco94104, w_eco94105, w_eco94106, w_eco94107, w_eco94108, w_eco94109, w_eco94110, w_eco94111, w_eco94112, w_eco94113, w_eco94114, w_eco94115, w_eco94116, w_eco94117, w_eco94118, w_eco94119, w_eco94120, w_eco94121, w_eco94122, w_eco94123, w_eco94124, w_eco94125, w_eco94126, w_eco94127, w_eco94128, w_eco94129, w_eco94130, w_eco94131, w_eco94132, w_eco94133, w_eco94134, w_eco94135, w_eco94136, w_eco94137, w_eco94138, w_eco94139, w_eco94140, w_eco94141, w_eco94142, w_eco94143, w_eco94144, w_eco94145, w_eco94146, w_eco94147, w_eco94148, w_eco94149, w_eco94150, w_eco94151, w_eco94152, w_eco94153, w_eco94154, w_eco94155, w_eco94156, w_eco94157, w_eco94158, w_eco94159, w_eco94160, w_eco94161, w_eco94162, w_eco94163, w_eco94164, w_eco94165, w_eco94166, w_eco94167, w_eco94168, w_eco94169, w_eco94170, w_eco94171, w_eco94172, w_eco94173, w_eco94174, w_eco94175, w_eco94176, w_eco94177, w_eco94178, w_eco94179, w_eco94180, w_eco94181, w_eco94182, w_eco94183, w_eco94184, w_eco94185, w_eco94186, w_eco94187, w_eco94188, w_eco94189, w_eco94190, w_eco94191, w_eco94192, w_eco94193, w_eco94194, w_eco94195, w_eco94196, w_eco94197, w_eco94198, w_eco94199, w_eco94200, w_eco94201, w_eco94202, w_eco94203, w_eco94204, w_eco94205, w_eco94206, w_eco94207, w_eco94208, w_eco94209, w_eco94210, w_eco94211, w_eco94212, w_eco94213, w_eco94214, w_eco94215, w_eco94216, w_eco94217, w_eco94218, w_eco94219, w_eco94220, w_eco94221, w_eco94222, w_eco94223, w_eco94224, w_eco94225, w_eco94226, w_eco94227, w_eco94228, w_eco94229, w_eco94230, w_eco94231, w_eco94232, w_eco94233, w_eco94234, w_eco94235, w_eco94236, w_eco94237, w_eco94238, w_eco94239, w_eco94240, w_eco94241, w_eco94242, w_eco94243, w_eco94244, w_eco94245, w_eco94246, w_eco94247, w_eco94248, w_eco94249, w_eco94250, w_eco94251, w_eco94252, w_eco94253, w_eco94254, w_eco94255, w_eco94256, w_eco94257, w_eco94258, w_eco94259, w_eco94260, w_eco94261, w_eco94262, w_eco94263, w_eco94264, w_eco94265, w_eco94266, w_eco94267, w_eco94268, w_eco94269, w_eco94270, w_eco94271, w_eco94272, w_eco94273, w_eco94274, w_eco94275, w_eco94276, w_eco94277, w_eco94278, w_eco94279, w_eco94280, w_eco94281, w_eco94282, w_eco94283, w_eco94284, w_eco94285, w_eco94286, w_eco94287, w_eco94288, w_eco94289, w_eco94290, w_eco94291, w_eco94292, w_eco94293, w_eco94294, w_eco94295, w_eco94296, w_eco94297, w_eco94298, w_eco94299, w_eco94300, w_eco94301, w_eco94302, w_eco94303, w_eco94304, w_eco94305, w_eco94306, w_eco94307, w_eco94308, w_eco94309, w_eco94310, w_eco94311, w_eco94312, w_eco94313, w_eco94314, w_eco94315, w_eco94316, w_eco94317, w_eco94318, w_eco94319, w_eco94320, w_eco94321, w_eco94322, w_eco94323, w_eco94324, w_eco94325, w_eco94326, w_eco94327, w_eco94328, w_eco94329, w_eco94330, w_eco94331, w_eco94332, w_eco94333, w_eco94334, w_eco94335, w_eco94336, w_eco94337, w_eco94338, w_eco94339, w_eco94340, w_eco94341, w_eco94342, w_eco94343, w_eco94344, w_eco94345, w_eco94346, w_eco94347, w_eco94348, w_eco94349, w_eco94350, w_eco94351, w_eco94352, w_eco94353, w_eco94354, w_eco94355, w_eco94356, w_eco94357, w_eco94358, w_eco94359, w_eco94360, w_eco94361, w_eco94362, w_eco94363, w_eco94364, w_eco94365, w_eco94366, w_eco94367, w_eco94368, w_eco94369, w_eco94370, w_eco94371, w_eco94372, w_eco94373, w_eco94374, w_eco94375, w_eco94376, w_eco94377, w_eco94378, w_eco94379, w_eco94380, w_eco94381, w_eco94382, w_eco94383, w_eco94384, w_eco94385, w_eco94386, w_eco94387, w_eco94388, w_eco94389, w_eco94390, w_eco94391, w_eco94392, w_eco94393, w_eco94394, w_eco94395, w_eco94396, w_eco94397, w_eco94398, w_eco94399, w_eco94400, w_eco94401, w_eco94402, w_eco94403, w_eco94404, w_eco94405, w_eco94406, w_eco94407, w_eco94408, w_eco94409, w_eco94410, w_eco94411, w_eco94412, w_eco94413, w_eco94414, w_eco94415, w_eco94416, w_eco94417, w_eco94418, w_eco94419, w_eco94420, w_eco94421, w_eco94422, w_eco94423, w_eco94424, w_eco94425, w_eco94426, w_eco94427, w_eco94428, w_eco94429, w_eco94430, w_eco94431, w_eco94432, w_eco94433, w_eco94434, w_eco94435, w_eco94436, w_eco94437, w_eco94438, w_eco94439, w_eco94440, w_eco94441, w_eco94442, w_eco94443, w_eco94444, w_eco94445, w_eco94446, w_eco94447, w_eco94448, w_eco94449, w_eco94450, w_eco94451, w_eco94452, w_eco94453, w_eco94454, w_eco94455, w_eco94456, w_eco94457, w_eco94458, w_eco94459, w_eco94460, w_eco94461, w_eco94462, w_eco94463, w_eco94464, w_eco94465, w_eco94466, w_eco94467, w_eco94468, w_eco94469, w_eco94470, w_eco94471, w_eco94472, w_eco94473, w_eco94474, w_eco94475, w_eco94476, w_eco94477, w_eco94478, w_eco94479, w_eco94480, w_eco94481, w_eco94482, w_eco94483, w_eco94484, w_eco94485, w_eco94486, w_eco94487, w_eco94488, w_eco94489, w_eco94490, w_eco94491, w_eco94492, w_eco94493, w_eco94494, w_eco94495, w_eco94496, w_eco94497, w_eco94498, w_eco94499, w_eco94500, w_eco94501, w_eco94502, w_eco94503, w_eco94504, w_eco94505, w_eco94506, w_eco94507, w_eco94508, w_eco94509, w_eco94510, w_eco94511, w_eco94512, w_eco94513, w_eco94514, w_eco94515, w_eco94516, w_eco94517, w_eco94518, w_eco94519, w_eco94520, w_eco94521, w_eco94522, w_eco94523, w_eco94524, w_eco94525, w_eco94526, w_eco94527, w_eco94528, w_eco94529, w_eco94530, w_eco94531, w_eco94532, w_eco94533, w_eco94534, w_eco94535, w_eco94536, w_eco94537, w_eco94538, w_eco94539, w_eco94540, w_eco94541, w_eco94542, w_eco94543, w_eco94544, w_eco94545, w_eco94546, w_eco94547, w_eco94548, w_eco94549, w_eco94550, w_eco94551, w_eco94552, w_eco94553, w_eco94554, w_eco94555, w_eco94556, w_eco94557, w_eco94558, w_eco94559, w_eco94560, w_eco94561, w_eco94562, w_eco94563, w_eco94564, w_eco94565, w_eco94566, w_eco94567, w_eco94568, w_eco94569, w_eco94570, w_eco94571, w_eco94572, w_eco94573, w_eco94574, w_eco94575, w_eco94576, w_eco94577, w_eco94578, w_eco94579, w_eco94580, w_eco94581, w_eco94582, w_eco94583, w_eco94584, w_eco94585, w_eco94586, w_eco94587, w_eco94588, w_eco94589, w_eco94590, w_eco94591, w_eco94592, w_eco94593, w_eco94594, w_eco94595, w_eco94596, w_eco94597, w_eco94598, w_eco94599, w_eco94600, w_eco94601, w_eco94602, w_eco94603, w_eco94604, w_eco94605, w_eco94606, w_eco94607, w_eco94608, w_eco94609, w_eco94610, w_eco94611, w_eco94612, w_eco94613, w_eco94614, w_eco94615, w_eco94616, w_eco94617, w_eco94618, w_eco94619, w_eco94620, w_eco94621, w_eco94622, w_eco94623, w_eco94624, w_eco94625, w_eco94626, w_eco94627, w_eco94628, w_eco94629, w_eco94630, w_eco94631, w_eco94632, w_eco94633, w_eco94634, w_eco94635, w_eco94636, w_eco94637, w_eco94638, w_eco94639, w_eco94640, w_eco94641, w_eco94642, w_eco94643, w_eco94644, w_eco94645, w_eco94646, w_eco94647, w_eco94648, w_eco94649, w_eco94650, w_eco94651, w_eco94652, w_eco94653, w_eco94654, w_eco94655, w_eco94656, w_eco94657, w_eco94658, w_eco94659, w_eco94660, w_eco94661, w_eco94662, w_eco94663, w_eco94664, w_eco94665, w_eco94666, w_eco94667, w_eco94668, w_eco94669, w_eco94670, w_eco94671, w_eco94672, w_eco94673, w_eco94674, w_eco94675, w_eco94676, w_eco94677, w_eco94678, w_eco94679, w_eco94680, w_eco94681, w_eco94682, w_eco94683, w_eco94684, w_eco94685, w_eco94686, w_eco94687, w_eco94688, w_eco94689, w_eco94690, w_eco94691, w_eco94692, w_eco94693, w_eco94694, w_eco94695, w_eco94696, w_eco94697, w_eco94698, w_eco94699, w_eco94700, w_eco94701, w_eco94702, w_eco94703, w_eco94704, w_eco94705, w_eco94706, w_eco94707, w_eco94708, w_eco94709, w_eco94710, w_eco94711, w_eco94712, w_eco94713, w_eco94714, w_eco94715, w_eco94716, w_eco94717, w_eco94718, w_eco94719, w_eco94720, w_eco94721, w_eco94722, w_eco94723, w_eco94724, w_eco94725, w_eco94726, w_eco94727, w_eco94728, w_eco94729, w_eco94730, w_eco94731, w_eco94732, w_eco94733, w_eco94734, w_eco94735, w_eco94736, w_eco94737, w_eco94738, w_eco94739, w_eco94740, w_eco94741, w_eco94742, w_eco94743, w_eco94744, w_eco94745, w_eco94746, w_eco94747, w_eco94748, w_eco94749, w_eco94750, w_eco94751, w_eco94752, w_eco94753, w_eco94754, w_eco94755, w_eco94756, w_eco94757, w_eco94758, w_eco94759, w_eco94760, w_eco94761, w_eco94762, w_eco94763, w_eco94764, w_eco94765, w_eco94766, w_eco94767, w_eco94768, w_eco94769, w_eco94770, w_eco94771, w_eco94772, w_eco94773, w_eco94774, w_eco94775, w_eco94776, w_eco94777, w_eco94778, w_eco94779, w_eco94780, w_eco94781, w_eco94782, w_eco94783, w_eco94784, w_eco94785, w_eco94786, w_eco94787, w_eco94788, w_eco94789, w_eco94790, w_eco94791, w_eco94792, w_eco94793, w_eco94794, w_eco94795, w_eco94796, w_eco94797, w_eco94798, w_eco94799, w_eco94800, w_eco94801, w_eco94802, w_eco94803, w_eco94804, w_eco94805, w_eco94806, w_eco94807, w_eco94808, w_eco94809, w_eco94810, w_eco94811, w_eco94812, w_eco94813, w_eco94814, w_eco94815, w_eco94816, w_eco94817, w_eco94818, w_eco94819, w_eco94820, w_eco94821, w_eco94822, w_eco94823, w_eco94824, w_eco94825, w_eco94826, w_eco94827, w_eco94828, w_eco94829, w_eco94830, w_eco94831, w_eco94832, w_eco94833, w_eco94834, w_eco94835, w_eco94836, w_eco94837, w_eco94838, w_eco94839, w_eco94840, w_eco94841, w_eco94842, w_eco94843, w_eco94844, w_eco94845, w_eco94846, w_eco94847, w_eco94848, w_eco94849, w_eco94850, w_eco94851, w_eco94852, w_eco94853, w_eco94854, w_eco94855, w_eco94856, w_eco94857, w_eco94858, w_eco94859, w_eco94860, w_eco94861, w_eco94862, w_eco94863, w_eco94864, w_eco94865, w_eco94866, w_eco94867, w_eco94868, w_eco94869, w_eco94870, w_eco94871, w_eco94872, w_eco94873, w_eco94874, w_eco94875, w_eco94876, w_eco94877, w_eco94878, w_eco94879, w_eco94880, w_eco94881, w_eco94882, w_eco94883, w_eco94884, w_eco94885, w_eco94886, w_eco94887, w_eco94888, w_eco94889, w_eco94890, w_eco94891, w_eco94892, w_eco94893, w_eco94894, w_eco94895, w_eco94896, w_eco94897, w_eco94898, w_eco94899, w_eco94900, w_eco94901, w_eco94902, w_eco94903, w_eco94904, w_eco94905, w_eco94906, w_eco94907, w_eco94908, w_eco94909, w_eco94910, w_eco94911, w_eco94912, w_eco94913, w_eco94914, w_eco94915, w_eco94916, w_eco94917, w_eco94918, w_eco94919, w_eco94920, w_eco94921, w_eco94922, w_eco94923, w_eco94924, w_eco94925, w_eco94926, w_eco94927, w_eco94928, w_eco94929, w_eco94930, w_eco94931, w_eco94932, w_eco94933, w_eco94934, w_eco94935, w_eco94936, w_eco94937, w_eco94938, w_eco94939, w_eco94940, w_eco94941, w_eco94942, w_eco94943, w_eco94944, w_eco94945, w_eco94946, w_eco94947, w_eco94948, w_eco94949, w_eco94950, w_eco94951, w_eco94952, w_eco94953, w_eco94954, w_eco94955, w_eco94956, w_eco94957, w_eco94958, w_eco94959, w_eco94960, w_eco94961, w_eco94962, w_eco94963, w_eco94964, w_eco94965, w_eco94966, w_eco94967, w_eco94968, w_eco94969, w_eco94970, w_eco94971, w_eco94972, w_eco94973, w_eco94974, w_eco94975, w_eco94976, w_eco94977, w_eco94978, w_eco94979, w_eco94980, w_eco94981, w_eco94982, w_eco94983, w_eco94984, w_eco94985, w_eco94986, w_eco94987, w_eco94988, w_eco94989, w_eco94990, w_eco94991, w_eco94992, w_eco94993, w_eco94994, w_eco94995, w_eco94996, w_eco94997, w_eco94998, w_eco94999, w_eco95000, w_eco95001, w_eco95002, w_eco95003, w_eco95004, w_eco95005, w_eco95006, w_eco95007, w_eco95008, w_eco95009, w_eco95010, w_eco95011, w_eco95012, w_eco95013, w_eco95014, w_eco95015, w_eco95016, w_eco95017, w_eco95018, w_eco95019, w_eco95020, w_eco95021, w_eco95022, w_eco95023, w_eco95024, w_eco95025, w_eco95026, w_eco95027, w_eco95028, w_eco95029, w_eco95030, w_eco95031, w_eco95032, w_eco95033, w_eco95034, w_eco95035, w_eco95036, w_eco95037, w_eco95038, w_eco95039, w_eco95040, w_eco95041, w_eco95042, w_eco95043, w_eco95044, w_eco95045, w_eco95046, w_eco95047, w_eco95048, w_eco95049, w_eco95050, w_eco95051, w_eco95052, w_eco95053, w_eco95054, w_eco95055, w_eco95056, w_eco95057, w_eco95058, w_eco95059, w_eco95060, w_eco95061, w_eco95062, w_eco95063, w_eco95064, w_eco95065, w_eco95066, w_eco95067, w_eco95068, w_eco95069, w_eco95070, w_eco95071, w_eco95072, w_eco95073, w_eco95074, w_eco95075, w_eco95076, w_eco95077, w_eco95078, w_eco95079, w_eco95080, w_eco95081, w_eco95082, w_eco95083, w_eco95084, w_eco95085, w_eco95086, w_eco95087, w_eco95088, w_eco95089, w_eco95090, w_eco95091, w_eco95092, w_eco95093, w_eco95094, w_eco95095, w_eco95096, w_eco95097, w_eco95098, w_eco95099, w_eco95100, w_eco95101, w_eco95102, w_eco95103, w_eco95104, w_eco95105, w_eco95106, w_eco95107, w_eco95108, w_eco95109, w_eco95110, w_eco95111, w_eco95112, w_eco95113, w_eco95114, w_eco95115, w_eco95116, w_eco95117, w_eco95118, w_eco95119, w_eco95120, w_eco95121, w_eco95122, w_eco95123, w_eco95124, w_eco95125, w_eco95126, w_eco95127, w_eco95128, w_eco95129, w_eco95130, w_eco95131, w_eco95132, w_eco95133, w_eco95134, w_eco95135, w_eco95136, w_eco95137, w_eco95138, w_eco95139, w_eco95140, w_eco95141, w_eco95142, w_eco95143, w_eco95144, w_eco95145, w_eco95146, w_eco95147, w_eco95148, w_eco95149, w_eco95150, w_eco95151, w_eco95152, w_eco95153, w_eco95154, w_eco95155, w_eco95156, w_eco95157, w_eco95158, w_eco95159, w_eco95160, w_eco95161, w_eco95162, w_eco95163, w_eco95164, w_eco95165, w_eco95166, w_eco95167, w_eco95168, w_eco95169, w_eco95170, w_eco95171, w_eco95172, w_eco95173, w_eco95174, w_eco95175, w_eco95176, w_eco95177, w_eco95178, w_eco95179, w_eco95180, w_eco95181, w_eco95182, w_eco95183, w_eco95184, w_eco95185, w_eco95186, w_eco95187, w_eco95188, w_eco95189, w_eco95190, w_eco95191, w_eco95192, w_eco95193, w_eco95194, w_eco95195, w_eco95196, w_eco95197, w_eco95198, w_eco95199, w_eco95200, w_eco95201, w_eco95202, w_eco95203, w_eco95204, w_eco95205, w_eco95206, w_eco95207, w_eco95208, w_eco95209, w_eco95210, w_eco95211, w_eco95212, w_eco95213, w_eco95214, w_eco95215, w_eco95216, w_eco95217, w_eco95218, w_eco95219, w_eco95220, w_eco95221, w_eco95222, w_eco95223, w_eco95224, w_eco95225, w_eco95226, w_eco95227, w_eco95228, w_eco95229, w_eco95230, w_eco95231, w_eco95232, w_eco95233, w_eco95234, w_eco95235, w_eco95236, w_eco95237, w_eco95238, w_eco95239, w_eco95240, w_eco95241, w_eco95242, w_eco95243, w_eco95244, w_eco95245, w_eco95246, w_eco95247, w_eco95248, w_eco95249, w_eco95250, w_eco95251, w_eco95252, w_eco95253, w_eco95254, w_eco95255, w_eco95256, w_eco95257, w_eco95258, w_eco95259, w_eco95260, w_eco95261, w_eco95262, w_eco95263, w_eco95264, w_eco95265, w_eco95266, w_eco95267, w_eco95268, w_eco95269, w_eco95270, w_eco95271, w_eco95272, w_eco95273, w_eco95274, w_eco95275, w_eco95276, w_eco95277, w_eco95278, w_eco95279, w_eco95280, w_eco95281, w_eco95282, w_eco95283, w_eco95284, w_eco95285, w_eco95286, w_eco95287, w_eco95288, w_eco95289, w_eco95290, w_eco95291, w_eco95292, w_eco95293, w_eco95294, w_eco95295, w_eco95296, w_eco95297, w_eco95298, w_eco95299, w_eco95300, w_eco95301, w_eco95302, w_eco95303, w_eco95304, w_eco95305, w_eco95306, w_eco95307, w_eco95308, w_eco95309, w_eco95310, w_eco95311, w_eco95312, w_eco95313, w_eco95314, w_eco95315, w_eco95316, w_eco95317, w_eco95318, w_eco95319, w_eco95320, w_eco95321, w_eco95322, w_eco95323, w_eco95324, w_eco95325, w_eco95326, w_eco95327, w_eco95328, w_eco95329, w_eco95330, w_eco95331, w_eco95332, w_eco95333, w_eco95334, w_eco95335, w_eco95336, w_eco95337, w_eco95338, w_eco95339, w_eco95340, w_eco95341, w_eco95342, w_eco95343, w_eco95344, w_eco95345, w_eco95346, w_eco95347, w_eco95348, w_eco95349, w_eco95350, w_eco95351, w_eco95352, w_eco95353, w_eco95354, w_eco95355, w_eco95356, w_eco95357, w_eco95358, w_eco95359, w_eco95360, w_eco95361, w_eco95362, w_eco95363, w_eco95364, w_eco95365, w_eco95366, w_eco95367, w_eco95368, w_eco95369, w_eco95370, w_eco95371, w_eco95372, w_eco95373, w_eco95374, w_eco95375, w_eco95376, w_eco95377, w_eco95378, w_eco95379, w_eco95380, w_eco95381, w_eco95382, w_eco95383, w_eco95384, w_eco95385, w_eco95386, w_eco95387, w_eco95388, w_eco95389, w_eco95390, w_eco95391, w_eco95392, w_eco95393, w_eco95394, w_eco95395, w_eco95396, w_eco95397, w_eco95398, w_eco95399, w_eco95400, w_eco95401, w_eco95402, w_eco95403, w_eco95404, w_eco95405, w_eco95406, w_eco95407, w_eco95408, w_eco95409, w_eco95410, w_eco95411, w_eco95412, w_eco95413, w_eco95414, w_eco95415, w_eco95416, w_eco95417, w_eco95418, w_eco95419, w_eco95420, w_eco95421, w_eco95422, w_eco95423, w_eco95424, w_eco95425, w_eco95426, w_eco95427, w_eco95428, w_eco95429, w_eco95430, w_eco95431, w_eco95432, w_eco95433, w_eco95434, w_eco95435, w_eco95436, w_eco95437, w_eco95438, w_eco95439, w_eco95440, w_eco95441, w_eco95442, w_eco95443, w_eco95444, w_eco95445, w_eco95446, w_eco95447, w_eco95448, w_eco95449, w_eco95450, w_eco95451, w_eco95452, w_eco95453, w_eco95454, w_eco95455, w_eco95456, w_eco95457, w_eco95458, w_eco95459, w_eco95460, w_eco95461, w_eco95462, w_eco95463, w_eco95464, w_eco95465, w_eco95466, w_eco95467, w_eco95468, w_eco95469, w_eco95470, w_eco95471, w_eco95472, w_eco95473, w_eco95474, w_eco95475, w_eco95476, w_eco95477, w_eco95478, w_eco95479, w_eco95480, w_eco95481, w_eco95482, w_eco95483, w_eco95484, w_eco95485, w_eco95486, w_eco95487, w_eco95488, w_eco95489, w_eco95490, w_eco95491, w_eco95492, w_eco95493, w_eco95494, w_eco95495, w_eco95496, w_eco95497, w_eco95498, w_eco95499, w_eco95500, w_eco95501, w_eco95502, w_eco95503, w_eco95504, w_eco95505, w_eco95506, w_eco95507, w_eco95508, w_eco95509, w_eco95510, w_eco95511, w_eco95512, w_eco95513, w_eco95514, w_eco95515, w_eco95516, w_eco95517, w_eco95518, w_eco95519, w_eco95520, w_eco95521, w_eco95522, w_eco95523, w_eco95524, w_eco95525, w_eco95526, w_eco95527, w_eco95528, w_eco95529, w_eco95530, w_eco95531, w_eco95532, w_eco95533, w_eco95534, w_eco95535, w_eco95536, w_eco95537, w_eco95538, w_eco95539, w_eco95540, w_eco95541, w_eco95542, w_eco95543, w_eco95544, w_eco95545, w_eco95546, w_eco95547, w_eco95548, w_eco95549, w_eco95550, w_eco95551, w_eco95552, w_eco95553, w_eco95554, w_eco95555, w_eco95556, w_eco95557, w_eco95558, w_eco95559, w_eco95560, w_eco95561, w_eco95562, w_eco95563, w_eco95564, w_eco95565, w_eco95566, w_eco95567, w_eco95568, w_eco95569, w_eco95570, w_eco95571, w_eco95572, w_eco95573, w_eco95574, w_eco95575, w_eco95576, w_eco95577, w_eco95578, w_eco95579, w_eco95580, w_eco95581, w_eco95582, w_eco95583, w_eco95584, w_eco95585, w_eco95586, w_eco95587, w_eco95588, w_eco95589, w_eco95590, w_eco95591, w_eco95592, w_eco95593, w_eco95594, w_eco95595, w_eco95596, w_eco95597, w_eco95598, w_eco95599, w_eco95600, w_eco95601, w_eco95602, w_eco95603, w_eco95604, w_eco95605, w_eco95606, w_eco95607, w_eco95608, w_eco95609, w_eco95610, w_eco95611, w_eco95612, w_eco95613, w_eco95614, w_eco95615, w_eco95616, w_eco95617, w_eco95618, w_eco95619, w_eco95620, w_eco95621, w_eco95622, w_eco95623, w_eco95624, w_eco95625, w_eco95626, w_eco95627, w_eco95628, w_eco95629, w_eco95630, w_eco95631, w_eco95632, w_eco95633, w_eco95634, w_eco95635, w_eco95636, w_eco95637, w_eco95638, w_eco95639, w_eco95640, w_eco95641, w_eco95642, w_eco95643, w_eco95644, w_eco95645, w_eco95646, w_eco95647, w_eco95648, w_eco95649, w_eco95650, w_eco95651, w_eco95652, w_eco95653, w_eco95654, w_eco95655, w_eco95656, w_eco95657, w_eco95658, w_eco95659, w_eco95660, w_eco95661, w_eco95662, w_eco95663, w_eco95664, w_eco95665, w_eco95666, w_eco95667, w_eco95668, w_eco95669, w_eco95670, w_eco95671, w_eco95672, w_eco95673, w_eco95674, w_eco95675, w_eco95676, w_eco95677, w_eco95678, w_eco95679, w_eco95680, w_eco95681, w_eco95682, w_eco95683, w_eco95684, w_eco95685, w_eco95686, w_eco95687, w_eco95688, w_eco95689, w_eco95690, w_eco95691, w_eco95692, w_eco95693, w_eco95694, w_eco95695, w_eco95696, w_eco95697, w_eco95698, w_eco95699, w_eco95700, w_eco95701, w_eco95702, w_eco95703, w_eco95704, w_eco95705, w_eco95706, w_eco95707, w_eco95708, w_eco95709, w_eco95710, w_eco95711, w_eco95712, w_eco95713, w_eco95714, w_eco95715, w_eco95716, w_eco95717, w_eco95718, w_eco95719, w_eco95720, w_eco95721, w_eco95722, w_eco95723, w_eco95724, w_eco95725, w_eco95726, w_eco95727, w_eco95728, w_eco95729, w_eco95730, w_eco95731, w_eco95732, w_eco95733, w_eco95734, w_eco95735, w_eco95736, w_eco95737, w_eco95738, w_eco95739, w_eco95740, w_eco95741, w_eco95742, w_eco95743, w_eco95744, w_eco95745, w_eco95746, w_eco95747, w_eco95748, w_eco95749, w_eco95750, w_eco95751, w_eco95752, w_eco95753, w_eco95754, w_eco95755, w_eco95756, w_eco95757, w_eco95758, w_eco95759, w_eco95760, w_eco95761, w_eco95762, w_eco95763, w_eco95764, w_eco95765, w_eco95766, w_eco95767, w_eco95768, w_eco95769, w_eco95770, w_eco95771, w_eco95772, w_eco95773, w_eco95774, w_eco95775, w_eco95776, w_eco95777, w_eco95778, w_eco95779, w_eco95780, w_eco95781, w_eco95782, w_eco95783, w_eco95784, w_eco95785, w_eco95786, w_eco95787, w_eco95788, w_eco95789, w_eco95790, w_eco95791, w_eco95792, w_eco95793, w_eco95794, w_eco95795, w_eco95796, w_eco95797, w_eco95798, w_eco95799, w_eco95800, w_eco95801, w_eco95802, w_eco95803, w_eco95804, w_eco95805, w_eco95806, w_eco95807, w_eco95808, w_eco95809, w_eco95810, w_eco95811, w_eco95812, w_eco95813, w_eco95814, w_eco95815, w_eco95816, w_eco95817, w_eco95818, w_eco95819, w_eco95820, w_eco95821, w_eco95822, w_eco95823, w_eco95824, w_eco95825, w_eco95826, w_eco95827, w_eco95828, w_eco95829, w_eco95830, w_eco95831, w_eco95832, w_eco95833, w_eco95834, w_eco95835, w_eco95836, w_eco95837, w_eco95838, w_eco95839, w_eco95840, w_eco95841, w_eco95842, w_eco95843, w_eco95844, w_eco95845, w_eco95846, w_eco95847, w_eco95848, w_eco95849, w_eco95850, w_eco95851, w_eco95852, w_eco95853, w_eco95854, w_eco95855, w_eco95856, w_eco95857, w_eco95858, w_eco95859, w_eco95860, w_eco95861, w_eco95862, w_eco95863, w_eco95864, w_eco95865, w_eco95866, w_eco95867, w_eco95868, w_eco95869, w_eco95870, w_eco95871, w_eco95872, w_eco95873, w_eco95874, w_eco95875, w_eco95876, w_eco95877, w_eco95878, w_eco95879, w_eco95880, w_eco95881, w_eco95882, w_eco95883, w_eco95884, w_eco95885, w_eco95886, w_eco95887, w_eco95888, w_eco95889, w_eco95890, w_eco95891, w_eco95892, w_eco95893, w_eco95894, w_eco95895, w_eco95896, w_eco95897, w_eco95898, w_eco95899, w_eco95900, w_eco95901, w_eco95902, w_eco95903, w_eco95904, w_eco95905, w_eco95906, w_eco95907, w_eco95908, w_eco95909, w_eco95910, w_eco95911, w_eco95912, w_eco95913, w_eco95914, w_eco95915, w_eco95916, w_eco95917, w_eco95918, w_eco95919, w_eco95920, w_eco95921, w_eco95922, w_eco95923, w_eco95924, w_eco95925, w_eco95926, w_eco95927, w_eco95928, w_eco95929, w_eco95930, w_eco95931, w_eco95932, w_eco95933, w_eco95934, w_eco95935, w_eco95936, w_eco95937, w_eco95938, w_eco95939, w_eco95940, w_eco95941, w_eco95942, w_eco95943, w_eco95944, w_eco95945, w_eco95946, w_eco95947, w_eco95948, w_eco95949, w_eco95950, w_eco95951, w_eco95952, w_eco95953, w_eco95954, w_eco95955, w_eco95956, w_eco95957, w_eco95958, w_eco95959, w_eco95960, w_eco95961, w_eco95962, w_eco95963, w_eco95964, w_eco95965, w_eco95966, w_eco95967, w_eco95968, w_eco95969, w_eco95970, w_eco95971, w_eco95972, w_eco95973, w_eco95974, w_eco95975, w_eco95976, w_eco95977, w_eco95978, w_eco95979, w_eco95980, w_eco95981, w_eco95982, w_eco95983, w_eco95984, w_eco95985, w_eco95986, w_eco95987, w_eco95988, w_eco95989, w_eco95990, w_eco95991, w_eco95992, w_eco95993, w_eco95994, w_eco95995, w_eco95996, w_eco95997, w_eco95998, w_eco95999, w_eco96000, w_eco96001, w_eco96002, w_eco96003, w_eco96004, w_eco96005, w_eco96006, w_eco96007, w_eco96008, w_eco96009, w_eco96010, w_eco96011, w_eco96012, w_eco96013, w_eco96014, w_eco96015, w_eco96016, w_eco96017, w_eco96018, w_eco96019, w_eco96020, w_eco96021, w_eco96022, w_eco96023, w_eco96024, w_eco96025, w_eco96026, w_eco96027, w_eco96028, w_eco96029, w_eco96030, w_eco96031, w_eco96032, w_eco96033, w_eco96034, w_eco96035, w_eco96036, w_eco96037, w_eco96038, w_eco96039, w_eco96040, w_eco96041, w_eco96042, w_eco96043, w_eco96044, w_eco96045, w_eco96046, w_eco96047, w_eco96048, w_eco96049, w_eco96050, w_eco96051, w_eco96052, w_eco96053, w_eco96054, w_eco96055, w_eco96056, w_eco96057, w_eco96058, w_eco96059, w_eco96060, w_eco96061, w_eco96062, w_eco96063, w_eco96064, w_eco96065, w_eco96066, w_eco96067, w_eco96068, w_eco96069, w_eco96070, w_eco96071, w_eco96072, w_eco96073, w_eco96074, w_eco96075, w_eco96076, w_eco96077, w_eco96078, w_eco96079, w_eco96080, w_eco96081, w_eco96082, w_eco96083, w_eco96084, w_eco96085, w_eco96086, w_eco96087, w_eco96088, w_eco96089, w_eco96090, w_eco96091, w_eco96092, w_eco96093, w_eco96094, w_eco96095, w_eco96096, w_eco96097, w_eco96098, w_eco96099, w_eco96100, w_eco96101, w_eco96102, w_eco96103, w_eco96104, w_eco96105, w_eco96106, w_eco96107, w_eco96108, w_eco96109, w_eco96110, w_eco96111, w_eco96112, w_eco96113, w_eco96114, w_eco96115, w_eco96116, w_eco96117, w_eco96118, w_eco96119, w_eco96120, w_eco96121, w_eco96122, w_eco96123, w_eco96124, w_eco96125, w_eco96126, w_eco96127, w_eco96128, w_eco96129, w_eco96130, w_eco96131, w_eco96132, w_eco96133, w_eco96134, w_eco96135, w_eco96136, w_eco96137, w_eco96138, w_eco96139, w_eco96140, w_eco96141, w_eco96142, w_eco96143, w_eco96144, w_eco96145, w_eco96146, w_eco96147, w_eco96148, w_eco96149, w_eco96150, w_eco96151, w_eco96152, w_eco96153, w_eco96154, w_eco96155, w_eco96156, w_eco96157, w_eco96158, w_eco96159, w_eco96160, w_eco96161, w_eco96162, w_eco96163, w_eco96164, w_eco96165, w_eco96166, w_eco96167, w_eco96168, w_eco96169, w_eco96170, w_eco96171, w_eco96172, w_eco96173, w_eco96174, w_eco96175, w_eco96176, w_eco96177, w_eco96178, w_eco96179, w_eco96180, w_eco96181, w_eco96182, w_eco96183, w_eco96184, w_eco96185, w_eco96186, w_eco96187, w_eco96188, w_eco96189, w_eco96190, w_eco96191, w_eco96192, w_eco96193, w_eco96194, w_eco96195, w_eco96196, w_eco96197, w_eco96198, w_eco96199, w_eco96200, w_eco96201, w_eco96202, w_eco96203, w_eco96204, w_eco96205, w_eco96206, w_eco96207, w_eco96208, w_eco96209, w_eco96210, w_eco96211, w_eco96212, w_eco96213, w_eco96214, w_eco96215, w_eco96216, w_eco96217, w_eco96218, w_eco96219, w_eco96220, w_eco96221, w_eco96222, w_eco96223, w_eco96224, w_eco96225, w_eco96226, w_eco96227, w_eco96228, w_eco96229, w_eco96230, w_eco96231, w_eco96232, w_eco96233, w_eco96234, w_eco96235, w_eco96236, w_eco96237, w_eco96238, w_eco96239, w_eco96240, w_eco96241, w_eco96242, w_eco96243, w_eco96244, w_eco96245, w_eco96246, w_eco96247, w_eco96248, w_eco96249, w_eco96250, w_eco96251, w_eco96252, w_eco96253, w_eco96254, w_eco96255, w_eco96256, w_eco96257, w_eco96258, w_eco96259, w_eco96260, w_eco96261, w_eco96262, w_eco96263, w_eco96264, w_eco96265, w_eco96266, w_eco96267, w_eco96268, w_eco96269, w_eco96270, w_eco96271, w_eco96272, w_eco96273, w_eco96274, w_eco96275, w_eco96276, w_eco96277, w_eco96278, w_eco96279, w_eco96280, w_eco96281, w_eco96282, w_eco96283, w_eco96284, w_eco96285, w_eco96286, w_eco96287, w_eco96288, w_eco96289, w_eco96290, w_eco96291, w_eco96292, w_eco96293, w_eco96294, w_eco96295, w_eco96296, w_eco96297, w_eco96298, w_eco96299, w_eco96300, w_eco96301, w_eco96302, w_eco96303, w_eco96304, w_eco96305, w_eco96306, w_eco96307, w_eco96308, w_eco96309, w_eco96310, w_eco96311, w_eco96312, w_eco96313, w_eco96314, w_eco96315, w_eco96316, w_eco96317, w_eco96318, w_eco96319, w_eco96320, w_eco96321, w_eco96322, w_eco96323, w_eco96324, w_eco96325, w_eco96326, w_eco96327, w_eco96328, w_eco96329, w_eco96330, w_eco96331, w_eco96332, w_eco96333, w_eco96334, w_eco96335, w_eco96336, w_eco96337, w_eco96338, w_eco96339, w_eco96340, w_eco96341, w_eco96342, w_eco96343, w_eco96344, w_eco96345, w_eco96346, w_eco96347, w_eco96348, w_eco96349, w_eco96350, w_eco96351, w_eco96352, w_eco96353, w_eco96354, w_eco96355, w_eco96356, w_eco96357, w_eco96358, w_eco96359, w_eco96360, w_eco96361, w_eco96362, w_eco96363, w_eco96364, w_eco96365, w_eco96366, w_eco96367, w_eco96368, w_eco96369, w_eco96370, w_eco96371, w_eco96372, w_eco96373, w_eco96374, w_eco96375, w_eco96376, w_eco96377, w_eco96378, w_eco96379, w_eco96380, w_eco96381, w_eco96382, w_eco96383, w_eco96384, w_eco96385, w_eco96386, w_eco96387, w_eco96388, w_eco96389, w_eco96390, w_eco96391, w_eco96392, w_eco96393, w_eco96394, w_eco96395, w_eco96396, w_eco96397, w_eco96398, w_eco96399, w_eco96400, w_eco96401, w_eco96402, w_eco96403, w_eco96404, w_eco96405, w_eco96406, w_eco96407, w_eco96408, w_eco96409, w_eco96410, w_eco96411, w_eco96412, w_eco96413, w_eco96414, w_eco96415, w_eco96416, w_eco96417, w_eco96418, w_eco96419, w_eco96420, w_eco96421, w_eco96422, w_eco96423, w_eco96424, w_eco96425, w_eco96426, w_eco96427, w_eco96428, w_eco96429, w_eco96430, w_eco96431, w_eco96432, w_eco96433, w_eco96434, w_eco96435, w_eco96436, w_eco96437, w_eco96438, w_eco96439, w_eco96440, w_eco96441, w_eco96442, w_eco96443, w_eco96444, w_eco96445, w_eco96446, w_eco96447, w_eco96448, w_eco96449, w_eco96450, w_eco96451, w_eco96452, w_eco96453, w_eco96454, w_eco96455, w_eco96456, w_eco96457, w_eco96458, w_eco96459, w_eco96460, w_eco96461, w_eco96462, w_eco96463, w_eco96464, w_eco96465, w_eco96466, w_eco96467, w_eco96468, w_eco96469, w_eco96470, w_eco96471, w_eco96472, w_eco96473, w_eco96474, w_eco96475, w_eco96476, w_eco96477, w_eco96478, w_eco96479, w_eco96480, w_eco96481, w_eco96482, w_eco96483, w_eco96484, w_eco96485, w_eco96486, w_eco96487, w_eco96488, w_eco96489, w_eco96490, w_eco96491, w_eco96492, w_eco96493, w_eco96494, w_eco96495, w_eco96496, w_eco96497, w_eco96498, w_eco96499, w_eco96500, w_eco96501, w_eco96502, w_eco96503, w_eco96504, w_eco96505, w_eco96506, w_eco96507, w_eco96508, w_eco96509, w_eco96510, w_eco96511, w_eco96512, w_eco96513, w_eco96514, w_eco96515, w_eco96516, w_eco96517, w_eco96518, w_eco96519, w_eco96520, w_eco96521, w_eco96522, w_eco96523, w_eco96524, w_eco96525, w_eco96526, w_eco96527, w_eco96528, w_eco96529, w_eco96530, w_eco96531, w_eco96532, w_eco96533, w_eco96534, w_eco96535, w_eco96536, w_eco96537, w_eco96538, w_eco96539, w_eco96540, w_eco96541, w_eco96542, w_eco96543, w_eco96544, w_eco96545, w_eco96546, w_eco96547, w_eco96548, w_eco96549, w_eco96550, w_eco96551, w_eco96552, w_eco96553, w_eco96554, w_eco96555, w_eco96556, w_eco96557, w_eco96558, w_eco96559, w_eco96560, w_eco96561, w_eco96562, w_eco96563, w_eco96564, w_eco96565, w_eco96566, w_eco96567, w_eco96568, w_eco96569, w_eco96570, w_eco96571, w_eco96572, w_eco96573, w_eco96574, w_eco96575, w_eco96576, w_eco96577, w_eco96578, w_eco96579, w_eco96580, w_eco96581, w_eco96582, w_eco96583, w_eco96584, w_eco96585, w_eco96586, w_eco96587, w_eco96588, w_eco96589, w_eco96590, w_eco96591, w_eco96592, w_eco96593, w_eco96594, w_eco96595, w_eco96596, w_eco96597, w_eco96598, w_eco96599, w_eco96600, w_eco96601, w_eco96602, w_eco96603, w_eco96604, w_eco96605, w_eco96606, w_eco96607, w_eco96608, w_eco96609, w_eco96610, w_eco96611, w_eco96612, w_eco96613, w_eco96614, w_eco96615, w_eco96616, w_eco96617, w_eco96618, w_eco96619, w_eco96620, w_eco96621, w_eco96622, w_eco96623, w_eco96624, w_eco96625, w_eco96626, w_eco96627, w_eco96628, w_eco96629, w_eco96630, w_eco96631, w_eco96632, w_eco96633, w_eco96634, w_eco96635, w_eco96636, w_eco96637, w_eco96638, w_eco96639, w_eco96640, w_eco96641, w_eco96642, w_eco96643, w_eco96644, w_eco96645, w_eco96646, w_eco96647, w_eco96648, w_eco96649, w_eco96650, w_eco96651, w_eco96652, w_eco96653, w_eco96654, w_eco96655, w_eco96656, w_eco96657, w_eco96658, w_eco96659, w_eco96660, w_eco96661, w_eco96662, w_eco96663, w_eco96664, w_eco96665, w_eco96666, w_eco96667, w_eco96668, w_eco96669, w_eco96670, w_eco96671, w_eco96672, w_eco96673, w_eco96674, w_eco96675, w_eco96676, w_eco96677, w_eco96678, w_eco96679, w_eco96680, w_eco96681, w_eco96682, w_eco96683, w_eco96684, w_eco96685, w_eco96686, w_eco96687, w_eco96688, w_eco96689, w_eco96690, w_eco96691, w_eco96692, w_eco96693, w_eco96694, w_eco96695, w_eco96696, w_eco96697, w_eco96698, w_eco96699, w_eco96700, w_eco96701, w_eco96702, w_eco96703, w_eco96704, w_eco96705, w_eco96706, w_eco96707, w_eco96708, w_eco96709, w_eco96710, w_eco96711, w_eco96712, w_eco96713, w_eco96714, w_eco96715, w_eco96716, w_eco96717, w_eco96718, w_eco96719, w_eco96720, w_eco96721, w_eco96722, w_eco96723, w_eco96724, w_eco96725, w_eco96726, w_eco96727, w_eco96728, w_eco96729, w_eco96730, w_eco96731, w_eco96732, w_eco96733, w_eco96734, w_eco96735, w_eco96736, w_eco96737, w_eco96738, w_eco96739, w_eco96740, w_eco96741, w_eco96742, w_eco96743, w_eco96744, w_eco96745, w_eco96746, w_eco96747, w_eco96748, w_eco96749, w_eco96750, w_eco96751, w_eco96752, w_eco96753, w_eco96754, w_eco96755, w_eco96756, w_eco96757, w_eco96758, w_eco96759, w_eco96760, w_eco96761, w_eco96762, w_eco96763, w_eco96764, w_eco96765, w_eco96766, w_eco96767, w_eco96768, w_eco96769, w_eco96770, w_eco96771, w_eco96772, w_eco96773, w_eco96774, w_eco96775, w_eco96776, w_eco96777, w_eco96778, w_eco96779, w_eco96780, w_eco96781, w_eco96782, w_eco96783, w_eco96784, w_eco96785, w_eco96786, w_eco96787, w_eco96788, w_eco96789, w_eco96790, w_eco96791, w_eco96792, w_eco96793, w_eco96794, w_eco96795, w_eco96796, w_eco96797, w_eco96798, w_eco96799, w_eco96800, w_eco96801, w_eco96802, w_eco96803, w_eco96804, w_eco96805, w_eco96806, w_eco96807, w_eco96808, w_eco96809, w_eco96810, w_eco96811, w_eco96812, w_eco96813, w_eco96814, w_eco96815, w_eco96816, w_eco96817, w_eco96818, w_eco96819, w_eco96820, w_eco96821, w_eco96822, w_eco96823, w_eco96824, w_eco96825, w_eco96826, w_eco96827, w_eco96828, w_eco96829, w_eco96830, w_eco96831, w_eco96832, w_eco96833, w_eco96834, w_eco96835, w_eco96836, w_eco96837, w_eco96838, w_eco96839, w_eco96840, w_eco96841, w_eco96842, w_eco96843, w_eco96844, w_eco96845, w_eco96846, w_eco96847, w_eco96848, w_eco96849, w_eco96850, w_eco96851, w_eco96852, w_eco96853, w_eco96854, w_eco96855, w_eco96856, w_eco96857, w_eco96858, w_eco96859, w_eco96860, w_eco96861, w_eco96862, w_eco96863, w_eco96864, w_eco96865, w_eco96866, w_eco96867, w_eco96868, w_eco96869, w_eco96870, w_eco96871, w_eco96872, w_eco96873, w_eco96874, w_eco96875, w_eco96876, w_eco96877, w_eco96878, w_eco96879, w_eco96880, w_eco96881, w_eco96882, w_eco96883, w_eco96884, w_eco96885, w_eco96886, w_eco96887, w_eco96888, w_eco96889, w_eco96890, w_eco96891, w_eco96892, w_eco96893, w_eco96894, w_eco96895, w_eco96896, w_eco96897, w_eco96898, w_eco96899, w_eco96900, w_eco96901, w_eco96902, w_eco96903, w_eco96904, w_eco96905, w_eco96906, w_eco96907, w_eco96908, w_eco96909, w_eco96910, w_eco96911, w_eco96912, w_eco96913, w_eco96914, w_eco96915, w_eco96916, w_eco96917, w_eco96918, w_eco96919, w_eco96920, w_eco96921, w_eco96922, w_eco96923, w_eco96924, w_eco96925, w_eco96926, w_eco96927, w_eco96928, w_eco96929, w_eco96930, w_eco96931, w_eco96932, w_eco96933, w_eco96934, w_eco96935, w_eco96936, w_eco96937, w_eco96938, w_eco96939, w_eco96940, w_eco96941, w_eco96942, w_eco96943, w_eco96944, w_eco96945, w_eco96946, w_eco96947, w_eco96948, w_eco96949, w_eco96950, w_eco96951, w_eco96952, w_eco96953, w_eco96954, w_eco96955, w_eco96956, w_eco96957, w_eco96958, w_eco96959, w_eco96960, w_eco96961, w_eco96962, w_eco96963, w_eco96964, w_eco96965, w_eco96966, w_eco96967, w_eco96968, w_eco96969, w_eco96970, w_eco96971, w_eco96972, w_eco96973, w_eco96974, w_eco96975, w_eco96976, w_eco96977, w_eco96978, w_eco96979, w_eco96980, w_eco96981, w_eco96982, w_eco96983, w_eco96984, w_eco96985, w_eco96986, w_eco96987, w_eco96988, w_eco96989, w_eco96990, w_eco96991, w_eco96992, w_eco96993, w_eco96994, w_eco96995, w_eco96996, w_eco96997, w_eco96998, w_eco96999, w_eco97000, w_eco97001, w_eco97002, w_eco97003, w_eco97004, w_eco97005, w_eco97006, w_eco97007, w_eco97008, w_eco97009, w_eco97010, w_eco97011, w_eco97012, w_eco97013, w_eco97014, w_eco97015, w_eco97016, w_eco97017, w_eco97018, w_eco97019, w_eco97020, w_eco97021, w_eco97022, w_eco97023, w_eco97024, w_eco97025, w_eco97026, w_eco97027, w_eco97028, w_eco97029, w_eco97030, w_eco97031, w_eco97032, w_eco97033, w_eco97034, w_eco97035, w_eco97036, w_eco97037, w_eco97038, w_eco97039, w_eco97040, w_eco97041, w_eco97042, w_eco97043, w_eco97044, w_eco97045, w_eco97046, w_eco97047, w_eco97048, w_eco97049, w_eco97050, w_eco97051, w_eco97052, w_eco97053, w_eco97054, w_eco97055, w_eco97056, w_eco97057, w_eco97058, w_eco97059, w_eco97060, w_eco97061, w_eco97062, w_eco97063, w_eco97064, w_eco97065, w_eco97066, w_eco97067, w_eco97068, w_eco97069, w_eco97070, w_eco97071, w_eco97072, w_eco97073, w_eco97074, w_eco97075, w_eco97076, w_eco97077, w_eco97078, w_eco97079, w_eco97080, w_eco97081, w_eco97082, w_eco97083, w_eco97084, w_eco97085, w_eco97086, w_eco97087, w_eco97088, w_eco97089, w_eco97090, w_eco97091, w_eco97092, w_eco97093, w_eco97094, w_eco97095, w_eco97096, w_eco97097, w_eco97098, w_eco97099, w_eco97100, w_eco97101, w_eco97102, w_eco97103, w_eco97104, w_eco97105, w_eco97106, w_eco97107, w_eco97108, w_eco97109, w_eco97110, w_eco97111, w_eco97112, w_eco97113, w_eco97114, w_eco97115, w_eco97116, w_eco97117, w_eco97118, w_eco97119, w_eco97120, w_eco97121, w_eco97122, w_eco97123, w_eco97124, w_eco97125, w_eco97126, w_eco97127, w_eco97128, w_eco97129, w_eco97130, w_eco97131, w_eco97132, w_eco97133, w_eco97134, w_eco97135, w_eco97136, w_eco97137, w_eco97138, w_eco97139, w_eco97140, w_eco97141, w_eco97142, w_eco97143, w_eco97144, w_eco97145, w_eco97146, w_eco97147, w_eco97148, w_eco97149, w_eco97150, w_eco97151, w_eco97152, w_eco97153, w_eco97154, w_eco97155, w_eco97156, w_eco97157, w_eco97158, w_eco97159, w_eco97160, w_eco97161, w_eco97162, w_eco97163, w_eco97164, w_eco97165, w_eco97166, w_eco97167, w_eco97168, w_eco97169, w_eco97170, w_eco97171, w_eco97172, w_eco97173, w_eco97174, w_eco97175, w_eco97176, w_eco97177, w_eco97178, w_eco97179, w_eco97180, w_eco97181, w_eco97182, w_eco97183, w_eco97184, w_eco97185, w_eco97186, w_eco97187, w_eco97188, w_eco97189, w_eco97190, w_eco97191, w_eco97192, w_eco97193, w_eco97194, w_eco97195, w_eco97196, w_eco97197, w_eco97198, w_eco97199, w_eco97200, w_eco97201, w_eco97202, w_eco97203, w_eco97204, w_eco97205, w_eco97206, w_eco97207, w_eco97208, w_eco97209, w_eco97210, w_eco97211, w_eco97212, w_eco97213, w_eco97214, w_eco97215, w_eco97216, w_eco97217, w_eco97218, w_eco97219, w_eco97220, w_eco97221, w_eco97222, w_eco97223, w_eco97224, w_eco97225, w_eco97226, w_eco97227, w_eco97228, w_eco97229, w_eco97230, w_eco97231, w_eco97232, w_eco97233, w_eco97234, w_eco97235, w_eco97236, w_eco97237, w_eco97238, w_eco97239, w_eco97240, w_eco97241, w_eco97242, w_eco97243, w_eco97244, w_eco97245, w_eco97246, w_eco97247, w_eco97248, w_eco97249, w_eco97250, w_eco97251, w_eco97252, w_eco97253, w_eco97254, w_eco97255, w_eco97256, w_eco97257, w_eco97258, w_eco97259, w_eco97260, w_eco97261, w_eco97262, w_eco97263, w_eco97264, w_eco97265, w_eco97266, w_eco97267, w_eco97268, w_eco97269, w_eco97270, w_eco97271, w_eco97272, w_eco97273, w_eco97274, w_eco97275, w_eco97276, w_eco97277, w_eco97278, w_eco97279, w_eco97280, w_eco97281, w_eco97282, w_eco97283, w_eco97284, w_eco97285, w_eco97286, w_eco97287, w_eco97288, w_eco97289, w_eco97290, w_eco97291, w_eco97292, w_eco97293, w_eco97294, w_eco97295, w_eco97296, w_eco97297, w_eco97298, w_eco97299, w_eco97300, w_eco97301, w_eco97302, w_eco97303, w_eco97304, w_eco97305, w_eco97306, w_eco97307, w_eco97308, w_eco97309, w_eco97310, w_eco97311, w_eco97312, w_eco97313, w_eco97314, w_eco97315, w_eco97316, w_eco97317, w_eco97318, w_eco97319, w_eco97320, w_eco97321, w_eco97322, w_eco97323, w_eco97324, w_eco97325, w_eco97326, w_eco97327, w_eco97328, w_eco97329, w_eco97330, w_eco97331, w_eco97332, w_eco97333, w_eco97334, w_eco97335, w_eco97336, w_eco97337, w_eco97338, w_eco97339, w_eco97340, w_eco97341, w_eco97342, w_eco97343, w_eco97344, w_eco97345, w_eco97346, w_eco97347, w_eco97348, w_eco97349, w_eco97350, w_eco97351, w_eco97352, w_eco97353, w_eco97354, w_eco97355, w_eco97356, w_eco97357, w_eco97358, w_eco97359, w_eco97360, w_eco97361, w_eco97362, w_eco97363, w_eco97364, w_eco97365, w_eco97366, w_eco97367, w_eco97368, w_eco97369, w_eco97370, w_eco97371, w_eco97372, w_eco97373, w_eco97374, w_eco97375, w_eco97376, w_eco97377, w_eco97378, w_eco97379, w_eco97380, w_eco97381, w_eco97382, w_eco97383, w_eco97384, w_eco97385, w_eco97386, w_eco97387, w_eco97388, w_eco97389, w_eco97390, w_eco97391, w_eco97392, w_eco97393, w_eco97394, w_eco97395, w_eco97396, w_eco97397, w_eco97398, w_eco97399, w_eco97400, w_eco97401, w_eco97402, w_eco97403, w_eco97404, w_eco97405, w_eco97406, w_eco97407, w_eco97408, w_eco97409, w_eco97410, w_eco97411, w_eco97412, w_eco97413, w_eco97414, w_eco97415, w_eco97416, w_eco97417, w_eco97418, w_eco97419, w_eco97420, w_eco97421, w_eco97422, w_eco97423, w_eco97424, w_eco97425, w_eco97426, w_eco97427, w_eco97428, w_eco97429, w_eco97430, w_eco97431, w_eco97432, w_eco97433, w_eco97434, w_eco97435, w_eco97436, w_eco97437, w_eco97438, w_eco97439, w_eco97440, w_eco97441, w_eco97442, w_eco97443, w_eco97444, w_eco97445, w_eco97446, w_eco97447, w_eco97448, w_eco97449, w_eco97450, w_eco97451, w_eco97452, w_eco97453, w_eco97454, w_eco97455, w_eco97456, w_eco97457, w_eco97458, w_eco97459, w_eco97460, w_eco97461, w_eco97462, w_eco97463, w_eco97464, w_eco97465, w_eco97466, w_eco97467, w_eco97468, w_eco97469, w_eco97470, w_eco97471, w_eco97472, w_eco97473, w_eco97474, w_eco97475, w_eco97476, w_eco97477, w_eco97478, w_eco97479, w_eco97480, w_eco97481, w_eco97482, w_eco97483, w_eco97484, w_eco97485, w_eco97486, w_eco97487, w_eco97488, w_eco97489, w_eco97490, w_eco97491, w_eco97492, w_eco97493, w_eco97494, w_eco97495, w_eco97496, w_eco97497, w_eco97498, w_eco97499, w_eco97500, w_eco97501, w_eco97502, w_eco97503, w_eco97504, w_eco97505, w_eco97506, w_eco97507, w_eco97508, w_eco97509, w_eco97510, w_eco97511, w_eco97512, w_eco97513, w_eco97514, w_eco97515, w_eco97516, w_eco97517, w_eco97518, w_eco97519, w_eco97520, w_eco97521, w_eco97522, w_eco97523, w_eco97524, w_eco97525, w_eco97526, w_eco97527, w_eco97528, w_eco97529, w_eco97530, w_eco97531, w_eco97532, w_eco97533, w_eco97534, w_eco97535, w_eco97536, w_eco97537, w_eco97538, w_eco97539, w_eco97540, w_eco97541, w_eco97542, w_eco97543, w_eco97544, w_eco97545, w_eco97546, w_eco97547, w_eco97548, w_eco97549, w_eco97550, w_eco97551, w_eco97552, w_eco97553, w_eco97554, w_eco97555, w_eco97556, w_eco97557, w_eco97558, w_eco97559, w_eco97560, w_eco97561, w_eco97562, w_eco97563, w_eco97564, w_eco97565, w_eco97566, w_eco97567, w_eco97568, w_eco97569, w_eco97570, w_eco97571, w_eco97572, w_eco97573, w_eco97574, w_eco97575, w_eco97576, w_eco97577, w_eco97578, w_eco97579, w_eco97580, w_eco97581, w_eco97582, w_eco97583, w_eco97584, w_eco97585, w_eco97586, w_eco97587, w_eco97588, w_eco97589, w_eco97590, w_eco97591, w_eco97592, w_eco97593, w_eco97594, w_eco97595, w_eco97596, w_eco97597, w_eco97598, w_eco97599, w_eco97600, w_eco97601, w_eco97602, w_eco97603, w_eco97604, w_eco97605, w_eco97606, w_eco97607, w_eco97608, w_eco97609, w_eco97610, w_eco97611, w_eco97612, w_eco97613, w_eco97614, w_eco97615, w_eco97616, w_eco97617, w_eco97618, w_eco97619, w_eco97620, w_eco97621, w_eco97622, w_eco97623, w_eco97624, w_eco97625, w_eco97626, w_eco97627, w_eco97628, w_eco97629, w_eco97630, w_eco97631, w_eco97632, w_eco97633, w_eco97634, w_eco97635, w_eco97636, w_eco97637, w_eco97638, w_eco97639, w_eco97640, w_eco97641, w_eco97642, w_eco97643, w_eco97644, w_eco97645, w_eco97646, w_eco97647, w_eco97648, w_eco97649, w_eco97650, w_eco97651, w_eco97652, w_eco97653, w_eco97654, w_eco97655, w_eco97656, w_eco97657, w_eco97658, w_eco97659, w_eco97660, w_eco97661, w_eco97662, w_eco97663, w_eco97664, w_eco97665, w_eco97666, w_eco97667, w_eco97668, w_eco97669, w_eco97670, w_eco97671, w_eco97672, w_eco97673, w_eco97674, w_eco97675, w_eco97676, w_eco97677, w_eco97678, w_eco97679, w_eco97680, w_eco97681, w_eco97682, w_eco97683, w_eco97684, w_eco97685, w_eco97686, w_eco97687, w_eco97688, w_eco97689, w_eco97690, w_eco97691, w_eco97692, w_eco97693, w_eco97694, w_eco97695, w_eco97696, w_eco97697, w_eco97698, w_eco97699, w_eco97700, w_eco97701, w_eco97702, w_eco97703, w_eco97704, w_eco97705, w_eco97706, w_eco97707, w_eco97708, w_eco97709, w_eco97710, w_eco97711, w_eco97712, w_eco97713, w_eco97714, w_eco97715, w_eco97716, w_eco97717, w_eco97718, w_eco97719, w_eco97720, w_eco97721, w_eco97722, w_eco97723, w_eco97724, w_eco97725, w_eco97726, w_eco97727, w_eco97728, w_eco97729, w_eco97730, w_eco97731, w_eco97732, w_eco97733, w_eco97734, w_eco97735, w_eco97736, w_eco97737, w_eco97738, w_eco97739, w_eco97740, w_eco97741, w_eco97742, w_eco97743, w_eco97744, w_eco97745, w_eco97746, w_eco97747, w_eco97748, w_eco97749, w_eco97750, w_eco97751, w_eco97752, w_eco97753, w_eco97754, w_eco97755, w_eco97756, w_eco97757, w_eco97758, w_eco97759, w_eco97760, w_eco97761, w_eco97762, w_eco97763, w_eco97764, w_eco97765, w_eco97766, w_eco97767, w_eco97768, w_eco97769, w_eco97770, w_eco97771, w_eco97772, w_eco97773, w_eco97774, w_eco97775, w_eco97776, w_eco97777, w_eco97778, w_eco97779, w_eco97780, w_eco97781, w_eco97782, w_eco97783, w_eco97784, w_eco97785, w_eco97786, w_eco97787, w_eco97788, w_eco97789, w_eco97790, w_eco97791, w_eco97792, w_eco97793, w_eco97794, w_eco97795, w_eco97796, w_eco97797, w_eco97798, w_eco97799, w_eco97800, w_eco97801, w_eco97802, w_eco97803, w_eco97804, w_eco97805, w_eco97806, w_eco97807, w_eco97808, w_eco97809, w_eco97810, w_eco97811, w_eco97812, w_eco97813, w_eco97814, w_eco97815, w_eco97816, w_eco97817, w_eco97818, w_eco97819, w_eco97820, w_eco97821, w_eco97822, w_eco97823, w_eco97824, w_eco97825, w_eco97826, w_eco97827, w_eco97828, w_eco97829, w_eco97830, w_eco97831, w_eco97832, w_eco97833, w_eco97834, w_eco97835, w_eco97836, w_eco97837, w_eco97838, w_eco97839, w_eco97840, w_eco97841, w_eco97842, w_eco97843, w_eco97844, w_eco97845, w_eco97846, w_eco97847, w_eco97848, w_eco97849, w_eco97850, w_eco97851, w_eco97852, w_eco97853, w_eco97854, w_eco97855, w_eco97856, w_eco97857, w_eco97858, w_eco97859, w_eco97860, w_eco97861, w_eco97862, w_eco97863, w_eco97864, w_eco97865, w_eco97866, w_eco97867, w_eco97868, w_eco97869, w_eco97870, w_eco97871, w_eco97872, w_eco97873, w_eco97874, w_eco97875, w_eco97876, w_eco97877, w_eco97878, w_eco97879, w_eco97880, w_eco97881, w_eco97882, w_eco97883, w_eco97884, w_eco97885, w_eco97886, w_eco97887, w_eco97888, w_eco97889, w_eco97890, w_eco97891, w_eco97892, w_eco97893, w_eco97894, w_eco97895, w_eco97896, w_eco97897, w_eco97898, w_eco97899, w_eco97900, w_eco97901, w_eco97902, w_eco97903, w_eco97904, w_eco97905, w_eco97906, w_eco97907, w_eco97908, w_eco97909, w_eco97910, w_eco97911, w_eco97912, w_eco97913, w_eco97914, w_eco97915, w_eco97916, w_eco97917, w_eco97918, w_eco97919, w_eco97920, w_eco97921, w_eco97922, w_eco97923, w_eco97924, w_eco97925, w_eco97926, w_eco97927, w_eco97928, w_eco97929, w_eco97930, w_eco97931, w_eco97932, w_eco97933, w_eco97934, w_eco97935, w_eco97936, w_eco97937, w_eco97938, w_eco97939, w_eco97940, w_eco97941, w_eco97942, w_eco97943, w_eco97944, w_eco97945, w_eco97946, w_eco97947, w_eco97948, w_eco97949, w_eco97950, w_eco97951, w_eco97952, w_eco97953, w_eco97954, w_eco97955, w_eco97956, w_eco97957, w_eco97958, w_eco97959, w_eco97960, w_eco97961, w_eco97962, w_eco97963, w_eco97964, w_eco97965, w_eco97966, w_eco97967, w_eco97968, w_eco97969, w_eco97970, w_eco97971, w_eco97972, w_eco97973, w_eco97974, w_eco97975, w_eco97976, w_eco97977, w_eco97978, w_eco97979, w_eco97980, w_eco97981, w_eco97982, w_eco97983, w_eco97984, w_eco97985, w_eco97986, w_eco97987, w_eco97988, w_eco97989, w_eco97990, w_eco97991, w_eco97992, w_eco97993, w_eco97994, w_eco97995, w_eco97996, w_eco97997, w_eco97998, w_eco97999, w_eco98000, w_eco98001, w_eco98002, w_eco98003, w_eco98004, w_eco98005, w_eco98006, w_eco98007, w_eco98008, w_eco98009, w_eco98010, w_eco98011, w_eco98012, w_eco98013, w_eco98014, w_eco98015, w_eco98016, w_eco98017, w_eco98018, w_eco98019, w_eco98020, w_eco98021, w_eco98022, w_eco98023, w_eco98024, w_eco98025, w_eco98026, w_eco98027, w_eco98028, w_eco98029, w_eco98030, w_eco98031, w_eco98032, w_eco98033, w_eco98034, w_eco98035, w_eco98036, w_eco98037, w_eco98038, w_eco98039, w_eco98040, w_eco98041, w_eco98042, w_eco98043, w_eco98044, w_eco98045, w_eco98046, w_eco98047, w_eco98048, w_eco98049, w_eco98050, w_eco98051, w_eco98052, w_eco98053, w_eco98054, w_eco98055, w_eco98056, w_eco98057, w_eco98058, w_eco98059, w_eco98060, w_eco98061, w_eco98062, w_eco98063, w_eco98064, w_eco98065, w_eco98066, w_eco98067, w_eco98068, w_eco98069, w_eco98070, w_eco98071, w_eco98072, w_eco98073, w_eco98074, w_eco98075, w_eco98076, w_eco98077, w_eco98078, w_eco98079, w_eco98080, w_eco98081, w_eco98082, w_eco98083, w_eco98084, w_eco98085, w_eco98086, w_eco98087, w_eco98088, w_eco98089, w_eco98090, w_eco98091, w_eco98092, w_eco98093, w_eco98094, w_eco98095, w_eco98096, w_eco98097, w_eco98098, w_eco98099, w_eco98100, w_eco98101, w_eco98102, w_eco98103, w_eco98104, w_eco98105, w_eco98106, w_eco98107, w_eco98108, w_eco98109, w_eco98110, w_eco98111, w_eco98112, w_eco98113, w_eco98114, w_eco98115, w_eco98116, w_eco98117, w_eco98118, w_eco98119, w_eco98120, w_eco98121, w_eco98122, w_eco98123, w_eco98124, w_eco98125, w_eco98126, w_eco98127, w_eco98128, w_eco98129, w_eco98130, w_eco98131, w_eco98132, w_eco98133, w_eco98134, w_eco98135, w_eco98136, w_eco98137, w_eco98138, w_eco98139, w_eco98140, w_eco98141, w_eco98142, w_eco98143, w_eco98144, w_eco98145, w_eco98146, w_eco98147, w_eco98148, w_eco98149, w_eco98150, w_eco98151, w_eco98152, w_eco98153, w_eco98154, w_eco98155, w_eco98156, w_eco98157, w_eco98158, w_eco98159, w_eco98160, w_eco98161, w_eco98162, w_eco98163, w_eco98164, w_eco98165, w_eco98166, w_eco98167, w_eco98168, w_eco98169, w_eco98170, w_eco98171, w_eco98172, w_eco98173, w_eco98174, w_eco98175, w_eco98176, w_eco98177, w_eco98178, w_eco98179, w_eco98180, w_eco98181, w_eco98182, w_eco98183, w_eco98184, w_eco98185, w_eco98186, w_eco98187, w_eco98188, w_eco98189, w_eco98190, w_eco98191, w_eco98192, w_eco98193, w_eco98194, w_eco98195, w_eco98196, w_eco98197, w_eco98198, w_eco98199, w_eco98200, w_eco98201, w_eco98202, w_eco98203, w_eco98204, w_eco98205, w_eco98206, w_eco98207, w_eco98208, w_eco98209, w_eco98210, w_eco98211, w_eco98212, w_eco98213, w_eco98214, w_eco98215, w_eco98216, w_eco98217, w_eco98218, w_eco98219, w_eco98220, w_eco98221, w_eco98222, w_eco98223, w_eco98224, w_eco98225, w_eco98226, w_eco98227, w_eco98228, w_eco98229, w_eco98230, w_eco98231, w_eco98232, w_eco98233, w_eco98234, w_eco98235, w_eco98236, w_eco98237, w_eco98238, w_eco98239, w_eco98240, w_eco98241, w_eco98242, w_eco98243, w_eco98244, w_eco98245, w_eco98246, w_eco98247, w_eco98248, w_eco98249, w_eco98250, w_eco98251, w_eco98252, w_eco98253, w_eco98254, w_eco98255, w_eco98256, w_eco98257, w_eco98258, w_eco98259, w_eco98260, w_eco98261, w_eco98262, w_eco98263, w_eco98264, w_eco98265, w_eco98266, w_eco98267, w_eco98268, w_eco98269, w_eco98270, w_eco98271, w_eco98272, w_eco98273, w_eco98274, w_eco98275, w_eco98276, w_eco98277, w_eco98278, w_eco98279, w_eco98280, w_eco98281, w_eco98282, w_eco98283, w_eco98284, w_eco98285, w_eco98286, w_eco98287, w_eco98288, w_eco98289, w_eco98290, w_eco98291, w_eco98292, w_eco98293, w_eco98294, w_eco98295, w_eco98296, w_eco98297, w_eco98298, w_eco98299, w_eco98300, w_eco98301, w_eco98302, w_eco98303, w_eco98304, w_eco98305, w_eco98306, w_eco98307, w_eco98308, w_eco98309, w_eco98310, w_eco98311, w_eco98312, w_eco98313, w_eco98314, w_eco98315, w_eco98316, w_eco98317, w_eco98318, w_eco98319, w_eco98320, w_eco98321, w_eco98322, w_eco98323, w_eco98324, w_eco98325, w_eco98326, w_eco98327, w_eco98328, w_eco98329, w_eco98330, w_eco98331, w_eco98332, w_eco98333, w_eco98334, w_eco98335, w_eco98336, w_eco98337, w_eco98338, w_eco98339, w_eco98340, w_eco98341, w_eco98342, w_eco98343, w_eco98344, w_eco98345, w_eco98346, w_eco98347, w_eco98348, w_eco98349, w_eco98350, w_eco98351, w_eco98352, w_eco98353, w_eco98354, w_eco98355, w_eco98356, w_eco98357, w_eco98358, w_eco98359, w_eco98360, w_eco98361, w_eco98362, w_eco98363, w_eco98364, w_eco98365, w_eco98366, w_eco98367, w_eco98368, w_eco98369, w_eco98370, w_eco98371, w_eco98372, w_eco98373, w_eco98374, w_eco98375, w_eco98376, w_eco98377, w_eco98378, w_eco98379, w_eco98380, w_eco98381, w_eco98382, w_eco98383, w_eco98384, w_eco98385, w_eco98386, w_eco98387, w_eco98388, w_eco98389, w_eco98390, w_eco98391, w_eco98392, w_eco98393, w_eco98394, w_eco98395, w_eco98396, w_eco98397, w_eco98398, w_eco98399, w_eco98400, w_eco98401, w_eco98402, w_eco98403, w_eco98404, w_eco98405, w_eco98406, w_eco98407, w_eco98408, w_eco98409, w_eco98410, w_eco98411, w_eco98412, w_eco98413, w_eco98414, w_eco98415, w_eco98416, w_eco98417, w_eco98418, w_eco98419, w_eco98420, w_eco98421, w_eco98422, w_eco98423, w_eco98424, w_eco98425, w_eco98426, w_eco98427, w_eco98428, w_eco98429, w_eco98430, w_eco98431, w_eco98432, w_eco98433, w_eco98434, w_eco98435, w_eco98436, w_eco98437, w_eco98438, w_eco98439, w_eco98440, w_eco98441, w_eco98442, w_eco98443, w_eco98444, w_eco98445, w_eco98446, w_eco98447, w_eco98448, w_eco98449, w_eco98450, w_eco98451, w_eco98452, w_eco98453, w_eco98454, w_eco98455, w_eco98456, w_eco98457, w_eco98458, w_eco98459, w_eco98460, w_eco98461, w_eco98462, w_eco98463, w_eco98464, w_eco98465, w_eco98466, w_eco98467, w_eco98468, w_eco98469, w_eco98470, w_eco98471, w_eco98472, w_eco98473, w_eco98474, w_eco98475, w_eco98476, w_eco98477, w_eco98478, w_eco98479, w_eco98480, w_eco98481, w_eco98482, w_eco98483, w_eco98484, w_eco98485, w_eco98486, w_eco98487, w_eco98488, w_eco98489, w_eco98490, w_eco98491, w_eco98492, w_eco98493, w_eco98494, w_eco98495, w_eco98496, w_eco98497, w_eco98498, w_eco98499, w_eco98500, w_eco98501, w_eco98502, w_eco98503, w_eco98504, w_eco98505, w_eco98506, w_eco98507, w_eco98508, w_eco98509, w_eco98510, w_eco98511, w_eco98512, w_eco98513, w_eco98514, w_eco98515, w_eco98516, w_eco98517, w_eco98518, w_eco98519, w_eco98520, w_eco98521, w_eco98522, w_eco98523, w_eco98524, w_eco98525, w_eco98526, w_eco98527, w_eco98528, w_eco98529, w_eco98530, w_eco98531, w_eco98532, w_eco98533, w_eco98534, w_eco98535, w_eco98536, w_eco98537, w_eco98538, w_eco98539, w_eco98540, w_eco98541, w_eco98542, w_eco98543, w_eco98544, w_eco98545, w_eco98546, w_eco98547, w_eco98548, w_eco98549, w_eco98550, w_eco98551, w_eco98552, w_eco98553, w_eco98554, w_eco98555, w_eco98556, w_eco98557, w_eco98558, w_eco98559, w_eco98560, w_eco98561, w_eco98562, w_eco98563, w_eco98564, w_eco98565, w_eco98566, w_eco98567, w_eco98568, w_eco98569, w_eco98570, w_eco98571, w_eco98572, w_eco98573, w_eco98574, w_eco98575, w_eco98576, w_eco98577, w_eco98578, w_eco98579, w_eco98580, w_eco98581, w_eco98582, w_eco98583, w_eco98584, w_eco98585, w_eco98586, w_eco98587, w_eco98588, w_eco98589, w_eco98590, w_eco98591, w_eco98592, w_eco98593, w_eco98594, w_eco98595, w_eco98596, w_eco98597, w_eco98598, w_eco98599, w_eco98600, w_eco98601, w_eco98602, w_eco98603, w_eco98604, w_eco98605, w_eco98606, w_eco98607, w_eco98608, w_eco98609, w_eco98610, w_eco98611, w_eco98612, w_eco98613, w_eco98614, w_eco98615, w_eco98616, w_eco98617, w_eco98618, w_eco98619, w_eco98620, w_eco98621, w_eco98622, w_eco98623, w_eco98624, w_eco98625, w_eco98626, w_eco98627, w_eco98628, w_eco98629, w_eco98630, w_eco98631, w_eco98632, w_eco98633, w_eco98634, w_eco98635, w_eco98636, w_eco98637, w_eco98638, w_eco98639, w_eco98640, w_eco98641, w_eco98642, w_eco98643, w_eco98644, w_eco98645, w_eco98646, w_eco98647, w_eco98648, w_eco98649, w_eco98650, w_eco98651, w_eco98652, w_eco98653, w_eco98654, w_eco98655, w_eco98656, w_eco98657, w_eco98658, w_eco98659, w_eco98660, w_eco98661, w_eco98662, w_eco98663, w_eco98664, w_eco98665, w_eco98666, w_eco98667, w_eco98668, w_eco98669, w_eco98670, w_eco98671, w_eco98672, w_eco98673, w_eco98674, w_eco98675, w_eco98676, w_eco98677, w_eco98678, w_eco98679, w_eco98680, w_eco98681, w_eco98682, w_eco98683, w_eco98684, w_eco98685, w_eco98686, w_eco98687, w_eco98688, w_eco98689, w_eco98690, w_eco98691, w_eco98692, w_eco98693, w_eco98694, w_eco98695, w_eco98696, w_eco98697, w_eco98698, w_eco98699, w_eco98700, w_eco98701, w_eco98702, w_eco98703, w_eco98704, w_eco98705, w_eco98706, w_eco98707, w_eco98708, w_eco98709, w_eco98710, w_eco98711, w_eco98712, w_eco98713, w_eco98714, w_eco98715, w_eco98716, w_eco98717, w_eco98718, w_eco98719, w_eco98720, w_eco98721, w_eco98722, w_eco98723, w_eco98724, w_eco98725, w_eco98726, w_eco98727, w_eco98728, w_eco98729, w_eco98730, w_eco98731, w_eco98732, w_eco98733, w_eco98734, w_eco98735, w_eco98736, w_eco98737, w_eco98738, w_eco98739, w_eco98740, w_eco98741, w_eco98742, w_eco98743, w_eco98744, w_eco98745, w_eco98746, w_eco98747, w_eco98748, w_eco98749, w_eco98750, w_eco98751, w_eco98752, w_eco98753, w_eco98754, w_eco98755, w_eco98756, w_eco98757, w_eco98758, w_eco98759, w_eco98760, w_eco98761, w_eco98762, w_eco98763, w_eco98764, w_eco98765, w_eco98766, w_eco98767, w_eco98768, w_eco98769, w_eco98770, w_eco98771, w_eco98772, w_eco98773, w_eco98774, w_eco98775, w_eco98776, w_eco98777, w_eco98778, w_eco98779, w_eco98780, w_eco98781, w_eco98782, w_eco98783, w_eco98784, w_eco98785, w_eco98786, w_eco98787, w_eco98788, w_eco98789, w_eco98790, w_eco98791, w_eco98792, w_eco98793, w_eco98794, w_eco98795, w_eco98796, w_eco98797, w_eco98798, w_eco98799, w_eco98800, w_eco98801, w_eco98802, w_eco98803, w_eco98804, w_eco98805, w_eco98806, w_eco98807, w_eco98808, w_eco98809, w_eco98810, w_eco98811, w_eco98812, w_eco98813, w_eco98814, w_eco98815, w_eco98816, w_eco98817, w_eco98818, w_eco98819, w_eco98820, w_eco98821, w_eco98822, w_eco98823, w_eco98824, w_eco98825, w_eco98826, w_eco98827, w_eco98828, w_eco98829, w_eco98830, w_eco98831, w_eco98832, w_eco98833, w_eco98834, w_eco98835, w_eco98836, w_eco98837, w_eco98838, w_eco98839, w_eco98840, w_eco98841, w_eco98842, w_eco98843, w_eco98844, w_eco98845, w_eco98846, w_eco98847, w_eco98848, w_eco98849, w_eco98850, w_eco98851, w_eco98852, w_eco98853, w_eco98854, w_eco98855, w_eco98856, w_eco98857, w_eco98858, w_eco98859, w_eco98860, w_eco98861, w_eco98862, w_eco98863, w_eco98864, w_eco98865, w_eco98866, w_eco98867, w_eco98868, w_eco98869, w_eco98870, w_eco98871, w_eco98872, w_eco98873, w_eco98874, w_eco98875, w_eco98876, w_eco98877, w_eco98878, w_eco98879, w_eco98880, w_eco98881, w_eco98882, w_eco98883, w_eco98884, w_eco98885, w_eco98886, w_eco98887, w_eco98888, w_eco98889, w_eco98890, w_eco98891, w_eco98892, w_eco98893, w_eco98894, w_eco98895, w_eco98896, w_eco98897, w_eco98898, w_eco98899, w_eco98900, w_eco98901, w_eco98902, w_eco98903, w_eco98904, w_eco98905, w_eco98906, w_eco98907, w_eco98908, w_eco98909, w_eco98910, w_eco98911, w_eco98912, w_eco98913, w_eco98914, w_eco98915, w_eco98916, w_eco98917, w_eco98918, w_eco98919, w_eco98920, w_eco98921, w_eco98922, w_eco98923, w_eco98924, w_eco98925, w_eco98926, w_eco98927, w_eco98928, w_eco98929, w_eco98930, w_eco98931, w_eco98932, w_eco98933, w_eco98934, w_eco98935, w_eco98936, w_eco98937, w_eco98938, w_eco98939, w_eco98940, w_eco98941, w_eco98942, w_eco98943, w_eco98944, w_eco98945, w_eco98946, w_eco98947, w_eco98948, w_eco98949, w_eco98950, w_eco98951, w_eco98952, w_eco98953, w_eco98954, w_eco98955, w_eco98956, w_eco98957, w_eco98958, w_eco98959, w_eco98960, w_eco98961, w_eco98962, w_eco98963, w_eco98964, w_eco98965, w_eco98966, w_eco98967, w_eco98968, w_eco98969, w_eco98970, w_eco98971, w_eco98972, w_eco98973, w_eco98974, w_eco98975, w_eco98976, w_eco98977, w_eco98978, w_eco98979, w_eco98980, w_eco98981, w_eco98982, w_eco98983, w_eco98984, w_eco98985, w_eco98986, w_eco98987, w_eco98988, w_eco98989, w_eco98990, w_eco98991, w_eco98992, w_eco98993, w_eco98994, w_eco98995, w_eco98996, w_eco98997, w_eco98998, w_eco98999, w_eco99000, w_eco99001, w_eco99002, w_eco99003, w_eco99004, w_eco99005, w_eco99006, w_eco99007, w_eco99008, w_eco99009, w_eco99010, w_eco99011, w_eco99012, w_eco99013, w_eco99014, w_eco99015, w_eco99016, w_eco99017, w_eco99018, w_eco99019, w_eco99020, w_eco99021, w_eco99022, w_eco99023, w_eco99024, w_eco99025, w_eco99026, w_eco99027, w_eco99028, w_eco99029, w_eco99030, w_eco99031, w_eco99032, w_eco99033, w_eco99034, w_eco99035, w_eco99036, w_eco99037, w_eco99038, w_eco99039, w_eco99040, w_eco99041, w_eco99042, w_eco99043, w_eco99044, w_eco99045, w_eco99046, w_eco99047, w_eco99048, w_eco99049, w_eco99050, w_eco99051, w_eco99052, w_eco99053, w_eco99054, w_eco99055, w_eco99056, w_eco99057, w_eco99058, w_eco99059, w_eco99060, w_eco99061, w_eco99062, w_eco99063, w_eco99064, w_eco99065, w_eco99066, w_eco99067, w_eco99068, w_eco99069, w_eco99070, w_eco99071, w_eco99072, w_eco99073, w_eco99074, w_eco99075, w_eco99076, w_eco99077, w_eco99078, w_eco99079, w_eco99080, w_eco99081, w_eco99082, w_eco99083, w_eco99084, w_eco99085, w_eco99086, w_eco99087, w_eco99088, w_eco99089, w_eco99090, w_eco99091, w_eco99092, w_eco99093, w_eco99094, w_eco99095, w_eco99096, w_eco99097, w_eco99098, w_eco99099, w_eco99100, w_eco99101, w_eco99102, w_eco99103, w_eco99104, w_eco99105, w_eco99106, w_eco99107, w_eco99108, w_eco99109, w_eco99110, w_eco99111, w_eco99112, w_eco99113, w_eco99114, w_eco99115, w_eco99116, w_eco99117, w_eco99118, w_eco99119, w_eco99120, w_eco99121, w_eco99122, w_eco99123, w_eco99124, w_eco99125, w_eco99126, w_eco99127, w_eco99128, w_eco99129, w_eco99130, w_eco99131, w_eco99132, w_eco99133, w_eco99134, w_eco99135, w_eco99136, w_eco99137, w_eco99138, w_eco99139, w_eco99140, w_eco99141, w_eco99142, w_eco99143, w_eco99144, w_eco99145, w_eco99146, w_eco99147, w_eco99148, w_eco99149, w_eco99150, w_eco99151, w_eco99152, w_eco99153, w_eco99154, w_eco99155, w_eco99156, w_eco99157, w_eco99158, w_eco99159, w_eco99160, w_eco99161, w_eco99162, w_eco99163, w_eco99164, w_eco99165, w_eco99166, w_eco99167, w_eco99168, w_eco99169, w_eco99170, w_eco99171, w_eco99172, w_eco99173, w_eco99174, w_eco99175, w_eco99176, w_eco99177, w_eco99178, w_eco99179, w_eco99180, w_eco99181, w_eco99182, w_eco99183, w_eco99184, w_eco99185, w_eco99186, w_eco99187, w_eco99188, w_eco99189, w_eco99190, w_eco99191, w_eco99192, w_eco99193, w_eco99194, w_eco99195, w_eco99196, w_eco99197, w_eco99198, w_eco99199, w_eco99200, w_eco99201, w_eco99202, w_eco99203, w_eco99204, w_eco99205, w_eco99206, w_eco99207, w_eco99208, w_eco99209, w_eco99210, w_eco99211, w_eco99212, w_eco99213, w_eco99214, w_eco99215, w_eco99216, w_eco99217, w_eco99218, w_eco99219, w_eco99220, w_eco99221, w_eco99222, w_eco99223, w_eco99224, w_eco99225, w_eco99226, w_eco99227, w_eco99228, w_eco99229, w_eco99230, w_eco99231, w_eco99232, w_eco99233, w_eco99234, w_eco99235, w_eco99236, w_eco99237, w_eco99238, w_eco99239, w_eco99240, w_eco99241, w_eco99242, w_eco99243, w_eco99244, w_eco99245, w_eco99246, w_eco99247, w_eco99248, w_eco99249, w_eco99250, w_eco99251, w_eco99252, w_eco99253, w_eco99254, w_eco99255, w_eco99256, w_eco99257, w_eco99258, w_eco99259, w_eco99260, w_eco99261, w_eco99262, w_eco99263, w_eco99264, w_eco99265, w_eco99266, w_eco99267, w_eco99268, w_eco99269, w_eco99270, w_eco99271, w_eco99272, w_eco99273, w_eco99274, w_eco99275, w_eco99276, w_eco99277, w_eco99278, w_eco99279, w_eco99280, w_eco99281, w_eco99282, w_eco99283, w_eco99284, w_eco99285, w_eco99286, w_eco99287, w_eco99288, w_eco99289, w_eco99290, w_eco99291, w_eco99292, w_eco99293, w_eco99294, w_eco99295, w_eco99296, w_eco99297, w_eco99298, w_eco99299, w_eco99300, w_eco99301, w_eco99302, w_eco99303, w_eco99304, w_eco99305, w_eco99306, w_eco99307, w_eco99308, w_eco99309, w_eco99310, w_eco99311, w_eco99312, w_eco99313, w_eco99314, w_eco99315, w_eco99316, w_eco99317, w_eco99318, w_eco99319, w_eco99320, w_eco99321, w_eco99322, w_eco99323, w_eco99324, w_eco99325, w_eco99326, w_eco99327, w_eco99328, w_eco99329, w_eco99330, w_eco99331, w_eco99332, w_eco99333, w_eco99334, w_eco99335, w_eco99336, w_eco99337, w_eco99338, w_eco99339, w_eco99340, w_eco99341, w_eco99342, w_eco99343, w_eco99344, w_eco99345, w_eco99346, w_eco99347, w_eco99348, w_eco99349, w_eco99350, w_eco99351, w_eco99352, w_eco99353, w_eco99354, w_eco99355, w_eco99356, w_eco99357, w_eco99358, w_eco99359, w_eco99360, w_eco99361, w_eco99362, w_eco99363, w_eco99364, w_eco99365, w_eco99366, w_eco99367, w_eco99368, w_eco99369, w_eco99370, w_eco99371, w_eco99372, w_eco99373, w_eco99374, w_eco99375, w_eco99376, w_eco99377, w_eco99378, w_eco99379, w_eco99380, w_eco99381, w_eco99382, w_eco99383, w_eco99384, w_eco99385, w_eco99386, w_eco99387, w_eco99388, w_eco99389, w_eco99390, w_eco99391, w_eco99392, w_eco99393, w_eco99394, w_eco99395, w_eco99396, w_eco99397, w_eco99398, w_eco99399, w_eco99400, w_eco99401, w_eco99402, w_eco99403, w_eco99404, w_eco99405, w_eco99406, w_eco99407, w_eco99408, w_eco99409, w_eco99410, w_eco99411, w_eco99412, w_eco99413, w_eco99414, w_eco99415, w_eco99416, w_eco99417, w_eco99418, w_eco99419, w_eco99420, w_eco99421, w_eco99422, w_eco99423, w_eco99424, w_eco99425, w_eco99426, w_eco99427, w_eco99428, w_eco99429, w_eco99430, w_eco99431, w_eco99432, w_eco99433, w_eco99434, w_eco99435, w_eco99436, w_eco99437, w_eco99438, w_eco99439, w_eco99440, w_eco99441, w_eco99442, w_eco99443, w_eco99444, w_eco99445, w_eco99446, w_eco99447, w_eco99448, w_eco99449, w_eco99450, w_eco99451, w_eco99452, w_eco99453, w_eco99454, w_eco99455, w_eco99456, w_eco99457, w_eco99458, w_eco99459, w_eco99460, w_eco99461, w_eco99462, w_eco99463, w_eco99464, w_eco99465, w_eco99466, w_eco99467, w_eco99468, w_eco99469, w_eco99470, w_eco99471, w_eco99472, w_eco99473, w_eco99474, w_eco99475, w_eco99476, w_eco99477, w_eco99478, w_eco99479, w_eco99480, w_eco99481, w_eco99482, w_eco99483, w_eco99484, w_eco99485, w_eco99486, w_eco99487, w_eco99488, w_eco99489, w_eco99490, w_eco99491, w_eco99492, w_eco99493, w_eco99494, w_eco99495, w_eco99496, w_eco99497, w_eco99498, w_eco99499, w_eco99500, w_eco99501, w_eco99502, w_eco99503, w_eco99504, w_eco99505, w_eco99506, w_eco99507, w_eco99508, w_eco99509, w_eco99510, w_eco99511, w_eco99512, w_eco99513, w_eco99514, w_eco99515, w_eco99516, w_eco99517, w_eco99518, w_eco99519, w_eco99520, w_eco99521, w_eco99522, w_eco99523, w_eco99524, w_eco99525, w_eco99526, w_eco99527, w_eco99528, w_eco99529, w_eco99530, w_eco99531, w_eco99532, w_eco99533, w_eco99534, w_eco99535, w_eco99536, w_eco99537, w_eco99538, w_eco99539, w_eco99540, w_eco99541, w_eco99542, w_eco99543, w_eco99544, w_eco99545, w_eco99546, w_eco99547, w_eco99548, w_eco99549, w_eco99550, w_eco99551, w_eco99552, w_eco99553, w_eco99554, w_eco99555, w_eco99556, w_eco99557, w_eco99558, w_eco99559, w_eco99560, w_eco99561, w_eco99562, w_eco99563, w_eco99564, w_eco99565, w_eco99566, w_eco99567, w_eco99568, w_eco99569, w_eco99570, w_eco99571, w_eco99572, w_eco99573, w_eco99574, w_eco99575, w_eco99576, w_eco99577, w_eco99578, w_eco99579, w_eco99580, w_eco99581, w_eco99582, w_eco99583, w_eco99584, w_eco99585, w_eco99586, w_eco99587, w_eco99588, w_eco99589, w_eco99590, w_eco99591, w_eco99592, w_eco99593, w_eco99594, w_eco99595, w_eco99596, w_eco99597, w_eco99598, w_eco99599, w_eco99600, w_eco99601, w_eco99602, w_eco99603, w_eco99604, w_eco99605, w_eco99606, w_eco99607, w_eco99608, w_eco99609, w_eco99610, w_eco99611, w_eco99612, w_eco99613, w_eco99614, w_eco99615, w_eco99616, w_eco99617, w_eco99618, w_eco99619, w_eco99620, w_eco99621, w_eco99622, w_eco99623, w_eco99624, w_eco99625, w_eco99626, w_eco99627, w_eco99628, w_eco99629, w_eco99630, w_eco99631, w_eco99632, w_eco99633, w_eco99634, w_eco99635, w_eco99636, w_eco99637, w_eco99638, w_eco99639, w_eco99640, w_eco99641, w_eco99642, w_eco99643, w_eco99644, w_eco99645, w_eco99646, w_eco99647, w_eco99648, w_eco99649, w_eco99650, w_eco99651, w_eco99652, w_eco99653, w_eco99654, w_eco99655, w_eco99656, w_eco99657, w_eco99658, w_eco99659, w_eco99660, w_eco99661, w_eco99662, w_eco99663, w_eco99664, w_eco99665, w_eco99666, w_eco99667, w_eco99668, w_eco99669, w_eco99670, w_eco99671, w_eco99672, w_eco99673, w_eco99674, w_eco99675, w_eco99676, w_eco99677, w_eco99678, w_eco99679, w_eco99680, w_eco99681, w_eco99682, w_eco99683, w_eco99684, w_eco99685, w_eco99686, w_eco99687, w_eco99688, w_eco99689, w_eco99690, w_eco99691, w_eco99692, w_eco99693, w_eco99694, w_eco99695, w_eco99696, w_eco99697, w_eco99698, w_eco99699, w_eco99700, w_eco99701, w_eco99702, w_eco99703, w_eco99704, w_eco99705, w_eco99706, w_eco99707, w_eco99708, w_eco99709, w_eco99710, w_eco99711, w_eco99712, w_eco99713, w_eco99714, w_eco99715, w_eco99716, w_eco99717, w_eco99718, w_eco99719, w_eco99720, w_eco99721, w_eco99722, w_eco99723, w_eco99724, w_eco99725, w_eco99726, w_eco99727, w_eco99728, w_eco99729, w_eco99730, w_eco99731, w_eco99732, w_eco99733, w_eco99734, w_eco99735, w_eco99736, w_eco99737, w_eco99738, w_eco99739, w_eco99740, w_eco99741, w_eco99742, w_eco99743, w_eco99744, w_eco99745, w_eco99746, w_eco99747, w_eco99748, w_eco99749, w_eco99750, w_eco99751, w_eco99752, w_eco99753, w_eco99754, w_eco99755, w_eco99756, w_eco99757, w_eco99758, w_eco99759, w_eco99760, w_eco99761, w_eco99762, w_eco99763, w_eco99764, w_eco99765, w_eco99766, w_eco99767, w_eco99768, w_eco99769, w_eco99770, w_eco99771, w_eco99772, w_eco99773, w_eco99774, w_eco99775, w_eco99776, w_eco99777, w_eco99778, w_eco99779, w_eco99780, w_eco99781, w_eco99782, w_eco99783, w_eco99784, w_eco99785, w_eco99786, w_eco99787, w_eco99788, w_eco99789, w_eco99790, w_eco99791, w_eco99792, w_eco99793, w_eco99794, w_eco99795, w_eco99796, w_eco99797, w_eco99798, w_eco99799, w_eco99800, w_eco99801, w_eco99802, w_eco99803, w_eco99804, w_eco99805, w_eco99806, w_eco99807, w_eco99808, w_eco99809, w_eco99810, w_eco99811, w_eco99812, w_eco99813, w_eco99814, w_eco99815, w_eco99816, w_eco99817, w_eco99818, w_eco99819, w_eco99820, w_eco99821, w_eco99822, w_eco99823, w_eco99824, w_eco99825, w_eco99826, w_eco99827, w_eco99828, w_eco99829, w_eco99830, w_eco99831, w_eco99832, w_eco99833, w_eco99834, w_eco99835, w_eco99836, w_eco99837, w_eco99838, w_eco99839, w_eco99840, w_eco99841, w_eco99842, w_eco99843, w_eco99844, w_eco99845, w_eco99846, w_eco99847, w_eco99848, w_eco99849, w_eco99850, w_eco99851, w_eco99852, w_eco99853, w_eco99854, w_eco99855, w_eco99856, w_eco99857, w_eco99858, w_eco99859, w_eco99860, w_eco99861, w_eco99862, w_eco99863, w_eco99864, w_eco99865, w_eco99866, w_eco99867, w_eco99868, w_eco99869, w_eco99870, w_eco99871, w_eco99872, w_eco99873, w_eco99874, w_eco99875, w_eco99876, w_eco99877, w_eco99878, w_eco99879, w_eco99880, w_eco99881, w_eco99882, w_eco99883, w_eco99884, w_eco99885, w_eco99886, w_eco99887, w_eco99888, w_eco99889, w_eco99890, w_eco99891, w_eco99892, w_eco99893, w_eco99894, w_eco99895, w_eco99896, w_eco99897, w_eco99898, w_eco99899, w_eco99900, w_eco99901, w_eco99902, w_eco99903, w_eco99904, w_eco99905, w_eco99906, w_eco99907, w_eco99908, w_eco99909, w_eco99910, w_eco99911, w_eco99912, w_eco99913, w_eco99914, w_eco99915, w_eco99916, w_eco99917, w_eco99918, w_eco99919, w_eco99920, w_eco99921, w_eco99922, w_eco99923, w_eco99924, w_eco99925, w_eco99926, w_eco99927, w_eco99928, w_eco99929, w_eco99930, w_eco99931, w_eco99932, w_eco99933, w_eco99934, w_eco99935, w_eco99936, w_eco99937, w_eco99938, w_eco99939, w_eco99940, w_eco99941, w_eco99942, w_eco99943, w_eco99944, w_eco99945, w_eco99946, w_eco99947, w_eco99948, w_eco99949, w_eco99950, w_eco99951, w_eco99952, w_eco99953, w_eco99954, w_eco99955, w_eco99956, w_eco99957, w_eco99958, w_eco99959, w_eco99960, w_eco99961, w_eco99962, w_eco99963, w_eco99964, w_eco99965, w_eco99966, w_eco99967, w_eco99968, w_eco99969, w_eco99970, w_eco99971, w_eco99972, w_eco99973, w_eco99974, w_eco99975, w_eco99976, w_eco99977, w_eco99978, w_eco99979, w_eco99980, w_eco99981, w_eco99982, w_eco99983, w_eco99984, w_eco99985, w_eco99986, w_eco99987, w_eco99988, w_eco99989, w_eco99990, w_eco99991, w_eco99992, w_eco99993, w_eco99994, w_eco99995, w_eco99996, w_eco99997, w_eco99998, w_eco99999, w_eco100000, w_eco100001, w_eco100002, w_eco100003, w_eco100004, w_eco100005, w_eco100006, w_eco100007, w_eco100008, w_eco100009, w_eco100010, w_eco100011, w_eco100012, w_eco100013, w_eco100014, w_eco100015, w_eco100016, w_eco100017, w_eco100018, w_eco100019, w_eco100020, w_eco100021, w_eco100022, w_eco100023, w_eco100024, w_eco100025, w_eco100026, w_eco100027, w_eco100028, w_eco100029, w_eco100030, w_eco100031, w_eco100032, w_eco100033, w_eco100034, w_eco100035, w_eco100036, w_eco100037, w_eco100038, w_eco100039, w_eco100040, w_eco100041, w_eco100042, w_eco100043, w_eco100044, w_eco100045, w_eco100046, w_eco100047, w_eco100048, w_eco100049, w_eco100050, w_eco100051, w_eco100052, w_eco100053, w_eco100054, w_eco100055, w_eco100056, w_eco100057, w_eco100058, w_eco100059, w_eco100060, w_eco100061, w_eco100062, w_eco100063, w_eco100064, w_eco100065, w_eco100066, w_eco100067, w_eco100068, w_eco100069, w_eco100070, w_eco100071, w_eco100072, w_eco100073, w_eco100074, w_eco100075, w_eco100076, w_eco100077, w_eco100078, w_eco100079, w_eco100080, w_eco100081, w_eco100082, w_eco100083, w_eco100084, w_eco100085, w_eco100086, w_eco100087, w_eco100088, w_eco100089, w_eco100090, w_eco100091, w_eco100092, w_eco100093, w_eco100094, w_eco100095, w_eco100096, w_eco100097, w_eco100098, w_eco100099, w_eco100100, w_eco100101, w_eco100102, w_eco100103, w_eco100104, w_eco100105, w_eco100106, w_eco100107, w_eco100108, w_eco100109, w_eco100110, w_eco100111, w_eco100112, w_eco100113, w_eco100114, w_eco100115, w_eco100116, w_eco100117, w_eco100118, w_eco100119, w_eco100120, w_eco100121, w_eco100122, w_eco100123, w_eco100124, w_eco100125, w_eco100126, w_eco100127, w_eco100128, w_eco100129, w_eco100130, w_eco100131, w_eco100132, w_eco100133, w_eco100134, w_eco100135, w_eco100136, w_eco100137, w_eco100138, w_eco100139, w_eco100140, w_eco100141, w_eco100142, w_eco100143, w_eco100144, w_eco100145, w_eco100146, w_eco100147, w_eco100148, w_eco100149, w_eco100150, w_eco100151, w_eco100152, w_eco100153, w_eco100154, w_eco100155, w_eco100156, w_eco100157, w_eco100158, w_eco100159, w_eco100160, w_eco100161, w_eco100162, w_eco100163, w_eco100164, w_eco100165, w_eco100166, w_eco100167, w_eco100168, w_eco100169, w_eco100170, w_eco100171, w_eco100172, w_eco100173, w_eco100174, w_eco100175, w_eco100176, w_eco100177, w_eco100178, w_eco100179, w_eco100180, w_eco100181, w_eco100182, w_eco100183, w_eco100184, w_eco100185, w_eco100186, w_eco100187, w_eco100188, w_eco100189, w_eco100190, w_eco100191, w_eco100192, w_eco100193, w_eco100194, w_eco100195, w_eco100196, w_eco100197, w_eco100198, w_eco100199, w_eco100200, w_eco100201, w_eco100202, w_eco100203, w_eco100204, w_eco100205, w_eco100206, w_eco100207, w_eco100208, w_eco100209, w_eco100210, w_eco100211, w_eco100212, w_eco100213, w_eco100214, w_eco100215, w_eco100216, w_eco100217, w_eco100218, w_eco100219, w_eco100220, w_eco100221, w_eco100222, w_eco100223, w_eco100224, w_eco100225, w_eco100226, w_eco100227, w_eco100228, w_eco100229, w_eco100230, w_eco100231, w_eco100232, w_eco100233, w_eco100234, w_eco100235, w_eco100236, w_eco100237, w_eco100238, w_eco100239, w_eco100240, w_eco100241, w_eco100242, w_eco100243, w_eco100244, w_eco100245, w_eco100246, w_eco100247, w_eco100248, w_eco100249, w_eco100250, w_eco100251, w_eco100252, w_eco100253, w_eco100254, w_eco100255, w_eco100256, w_eco100257, w_eco100258, w_eco100259, w_eco100260, w_eco100261, w_eco100262, w_eco100263, w_eco100264, w_eco100265, w_eco100266, w_eco100267, w_eco100268, w_eco100269, w_eco100270, w_eco100271, w_eco100272, w_eco100273, w_eco100274, w_eco100275, w_eco100276, w_eco100277, w_eco100278, w_eco100279, w_eco100280, w_eco100281, w_eco100282, w_eco100283, w_eco100284, w_eco100285, w_eco100286, w_eco100287, w_eco100288, w_eco100289, w_eco100290, w_eco100291, w_eco100292, w_eco100293, w_eco100294, w_eco100295, w_eco100296, w_eco100297, w_eco100298, w_eco100299, w_eco100300, w_eco100301, w_eco100302, w_eco100303, w_eco100304, w_eco100305, w_eco100306, w_eco100307, w_eco100308, w_eco100309, w_eco100310, w_eco100311, w_eco100312, w_eco100313, w_eco100314, w_eco100315, w_eco100316, w_eco100317, w_eco100318, w_eco100319, w_eco100320, w_eco100321, w_eco100322, w_eco100323, w_eco100324, w_eco100325, w_eco100326, w_eco100327, w_eco100328, w_eco100329, w_eco100330, w_eco100331, w_eco100332, w_eco100333, w_eco100334, w_eco100335, w_eco100336, w_eco100337, w_eco100338, w_eco100339, w_eco100340, w_eco100341, w_eco100342, w_eco100343, w_eco100344, w_eco100345, w_eco100346, w_eco100347, w_eco100348, w_eco100349, w_eco100350, w_eco100351, w_eco100352, w_eco100353, w_eco100354, w_eco100355, w_eco100356, w_eco100357, w_eco100358, w_eco100359, w_eco100360, w_eco100361, w_eco100362, w_eco100363, w_eco100364, w_eco100365, w_eco100366, w_eco100367, w_eco100368, w_eco100369, w_eco100370, w_eco100371, w_eco100372, w_eco100373, w_eco100374, w_eco100375, w_eco100376, w_eco100377, w_eco100378, w_eco100379, w_eco100380, w_eco100381, w_eco100382, w_eco100383, w_eco100384, w_eco100385, w_eco100386, w_eco100387, w_eco100388, w_eco100389, w_eco100390, w_eco100391, w_eco100392, w_eco100393, w_eco100394, w_eco100395, w_eco100396, w_eco100397, w_eco100398, w_eco100399, w_eco100400, w_eco100401, w_eco100402, w_eco100403, w_eco100404, w_eco100405, w_eco100406, w_eco100407, w_eco100408, w_eco100409, w_eco100410, w_eco100411, w_eco100412, w_eco100413, w_eco100414, w_eco100415, w_eco100416, w_eco100417, w_eco100418, w_eco100419, w_eco100420, w_eco100421, w_eco100422, w_eco100423, w_eco100424, w_eco100425, w_eco100426, w_eco100427, w_eco100428, w_eco100429, w_eco100430, w_eco100431, w_eco100432, w_eco100433, w_eco100434, w_eco100435, w_eco100436, w_eco100437, w_eco100438, w_eco100439, w_eco100440, w_eco100441, w_eco100442, w_eco100443, w_eco100444, w_eco100445, w_eco100446, w_eco100447, w_eco100448, w_eco100449, w_eco100450, w_eco100451, w_eco100452, w_eco100453, w_eco100454, w_eco100455, w_eco100456, w_eco100457, w_eco100458, w_eco100459, w_eco100460, w_eco100461, w_eco100462, w_eco100463, w_eco100464, w_eco100465, w_eco100466, w_eco100467, w_eco100468, w_eco100469, w_eco100470, w_eco100471, w_eco100472, w_eco100473, w_eco100474, w_eco100475, w_eco100476, w_eco100477, w_eco100478, w_eco100479, w_eco100480, w_eco100481, w_eco100482, w_eco100483, w_eco100484, w_eco100485, w_eco100486, w_eco100487, w_eco100488, w_eco100489, w_eco100490, w_eco100491, w_eco100492, w_eco100493, w_eco100494, w_eco100495, w_eco100496, w_eco100497, w_eco100498, w_eco100499, w_eco100500, w_eco100501, w_eco100502, w_eco100503, w_eco100504, w_eco100505, w_eco100506, w_eco100507, w_eco100508, w_eco100509, w_eco100510, w_eco100511, w_eco100512, w_eco100513, w_eco100514, w_eco100515, w_eco100516, w_eco100517, w_eco100518, w_eco100519, w_eco100520, w_eco100521, w_eco100522, w_eco100523, w_eco100524, w_eco100525, w_eco100526, w_eco100527, w_eco100528, w_eco100529, w_eco100530, w_eco100531, w_eco100532, w_eco100533, w_eco100534, w_eco100535, w_eco100536, w_eco100537, w_eco100538, w_eco100539, w_eco100540, w_eco100541, w_eco100542, w_eco100543, w_eco100544, w_eco100545, w_eco100546, w_eco100547, w_eco100548, w_eco100549, w_eco100550, w_eco100551, w_eco100552, w_eco100553, w_eco100554, w_eco100555, w_eco100556, w_eco100557, w_eco100558, w_eco100559, w_eco100560, w_eco100561, w_eco100562, w_eco100563, w_eco100564, w_eco100565, w_eco100566, w_eco100567, w_eco100568, w_eco100569, w_eco100570, w_eco100571, w_eco100572, w_eco100573, w_eco100574, w_eco100575, w_eco100576, w_eco100577, w_eco100578, w_eco100579, w_eco100580, w_eco100581, w_eco100582, w_eco100583, w_eco100584, w_eco100585, w_eco100586, w_eco100587, w_eco100588, w_eco100589, w_eco100590, w_eco100591, w_eco100592, w_eco100593, w_eco100594, w_eco100595, w_eco100596, w_eco100597, w_eco100598, w_eco100599, w_eco100600, w_eco100601, w_eco100602, w_eco100603, w_eco100604, w_eco100605, w_eco100606, w_eco100607, w_eco100608, w_eco100609, w_eco100610, w_eco100611, w_eco100612, w_eco100613, w_eco100614, w_eco100615, w_eco100616, w_eco100617, w_eco100618, w_eco100619, w_eco100620, w_eco100621, w_eco100622, w_eco100623, w_eco100624, w_eco100625, w_eco100626, w_eco100627, w_eco100628, w_eco100629, w_eco100630, w_eco100631, w_eco100632, w_eco100633, w_eco100634, w_eco100635, w_eco100636, w_eco100637, w_eco100638, w_eco100639, w_eco100640, w_eco100641, w_eco100642, w_eco100643, w_eco100644, w_eco100645, w_eco100646, w_eco100647, w_eco100648, w_eco100649, w_eco100650, w_eco100651, w_eco100652, w_eco100653, w_eco100654, w_eco100655, w_eco100656, w_eco100657, w_eco100658, w_eco100659, w_eco100660, w_eco100661, w_eco100662, w_eco100663, w_eco100664, w_eco100665, w_eco100666, w_eco100667, w_eco100668, w_eco100669, w_eco100670, w_eco100671, w_eco100672, w_eco100673, w_eco100674, w_eco100675, w_eco100676, w_eco100677, w_eco100678, w_eco100679, w_eco100680, w_eco100681, w_eco100682, w_eco100683, w_eco100684, w_eco100685, w_eco100686, w_eco100687, w_eco100688, w_eco100689, w_eco100690, w_eco100691, w_eco100692, w_eco100693, w_eco100694, w_eco100695, w_eco100696, w_eco100697, w_eco100698, w_eco100699, w_eco100700, w_eco100701, w_eco100702, w_eco100703, w_eco100704, w_eco100705, w_eco100706, w_eco100707, w_eco100708, w_eco100709, w_eco100710, w_eco100711, w_eco100712, w_eco100713, w_eco100714, w_eco100715, w_eco100716, w_eco100717, w_eco100718, w_eco100719, w_eco100720, w_eco100721, w_eco100722, w_eco100723, w_eco100724, w_eco100725, w_eco100726, w_eco100727, w_eco100728, w_eco100729, w_eco100730, w_eco100731, w_eco100732, w_eco100733, w_eco100734, w_eco100735, w_eco100736, w_eco100737, w_eco100738, w_eco100739, w_eco100740, w_eco100741, w_eco100742, w_eco100743, w_eco100744, w_eco100745, w_eco100746, w_eco100747, w_eco100748, w_eco100749, w_eco100750, w_eco100751, w_eco100752, w_eco100753, w_eco100754, w_eco100755, w_eco100756, w_eco100757, w_eco100758, w_eco100759, w_eco100760, w_eco100761, w_eco100762, w_eco100763, w_eco100764, w_eco100765, w_eco100766, w_eco100767, w_eco100768, w_eco100769, w_eco100770, w_eco100771, w_eco100772, w_eco100773, w_eco100774, w_eco100775, w_eco100776, w_eco100777, w_eco100778, w_eco100779, w_eco100780, w_eco100781, w_eco100782, w_eco100783, w_eco100784, w_eco100785, w_eco100786, w_eco100787, w_eco100788, w_eco100789, w_eco100790, w_eco100791, w_eco100792, w_eco100793, w_eco100794, w_eco100795, w_eco100796, w_eco100797, w_eco100798, w_eco100799, w_eco100800, w_eco100801, w_eco100802, w_eco100803, w_eco100804, w_eco100805, w_eco100806, w_eco100807, w_eco100808, w_eco100809, w_eco100810, w_eco100811, w_eco100812, w_eco100813, w_eco100814, w_eco100815, w_eco100816, w_eco100817, w_eco100818, w_eco100819, w_eco100820, w_eco100821, w_eco100822, w_eco100823, w_eco100824, w_eco100825, w_eco100826, w_eco100827, w_eco100828, w_eco100829, w_eco100830, w_eco100831, w_eco100832, w_eco100833, w_eco100834, w_eco100835, w_eco100836, w_eco100837, w_eco100838, w_eco100839, w_eco100840, w_eco100841, w_eco100842, w_eco100843, w_eco100844, w_eco100845, w_eco100846, w_eco100847, w_eco100848, w_eco100849, w_eco100850, w_eco100851, w_eco100852, w_eco100853, w_eco100854, w_eco100855, w_eco100856, w_eco100857, w_eco100858, w_eco100859, w_eco100860, w_eco100861, w_eco100862, w_eco100863, w_eco100864, w_eco100865, w_eco100866, w_eco100867, w_eco100868, w_eco100869, w_eco100870, w_eco100871, w_eco100872, w_eco100873, w_eco100874, w_eco100875, w_eco100876, w_eco100877, w_eco100878, w_eco100879, w_eco100880, w_eco100881, w_eco100882, w_eco100883, w_eco100884, w_eco100885, w_eco100886, w_eco100887, w_eco100888, w_eco100889, w_eco100890, w_eco100891, w_eco100892, w_eco100893, w_eco100894, w_eco100895, w_eco100896, w_eco100897, w_eco100898, w_eco100899, w_eco100900, w_eco100901, w_eco100902, w_eco100903, w_eco100904, w_eco100905, w_eco100906, w_eco100907, w_eco100908, w_eco100909, w_eco100910, w_eco100911, w_eco100912, w_eco100913, w_eco100914, w_eco100915, w_eco100916, w_eco100917, w_eco100918, w_eco100919, w_eco100920, w_eco100921, w_eco100922, w_eco100923, w_eco100924, w_eco100925, w_eco100926, w_eco100927, w_eco100928, w_eco100929, w_eco100930, w_eco100931, w_eco100932, w_eco100933, w_eco100934, w_eco100935, w_eco100936, w_eco100937, w_eco100938, w_eco100939, w_eco100940, w_eco100941, w_eco100942, w_eco100943, w_eco100944, w_eco100945, w_eco100946, w_eco100947, w_eco100948, w_eco100949, w_eco100950, w_eco100951, w_eco100952, w_eco100953, w_eco100954, w_eco100955, w_eco100956, w_eco100957, w_eco100958, w_eco100959, w_eco100960, w_eco100961, w_eco100962, w_eco100963, w_eco100964, w_eco100965, w_eco100966, w_eco100967, w_eco100968, w_eco100969, w_eco100970, w_eco100971, w_eco100972, w_eco100973, w_eco100974, w_eco100975, w_eco100976, w_eco100977, w_eco100978, w_eco100979, w_eco100980, w_eco100981, w_eco100982, w_eco100983, w_eco100984, w_eco100985, w_eco100986, w_eco100987, w_eco100988, w_eco100989, w_eco100990, w_eco100991, w_eco100992, w_eco100993, w_eco100994, w_eco100995, w_eco100996, w_eco100997, w_eco100998, w_eco100999, w_eco101000, w_eco101001, w_eco101002, w_eco101003, w_eco101004, w_eco101005, w_eco101006, w_eco101007, w_eco101008, w_eco101009, w_eco101010, w_eco101011, w_eco101012, w_eco101013, w_eco101014, w_eco101015, w_eco101016, w_eco101017, w_eco101018, w_eco101019, w_eco101020, w_eco101021, w_eco101022, w_eco101023, w_eco101024, w_eco101025, w_eco101026, w_eco101027, w_eco101028, w_eco101029, w_eco101030, w_eco101031, w_eco101032, w_eco101033, w_eco101034, w_eco101035, w_eco101036, w_eco101037, w_eco101038, w_eco101039, w_eco101040, w_eco101041, w_eco101042, w_eco101043, w_eco101044, w_eco101045, w_eco101046, w_eco101047, w_eco101048, w_eco101049, w_eco101050, w_eco101051, w_eco101052, w_eco101053, w_eco101054, w_eco101055, w_eco101056, w_eco101057, w_eco101058, w_eco101059, w_eco101060, w_eco101061, w_eco101062, w_eco101063, w_eco101064, w_eco101065, w_eco101066, w_eco101067, w_eco101068, w_eco101069, w_eco101070, w_eco101071, w_eco101072, w_eco101073, w_eco101074, w_eco101075, w_eco101076, w_eco101077, w_eco101078, w_eco101079, w_eco101080, w_eco101081, w_eco101082, w_eco101083, w_eco101084, w_eco101085, w_eco101086, w_eco101087, w_eco101088, w_eco101089, w_eco101090, w_eco101091, w_eco101092, w_eco101093, w_eco101094, w_eco101095, w_eco101096, w_eco101097, w_eco101098, w_eco101099, w_eco101100, w_eco101101, w_eco101102, w_eco101103, w_eco101104, w_eco101105, w_eco101106, w_eco101107, w_eco101108, w_eco101109, w_eco101110, w_eco101111, w_eco101112, w_eco101113, w_eco101114, w_eco101115, w_eco101116, w_eco101117, w_eco101118, w_eco101119, w_eco101120, w_eco101121, w_eco101122, w_eco101123, w_eco101124, w_eco101125, w_eco101126, w_eco101127, w_eco101128, w_eco101129, w_eco101130, w_eco101131, w_eco101132, w_eco101133, w_eco101134, w_eco101135, w_eco101136, w_eco101137, w_eco101138, w_eco101139, w_eco101140, w_eco101141, w_eco101142, w_eco101143, w_eco101144, w_eco101145, w_eco101146, w_eco101147, w_eco101148, w_eco101149, w_eco101150, w_eco101151, w_eco101152, w_eco101153, w_eco101154, w_eco101155, w_eco101156, w_eco101157, w_eco101158, w_eco101159, w_eco101160, w_eco101161, w_eco101162, w_eco101163, w_eco101164, w_eco101165, w_eco101166, w_eco101167, w_eco101168, w_eco101169, w_eco101170, w_eco101171, w_eco101172, w_eco101173, w_eco101174, w_eco101175, w_eco101176, w_eco101177, w_eco101178, w_eco101179, w_eco101180, w_eco101181, w_eco101182, w_eco101183, w_eco101184, w_eco101185, w_eco101186, w_eco101187, w_eco101188, w_eco101189, w_eco101190, w_eco101191, w_eco101192, w_eco101193, w_eco101194, w_eco101195, w_eco101196, w_eco101197, w_eco101198, w_eco101199, w_eco101200, w_eco101201, w_eco101202, w_eco101203, w_eco101204, w_eco101205, w_eco101206, w_eco101207, w_eco101208, w_eco101209, w_eco101210, w_eco101211, w_eco101212, w_eco101213, w_eco101214, w_eco101215, w_eco101216, w_eco101217, w_eco101218, w_eco101219, w_eco101220, w_eco101221, w_eco101222, w_eco101223, w_eco101224, w_eco101225, w_eco101226, w_eco101227, w_eco101228, w_eco101229, w_eco101230, w_eco101231, w_eco101232, w_eco101233, w_eco101234, w_eco101235, w_eco101236, w_eco101237, w_eco101238, w_eco101239, w_eco101240, w_eco101241, w_eco101242, w_eco101243, w_eco101244, w_eco101245, w_eco101246, w_eco101247, w_eco101248, w_eco101249, w_eco101250, w_eco101251, w_eco101252, w_eco101253, w_eco101254, w_eco101255, w_eco101256, w_eco101257, w_eco101258, w_eco101259, w_eco101260, w_eco101261, w_eco101262, w_eco101263, w_eco101264, w_eco101265, w_eco101266, w_eco101267, w_eco101268, w_eco101269, w_eco101270, w_eco101271, w_eco101272, w_eco101273, w_eco101274, w_eco101275, w_eco101276, w_eco101277, w_eco101278, w_eco101279, w_eco101280, w_eco101281, w_eco101282, w_eco101283, w_eco101284, w_eco101285, w_eco101286, w_eco101287, w_eco101288, w_eco101289, w_eco101290, w_eco101291, w_eco101292, w_eco101293, w_eco101294, w_eco101295, w_eco101296, w_eco101297, w_eco101298, w_eco101299, w_eco101300, w_eco101301, w_eco101302, w_eco101303, w_eco101304, w_eco101305, w_eco101306, w_eco101307, w_eco101308, w_eco101309, w_eco101310, w_eco101311, w_eco101312, w_eco101313, w_eco101314, w_eco101315, w_eco101316, w_eco101317, w_eco101318, w_eco101319, w_eco101320, w_eco101321, w_eco101322, w_eco101323, w_eco101324, w_eco101325, w_eco101326, w_eco101327, w_eco101328, w_eco101329, w_eco101330, w_eco101331, w_eco101332, w_eco101333, w_eco101334, w_eco101335, w_eco101336, w_eco101337, w_eco101338, w_eco101339, w_eco101340, w_eco101341, w_eco101342, w_eco101343, w_eco101344, w_eco101345, w_eco101346, w_eco101347, w_eco101348, w_eco101349, w_eco101350, w_eco101351, w_eco101352, w_eco101353, w_eco101354, w_eco101355, w_eco101356, w_eco101357, w_eco101358, w_eco101359, w_eco101360, w_eco101361, w_eco101362, w_eco101363, w_eco101364, w_eco101365, w_eco101366, w_eco101367, w_eco101368, w_eco101369, w_eco101370, w_eco101371, w_eco101372, w_eco101373, w_eco101374, w_eco101375, w_eco101376, w_eco101377, w_eco101378, w_eco101379, w_eco101380, w_eco101381, w_eco101382, w_eco101383, w_eco101384, w_eco101385, w_eco101386, w_eco101387, w_eco101388, w_eco101389, w_eco101390, w_eco101391, w_eco101392, w_eco101393, w_eco101394, w_eco101395, w_eco101396, w_eco101397, w_eco101398, w_eco101399, w_eco101400, w_eco101401, w_eco101402, w_eco101403, w_eco101404, w_eco101405, w_eco101406, w_eco101407, w_eco101408, w_eco101409, w_eco101410, w_eco101411, w_eco101412, w_eco101413, w_eco101414, w_eco101415, w_eco101416, w_eco101417, w_eco101418, w_eco101419, w_eco101420, w_eco101421, w_eco101422, w_eco101423, w_eco101424, w_eco101425, w_eco101426, w_eco101427, w_eco101428, w_eco101429, w_eco101430, w_eco101431, w_eco101432, w_eco101433, w_eco101434, w_eco101435, w_eco101436, w_eco101437, w_eco101438, w_eco101439, w_eco101440, w_eco101441, w_eco101442, w_eco101443, w_eco101444, w_eco101445, w_eco101446, w_eco101447, w_eco101448, w_eco101449, w_eco101450, w_eco101451, w_eco101452, w_eco101453, w_eco101454, w_eco101455, w_eco101456, w_eco101457, w_eco101458, w_eco101459, w_eco101460, w_eco101461, w_eco101462, w_eco101463, w_eco101464, w_eco101465, w_eco101466, w_eco101467, w_eco101468, w_eco101469, w_eco101470, w_eco101471, w_eco101472, w_eco101473, w_eco101474, w_eco101475, w_eco101476, w_eco101477, w_eco101478, w_eco101479, w_eco101480, w_eco101481, w_eco101482, w_eco101483, w_eco101484, w_eco101485, w_eco101486, w_eco101487, w_eco101488, w_eco101489, w_eco101490, w_eco101491, w_eco101492, w_eco101493, w_eco101494, w_eco101495, w_eco101496, w_eco101497, w_eco101498, w_eco101499, w_eco101500, w_eco101501, w_eco101502, w_eco101503, w_eco101504, w_eco101505, w_eco101506, w_eco101507, w_eco101508, w_eco101509, w_eco101510, w_eco101511, w_eco101512, w_eco101513, w_eco101514, w_eco101515, w_eco101516, w_eco101517, w_eco101518, w_eco101519, w_eco101520, w_eco101521, w_eco101522, w_eco101523, w_eco101524, w_eco101525, w_eco101526, w_eco101527, w_eco101528, w_eco101529, w_eco101530, w_eco101531, w_eco101532, w_eco101533, w_eco101534, w_eco101535, w_eco101536, w_eco101537, w_eco101538, w_eco101539, w_eco101540, w_eco101541, w_eco101542, w_eco101543, w_eco101544, w_eco101545, w_eco101546, w_eco101547, w_eco101548, w_eco101549, w_eco101550, w_eco101551, w_eco101552, w_eco101553, w_eco101554, w_eco101555, w_eco101556, w_eco101557, w_eco101558, w_eco101559, w_eco101560, w_eco101561, w_eco101562, w_eco101563, w_eco101564, w_eco101565, w_eco101566, w_eco101567, w_eco101568, w_eco101569, w_eco101570, w_eco101571, w_eco101572, w_eco101573, w_eco101574, w_eco101575, w_eco101576, w_eco101577, w_eco101578, w_eco101579, w_eco101580, w_eco101581, w_eco101582, w_eco101583, w_eco101584, w_eco101585, w_eco101586, w_eco101587, w_eco101588, w_eco101589, w_eco101590, w_eco101591, w_eco101592, w_eco101593, w_eco101594, w_eco101595, w_eco101596, w_eco101597, w_eco101598, w_eco101599, w_eco101600, w_eco101601, w_eco101602, w_eco101603, w_eco101604, w_eco101605, w_eco101606, w_eco101607, w_eco101608, w_eco101609, w_eco101610, w_eco101611, w_eco101612, w_eco101613, w_eco101614, w_eco101615, w_eco101616, w_eco101617, w_eco101618, w_eco101619, w_eco101620, w_eco101621, w_eco101622, w_eco101623, w_eco101624, w_eco101625, w_eco101626, w_eco101627, w_eco101628, w_eco101629, w_eco101630, w_eco101631, w_eco101632, w_eco101633, w_eco101634, w_eco101635, w_eco101636, w_eco101637, w_eco101638, w_eco101639, w_eco101640, w_eco101641, w_eco101642, w_eco101643, w_eco101644, w_eco101645, w_eco101646, w_eco101647, w_eco101648, w_eco101649, w_eco101650, w_eco101651, w_eco101652, w_eco101653, w_eco101654, w_eco101655, w_eco101656, w_eco101657, w_eco101658, w_eco101659, w_eco101660, w_eco101661, w_eco101662, w_eco101663, w_eco101664, w_eco101665, w_eco101666, w_eco101667, w_eco101668, w_eco101669, w_eco101670, w_eco101671, w_eco101672, w_eco101673, w_eco101674, w_eco101675, w_eco101676, w_eco101677, w_eco101678, w_eco101679, w_eco101680, w_eco101681, w_eco101682, w_eco101683, w_eco101684, w_eco101685, w_eco101686, w_eco101687, w_eco101688, w_eco101689, w_eco101690, w_eco101691, w_eco101692, w_eco101693, w_eco101694, w_eco101695, w_eco101696, w_eco101697, w_eco101698, w_eco101699, w_eco101700, w_eco101701, w_eco101702, w_eco101703, w_eco101704, w_eco101705, w_eco101706, w_eco101707, w_eco101708, w_eco101709, w_eco101710, w_eco101711, w_eco101712, w_eco101713, w_eco101714, w_eco101715, w_eco101716, w_eco101717, w_eco101718, w_eco101719, w_eco101720, w_eco101721, w_eco101722, w_eco101723, w_eco101724, w_eco101725, w_eco101726, w_eco101727, w_eco101728, w_eco101729, w_eco101730, w_eco101731, w_eco101732, w_eco101733, w_eco101734, w_eco101735, w_eco101736, w_eco101737, w_eco101738, w_eco101739, w_eco101740, w_eco101741, w_eco101742, w_eco101743, w_eco101744, w_eco101745, w_eco101746, w_eco101747, w_eco101748, w_eco101749, w_eco101750, w_eco101751, w_eco101752, w_eco101753, w_eco101754, w_eco101755, w_eco101756, w_eco101757, w_eco101758, w_eco101759, w_eco101760, w_eco101761, w_eco101762, w_eco101763, w_eco101764, w_eco101765, w_eco101766, w_eco101767, w_eco101768, w_eco101769, w_eco101770, w_eco101771, w_eco101772, w_eco101773, w_eco101774, w_eco101775, w_eco101776, w_eco101777, w_eco101778, w_eco101779, w_eco101780, w_eco101781, w_eco101782, w_eco101783, w_eco101784, w_eco101785, w_eco101786, w_eco101787, w_eco101788, w_eco101789, w_eco101790, w_eco101791, w_eco101792, w_eco101793, w_eco101794, w_eco101795, w_eco101796, w_eco101797, w_eco101798, w_eco101799, w_eco101800, w_eco101801, w_eco101802, w_eco101803, w_eco101804, w_eco101805, w_eco101806, w_eco101807, w_eco101808, w_eco101809, w_eco101810, w_eco101811, w_eco101812, w_eco101813, w_eco101814, w_eco101815, w_eco101816, w_eco101817, w_eco101818, w_eco101819, w_eco101820, w_eco101821, w_eco101822, w_eco101823, w_eco101824, w_eco101825, w_eco101826, w_eco101827, w_eco101828, w_eco101829, w_eco101830, w_eco101831, w_eco101832, w_eco101833, w_eco101834, w_eco101835, w_eco101836, w_eco101837, w_eco101838, w_eco101839, w_eco101840, w_eco101841, w_eco101842, w_eco101843, w_eco101844, w_eco101845, w_eco101846, w_eco101847, w_eco101848, w_eco101849, w_eco101850, w_eco101851, w_eco101852, w_eco101853, w_eco101854, w_eco101855, w_eco101856, w_eco101857, w_eco101858, w_eco101859, w_eco101860, w_eco101861, w_eco101862, w_eco101863, w_eco101864, w_eco101865, w_eco101866, w_eco101867, w_eco101868, w_eco101869, w_eco101870, w_eco101871, w_eco101872, w_eco101873, w_eco101874, w_eco101875, w_eco101876, w_eco101877, w_eco101878, w_eco101879, w_eco101880, w_eco101881, w_eco101882, w_eco101883, w_eco101884, w_eco101885, w_eco101886, w_eco101887, w_eco101888, w_eco101889, w_eco101890, w_eco101891, w_eco101892, w_eco101893, w_eco101894, w_eco101895, w_eco101896, w_eco101897, w_eco101898, w_eco101899, w_eco101900, w_eco101901, w_eco101902, w_eco101903, w_eco101904, w_eco101905, w_eco101906, w_eco101907, w_eco101908, w_eco101909, w_eco101910, w_eco101911, w_eco101912, w_eco101913, w_eco101914, w_eco101915, w_eco101916, w_eco101917, w_eco101918, w_eco101919, w_eco101920, w_eco101921, w_eco101922, w_eco101923, w_eco101924, w_eco101925, w_eco101926, w_eco101927, w_eco101928, w_eco101929, w_eco101930, w_eco101931, w_eco101932, w_eco101933, w_eco101934, w_eco101935, w_eco101936, w_eco101937, w_eco101938, w_eco101939, w_eco101940, w_eco101941, w_eco101942, w_eco101943, w_eco101944, w_eco101945, w_eco101946, w_eco101947, w_eco101948, w_eco101949, w_eco101950, w_eco101951, w_eco101952, w_eco101953, w_eco101954, w_eco101955, w_eco101956, w_eco101957, w_eco101958, w_eco101959, w_eco101960, w_eco101961, w_eco101962, w_eco101963, w_eco101964, w_eco101965, w_eco101966, w_eco101967, w_eco101968, w_eco101969, w_eco101970, w_eco101971, w_eco101972, w_eco101973, w_eco101974, w_eco101975, w_eco101976, w_eco101977, w_eco101978, w_eco101979, w_eco101980, w_eco101981, w_eco101982, w_eco101983, w_eco101984, w_eco101985, w_eco101986, w_eco101987, w_eco101988, w_eco101989, w_eco101990, w_eco101991, w_eco101992, w_eco101993, w_eco101994, w_eco101995, w_eco101996, w_eco101997, w_eco101998, w_eco101999, w_eco102000, w_eco102001, w_eco102002, w_eco102003, w_eco102004, w_eco102005, w_eco102006, w_eco102007, w_eco102008, w_eco102009, w_eco102010, w_eco102011, w_eco102012, w_eco102013, w_eco102014, w_eco102015, w_eco102016, w_eco102017, w_eco102018, w_eco102019, w_eco102020, w_eco102021, w_eco102022, w_eco102023, w_eco102024, w_eco102025, w_eco102026, w_eco102027, w_eco102028, w_eco102029, w_eco102030, w_eco102031, w_eco102032, w_eco102033, w_eco102034, w_eco102035, w_eco102036, w_eco102037, w_eco102038, w_eco102039, w_eco102040, w_eco102041, w_eco102042, w_eco102043, w_eco102044, w_eco102045, w_eco102046, w_eco102047, w_eco102048, w_eco102049, w_eco102050, w_eco102051, w_eco102052, w_eco102053, w_eco102054, w_eco102055, w_eco102056, w_eco102057, w_eco102058, w_eco102059, w_eco102060, w_eco102061, w_eco102062, w_eco102063, w_eco102064, w_eco102065, w_eco102066, w_eco102067, w_eco102068, w_eco102069, w_eco102070, w_eco102071, w_eco102072, w_eco102073, w_eco102074, w_eco102075, w_eco102076, w_eco102077, w_eco102078, w_eco102079, w_eco102080, w_eco102081, w_eco102082, w_eco102083, w_eco102084, w_eco102085, w_eco102086, w_eco102087, w_eco102088, w_eco102089, w_eco102090, w_eco102091, w_eco102092, w_eco102093, w_eco102094, w_eco102095, w_eco102096, w_eco102097, w_eco102098, w_eco102099, w_eco102100, w_eco102101, w_eco102102, w_eco102103, w_eco102104, w_eco102105, w_eco102106, w_eco102107, w_eco102108, w_eco102109, w_eco102110, w_eco102111, w_eco102112, w_eco102113, w_eco102114, w_eco102115, w_eco102116, w_eco102117, w_eco102118, w_eco102119, w_eco102120, w_eco102121, w_eco102122, w_eco102123, w_eco102124, w_eco102125, w_eco102126, w_eco102127, w_eco102128, w_eco102129, w_eco102130, w_eco102131, w_eco102132, w_eco102133, w_eco102134, w_eco102135, w_eco102136, w_eco102137, w_eco102138, w_eco102139, w_eco102140, w_eco102141, w_eco102142, w_eco102143, w_eco102144, w_eco102145, w_eco102146, w_eco102147, w_eco102148, w_eco102149, w_eco102150, w_eco102151, w_eco102152, w_eco102153, w_eco102154, w_eco102155, w_eco102156, w_eco102157, w_eco102158, w_eco102159, w_eco102160, w_eco102161, w_eco102162, w_eco102163, w_eco102164, w_eco102165, w_eco102166, w_eco102167, w_eco102168, w_eco102169, w_eco102170, w_eco102171, w_eco102172, w_eco102173, w_eco102174, w_eco102175, w_eco102176, w_eco102177, w_eco102178, w_eco102179, w_eco102180, w_eco102181, w_eco102182, w_eco102183, w_eco102184, w_eco102185, w_eco102186, w_eco102187, w_eco102188, w_eco102189, w_eco102190, w_eco102191, w_eco102192, w_eco102193, w_eco102194, w_eco102195, w_eco102196, w_eco102197, w_eco102198, w_eco102199, w_eco102200, w_eco102201, w_eco102202, w_eco102203, w_eco102204, w_eco102205, w_eco102206, w_eco102207, w_eco102208, w_eco102209, w_eco102210, w_eco102211, w_eco102212, w_eco102213, w_eco102214, w_eco102215, w_eco102216, w_eco102217, w_eco102218, w_eco102219, w_eco102220, w_eco102221, w_eco102222, w_eco102223, w_eco102224, w_eco102225, w_eco102226, w_eco102227, w_eco102228, w_eco102229, w_eco102230, w_eco102231, w_eco102232, w_eco102233, w_eco102234, w_eco102235, w_eco102236, w_eco102237, w_eco102238, w_eco102239, w_eco102240, w_eco102241, w_eco102242, w_eco102243, w_eco102244, w_eco102245, w_eco102246, w_eco102247, w_eco102248, w_eco102249, w_eco102250, w_eco102251, w_eco102252, w_eco102253, w_eco102254, w_eco102255, w_eco102256, w_eco102257, w_eco102258, w_eco102259, w_eco102260, w_eco102261, w_eco102262, w_eco102263, w_eco102264, w_eco102265, w_eco102266, w_eco102267, w_eco102268, w_eco102269, w_eco102270, w_eco102271, w_eco102272, w_eco102273, w_eco102274, w_eco102275, w_eco102276, w_eco102277, w_eco102278, w_eco102279, w_eco102280, w_eco102281, w_eco102282, w_eco102283, w_eco102284, w_eco102285, w_eco102286, w_eco102287, w_eco102288, w_eco102289, w_eco102290, w_eco102291, w_eco102292, w_eco102293, w_eco102294, w_eco102295, w_eco102296, w_eco102297, w_eco102298, w_eco102299, w_eco102300, w_eco102301, w_eco102302, w_eco102303, w_eco102304, w_eco102305, w_eco102306, w_eco102307, w_eco102308, w_eco102309, w_eco102310, w_eco102311, w_eco102312, w_eco102313, w_eco102314, w_eco102315, w_eco102316, w_eco102317, w_eco102318, w_eco102319, w_eco102320, w_eco102321, w_eco102322, w_eco102323, w_eco102324, w_eco102325, w_eco102326, w_eco102327, w_eco102328, w_eco102329, w_eco102330, w_eco102331, w_eco102332, w_eco102333, w_eco102334, w_eco102335, w_eco102336, w_eco102337, w_eco102338, w_eco102339, w_eco102340, w_eco102341, w_eco102342, w_eco102343, w_eco102344, w_eco102345, w_eco102346, w_eco102347, w_eco102348, w_eco102349, w_eco102350, w_eco102351, w_eco102352, w_eco102353, w_eco102354, w_eco102355, w_eco102356, w_eco102357, w_eco102358, w_eco102359, w_eco102360, w_eco102361, w_eco102362, w_eco102363, w_eco102364, w_eco102365, w_eco102366, w_eco102367, w_eco102368, w_eco102369, w_eco102370, w_eco102371, w_eco102372, w_eco102373, w_eco102374, w_eco102375, w_eco102376, w_eco102377, w_eco102378, w_eco102379, w_eco102380, w_eco102381, w_eco102382, w_eco102383, w_eco102384, w_eco102385, w_eco102386, w_eco102387, w_eco102388, w_eco102389, w_eco102390, w_eco102391, w_eco102392, w_eco102393, w_eco102394, w_eco102395, w_eco102396, w_eco102397, w_eco102398, w_eco102399, w_eco102400, w_eco102401, w_eco102402, w_eco102403, w_eco102404, w_eco102405, w_eco102406, w_eco102407, w_eco102408, w_eco102409, w_eco102410, w_eco102411, w_eco102412, w_eco102413, w_eco102414, w_eco102415, w_eco102416, w_eco102417, w_eco102418, w_eco102419, w_eco102420, w_eco102421, w_eco102422, w_eco102423, w_eco102424, w_eco102425, w_eco102426, w_eco102427, w_eco102428, w_eco102429, w_eco102430, w_eco102431, w_eco102432, w_eco102433, w_eco102434, w_eco102435, w_eco102436, w_eco102437, w_eco102438, w_eco102439, w_eco102440, w_eco102441, w_eco102442, w_eco102443, w_eco102444, w_eco102445, w_eco102446, w_eco102447, w_eco102448, w_eco102449, w_eco102450, w_eco102451, w_eco102452, w_eco102453, w_eco102454, w_eco102455, w_eco102456, w_eco102457, w_eco102458, w_eco102459, w_eco102460, w_eco102461, w_eco102462, w_eco102463, w_eco102464, w_eco102465, w_eco102466, w_eco102467, w_eco102468, w_eco102469, w_eco102470, w_eco102471, w_eco102472, w_eco102473, w_eco102474, w_eco102475, w_eco102476, w_eco102477, w_eco102478, w_eco102479, w_eco102480, w_eco102481, w_eco102482, w_eco102483, w_eco102484, w_eco102485, w_eco102486, w_eco102487, w_eco102488, w_eco102489, w_eco102490, w_eco102491, w_eco102492, w_eco102493, w_eco102494, w_eco102495, w_eco102496, w_eco102497, w_eco102498, w_eco102499, w_eco102500, w_eco102501, w_eco102502, w_eco102503, w_eco102504, w_eco102505, w_eco102506, w_eco102507, w_eco102508, w_eco102509, w_eco102510, w_eco102511, w_eco102512, w_eco102513, w_eco102514, w_eco102515, w_eco102516, w_eco102517, w_eco102518, w_eco102519, w_eco102520, w_eco102521, w_eco102522, w_eco102523, w_eco102524, w_eco102525, w_eco102526, w_eco102527, w_eco102528, w_eco102529, w_eco102530, w_eco102531, w_eco102532, w_eco102533, w_eco102534, w_eco102535, w_eco102536, w_eco102537, w_eco102538, w_eco102539, w_eco102540, w_eco102541, w_eco102542, w_eco102543, w_eco102544, w_eco102545, w_eco102546, w_eco102547, w_eco102548, w_eco102549, w_eco102550, w_eco102551, w_eco102552, w_eco102553, w_eco102554, w_eco102555, w_eco102556, w_eco102557, w_eco102558, w_eco102559, w_eco102560, w_eco102561, w_eco102562, w_eco102563, w_eco102564, w_eco102565, w_eco102566, w_eco102567, w_eco102568, w_eco102569, w_eco102570, w_eco102571, w_eco102572, w_eco102573, w_eco102574, w_eco102575, w_eco102576, w_eco102577, w_eco102578, w_eco102579, w_eco102580, w_eco102581, w_eco102582, w_eco102583, w_eco102584, w_eco102585, w_eco102586, w_eco102587, w_eco102588, w_eco102589, w_eco102590, w_eco102591, w_eco102592, w_eco102593, w_eco102594, w_eco102595, w_eco102596, w_eco102597, w_eco102598, w_eco102599, w_eco102600, w_eco102601, w_eco102602, w_eco102603, w_eco102604, w_eco102605, w_eco102606, w_eco102607, w_eco102608, w_eco102609, w_eco102610, w_eco102611, w_eco102612, w_eco102613, w_eco102614, w_eco102615, w_eco102616, w_eco102617, w_eco102618, w_eco102619, w_eco102620, w_eco102621, w_eco102622, w_eco102623, w_eco102624, w_eco102625, w_eco102626, w_eco102627, w_eco102628, w_eco102629, w_eco102630, w_eco102631, w_eco102632, w_eco102633, w_eco102634, w_eco102635, w_eco102636, w_eco102637, w_eco102638, w_eco102639, w_eco102640, w_eco102641, w_eco102642, w_eco102643, w_eco102644, w_eco102645, w_eco102646, w_eco102647, w_eco102648, w_eco102649, w_eco102650, w_eco102651, w_eco102652, w_eco102653, w_eco102654, w_eco102655, w_eco102656, w_eco102657, w_eco102658, w_eco102659, w_eco102660, w_eco102661, w_eco102662, w_eco102663, w_eco102664, w_eco102665, w_eco102666, w_eco102667, w_eco102668, w_eco102669, w_eco102670, w_eco102671, w_eco102672, w_eco102673, w_eco102674, w_eco102675, w_eco102676, w_eco102677, w_eco102678, w_eco102679, w_eco102680, w_eco102681, w_eco102682, w_eco102683, w_eco102684, w_eco102685, w_eco102686, w_eco102687, w_eco102688, w_eco102689, w_eco102690, w_eco102691, w_eco102692, w_eco102693, w_eco102694, w_eco102695, w_eco102696, w_eco102697, w_eco102698, w_eco102699, w_eco102700, w_eco102701, w_eco102702, w_eco102703, w_eco102704, w_eco102705, w_eco102706, w_eco102707, w_eco102708, w_eco102709, w_eco102710, w_eco102711, w_eco102712, w_eco102713, w_eco102714, w_eco102715, w_eco102716, w_eco102717, w_eco102718, w_eco102719, w_eco102720, w_eco102721, w_eco102722, w_eco102723, w_eco102724, w_eco102725, w_eco102726, w_eco102727, w_eco102728, w_eco102729, w_eco102730, w_eco102731, w_eco102732, w_eco102733, w_eco102734, w_eco102735, w_eco102736, w_eco102737, w_eco102738, w_eco102739, w_eco102740, w_eco102741, w_eco102742, w_eco102743, w_eco102744, w_eco102745, w_eco102746, w_eco102747, w_eco102748, w_eco102749, w_eco102750, w_eco102751, w_eco102752, w_eco102753, w_eco102754, w_eco102755, w_eco102756, w_eco102757, w_eco102758, w_eco102759, w_eco102760, w_eco102761, w_eco102762, w_eco102763, w_eco102764, w_eco102765, w_eco102766, w_eco102767, w_eco102768, w_eco102769, w_eco102770, w_eco102771, w_eco102772, w_eco102773, w_eco102774, w_eco102775, w_eco102776, w_eco102777, w_eco102778, w_eco102779, w_eco102780, w_eco102781, w_eco102782, w_eco102783, w_eco102784, w_eco102785, w_eco102786, w_eco102787, w_eco102788, w_eco102789, w_eco102790, w_eco102791, w_eco102792, w_eco102793, w_eco102794, w_eco102795, w_eco102796, w_eco102797, w_eco102798, w_eco102799, w_eco102800, w_eco102801, w_eco102802, w_eco102803, w_eco102804, w_eco102805, w_eco102806, w_eco102807, w_eco102808, w_eco102809, w_eco102810, w_eco102811, w_eco102812, w_eco102813, w_eco102814, w_eco102815, w_eco102816, w_eco102817, w_eco102818, w_eco102819, w_eco102820, w_eco102821, w_eco102822, w_eco102823, w_eco102824, w_eco102825, w_eco102826, w_eco102827, w_eco102828, w_eco102829, w_eco102830, w_eco102831, w_eco102832, w_eco102833, w_eco102834, w_eco102835, w_eco102836, w_eco102837, w_eco102838, w_eco102839, w_eco102840, w_eco102841, w_eco102842, w_eco102843, w_eco102844, w_eco102845, w_eco102846, w_eco102847, w_eco102848, w_eco102849, w_eco102850, w_eco102851, w_eco102852, w_eco102853, w_eco102854, w_eco102855, w_eco102856, w_eco102857, w_eco102858, w_eco102859, w_eco102860, w_eco102861, w_eco102862, w_eco102863, w_eco102864, w_eco102865, w_eco102866, w_eco102867, w_eco102868, w_eco102869, w_eco102870, w_eco102871, w_eco102872, w_eco102873, w_eco102874, w_eco102875, w_eco102876, w_eco102877, w_eco102878, w_eco102879, w_eco102880, w_eco102881, w_eco102882, w_eco102883, w_eco102884, w_eco102885, w_eco102886, w_eco102887, w_eco102888, w_eco102889, w_eco102890, w_eco102891, w_eco102892, w_eco102893, w_eco102894, w_eco102895, w_eco102896, w_eco102897, w_eco102898, w_eco102899, w_eco102900, w_eco102901, w_eco102902, w_eco102903, w_eco102904, w_eco102905, w_eco102906, w_eco102907, w_eco102908, w_eco102909, w_eco102910, w_eco102911, w_eco102912, w_eco102913, w_eco102914, w_eco102915, w_eco102916, w_eco102917, w_eco102918, w_eco102919, w_eco102920, w_eco102921, w_eco102922, w_eco102923, w_eco102924, w_eco102925, w_eco102926, w_eco102927, w_eco102928, w_eco102929, w_eco102930, w_eco102931, w_eco102932, w_eco102933, w_eco102934, w_eco102935, w_eco102936, w_eco102937, w_eco102938, w_eco102939, w_eco102940, w_eco102941, w_eco102942, w_eco102943, w_eco102944, w_eco102945, w_eco102946, w_eco102947, w_eco102948, w_eco102949, w_eco102950, w_eco102951, w_eco102952, w_eco102953, w_eco102954, w_eco102955, w_eco102956, w_eco102957, w_eco102958, w_eco102959, w_eco102960, w_eco102961, w_eco102962, w_eco102963, w_eco102964, w_eco102965, w_eco102966, w_eco102967, w_eco102968, w_eco102969, w_eco102970, w_eco102971, w_eco102972, w_eco102973, w_eco102974, w_eco102975, w_eco102976, w_eco102977, w_eco102978, w_eco102979, w_eco102980, w_eco102981, w_eco102982, w_eco102983, w_eco102984, w_eco102985, w_eco102986, w_eco102987, w_eco102988, w_eco102989, w_eco102990, w_eco102991, w_eco102992, w_eco102993, w_eco102994, w_eco102995, w_eco102996, w_eco102997, w_eco102998, w_eco102999, w_eco103000, w_eco103001, w_eco103002, w_eco103003, w_eco103004, w_eco103005, w_eco103006, w_eco103007, w_eco103008, w_eco103009, w_eco103010, w_eco103011, w_eco103012, w_eco103013, w_eco103014, w_eco103015, w_eco103016, w_eco103017, w_eco103018, w_eco103019, w_eco103020, w_eco103021, w_eco103022, w_eco103023, w_eco103024, w_eco103025, w_eco103026, w_eco103027, w_eco103028, w_eco103029, w_eco103030, w_eco103031, w_eco103032, w_eco103033, w_eco103034, w_eco103035, w_eco103036, w_eco103037, w_eco103038, w_eco103039, w_eco103040, w_eco103041, w_eco103042, w_eco103043, w_eco103044, w_eco103045, w_eco103046, w_eco103047, w_eco103048, w_eco103049, w_eco103050, w_eco103051, w_eco103052, w_eco103053, w_eco103054, w_eco103055, w_eco103056, w_eco103057, w_eco103058, w_eco103059, w_eco103060, w_eco103061, w_eco103062, w_eco103063, w_eco103064, w_eco103065, w_eco103066, w_eco103067, w_eco103068, w_eco103069, w_eco103070, w_eco103071, w_eco103072, w_eco103073, w_eco103074, w_eco103075, w_eco103076, w_eco103077, w_eco103078, w_eco103079, w_eco103080, w_eco103081, w_eco103082, w_eco103083, w_eco103084, w_eco103085, w_eco103086, w_eco103087, w_eco103088, w_eco103089, w_eco103090, w_eco103091, w_eco103092, w_eco103093, w_eco103094, w_eco103095, w_eco103096, w_eco103097, w_eco103098, w_eco103099, w_eco103100, w_eco103101, w_eco103102, w_eco103103, w_eco103104, w_eco103105, w_eco103106, w_eco103107, w_eco103108, w_eco103109, w_eco103110, w_eco103111, w_eco103112, w_eco103113, w_eco103114, w_eco103115, w_eco103116, w_eco103117, w_eco103118, w_eco103119, w_eco103120, w_eco103121, w_eco103122, w_eco103123, w_eco103124, w_eco103125, w_eco103126, w_eco103127, w_eco103128, w_eco103129, w_eco103130, w_eco103131, w_eco103132, w_eco103133, w_eco103134, w_eco103135, w_eco103136, w_eco103137, w_eco103138, w_eco103139, w_eco103140, w_eco103141, w_eco103142, w_eco103143, w_eco103144, w_eco103145, w_eco103146, w_eco103147, w_eco103148, w_eco103149, w_eco103150, w_eco103151, w_eco103152, w_eco103153, w_eco103154, w_eco103155, w_eco103156, w_eco103157, w_eco103158, w_eco103159, w_eco103160, w_eco103161, w_eco103162, w_eco103163, w_eco103164, w_eco103165, w_eco103166, w_eco103167, w_eco103168, w_eco103169, w_eco103170, w_eco103171, w_eco103172, w_eco103173, w_eco103174, w_eco103175, w_eco103176, w_eco103177, w_eco103178, w_eco103179, w_eco103180, w_eco103181, w_eco103182, w_eco103183, w_eco103184, w_eco103185, w_eco103186, w_eco103187, w_eco103188, w_eco103189, w_eco103190, w_eco103191, w_eco103192, w_eco103193, w_eco103194, w_eco103195, w_eco103196, w_eco103197, w_eco103198, w_eco103199, w_eco103200, w_eco103201, w_eco103202, w_eco103203, w_eco103204, w_eco103205, w_eco103206, w_eco103207, w_eco103208, w_eco103209, w_eco103210, w_eco103211, w_eco103212, w_eco103213, w_eco103214, w_eco103215, w_eco103216, w_eco103217, w_eco103218, w_eco103219, w_eco103220, w_eco103221, w_eco103222, w_eco103223, w_eco103224, w_eco103225, w_eco103226, w_eco103227, w_eco103228, w_eco103229, w_eco103230, w_eco103231, w_eco103232, w_eco103233, w_eco103234, w_eco103235, w_eco103236, w_eco103237, w_eco103238, w_eco103239, w_eco103240, w_eco103241, w_eco103242, w_eco103243, w_eco103244, w_eco103245, w_eco103246, w_eco103247, w_eco103248, w_eco103249, w_eco103250, w_eco103251, w_eco103252, w_eco103253, w_eco103254, w_eco103255, w_eco103256, w_eco103257, w_eco103258, w_eco103259, w_eco103260, w_eco103261, w_eco103262, w_eco103263, w_eco103264, w_eco103265, w_eco103266, w_eco103267, w_eco103268, w_eco103269, w_eco103270, w_eco103271, w_eco103272, w_eco103273, w_eco103274, w_eco103275, w_eco103276, w_eco103277, w_eco103278, w_eco103279, w_eco103280, w_eco103281, w_eco103282, w_eco103283, w_eco103284, w_eco103285, w_eco103286, w_eco103287, w_eco103288, w_eco103289, w_eco103290, w_eco103291, w_eco103292, w_eco103293, w_eco103294, w_eco103295, w_eco103296, w_eco103297, w_eco103298, w_eco103299, w_eco103300, w_eco103301, w_eco103302, w_eco103303, w_eco103304, w_eco103305, w_eco103306, w_eco103307, w_eco103308, w_eco103309, w_eco103310, w_eco103311, w_eco103312, w_eco103313, w_eco103314, w_eco103315, w_eco103316, w_eco103317, w_eco103318, w_eco103319, w_eco103320, w_eco103321, w_eco103322, w_eco103323, w_eco103324, w_eco103325, w_eco103326, w_eco103327, w_eco103328, w_eco103329, w_eco103330, w_eco103331, w_eco103332, w_eco103333, w_eco103334, w_eco103335, w_eco103336, w_eco103337, w_eco103338, w_eco103339, w_eco103340, w_eco103341, w_eco103342, w_eco103343, w_eco103344, w_eco103345, w_eco103346, w_eco103347, w_eco103348, w_eco103349, w_eco103350, w_eco103351, w_eco103352, w_eco103353, w_eco103354, w_eco103355, w_eco103356, w_eco103357, w_eco103358, w_eco103359, w_eco103360, w_eco103361, w_eco103362, w_eco103363, w_eco103364, w_eco103365, w_eco103366, w_eco103367, w_eco103368, w_eco103369, w_eco103370, w_eco103371, w_eco103372, w_eco103373, w_eco103374, w_eco103375, w_eco103376, w_eco103377, w_eco103378, w_eco103379, w_eco103380, w_eco103381, w_eco103382, w_eco103383, w_eco103384, w_eco103385, w_eco103386, w_eco103387, w_eco103388, w_eco103389, w_eco103390, w_eco103391, w_eco103392, w_eco103393, w_eco103394, w_eco103395, w_eco103396, w_eco103397, w_eco103398, w_eco103399, w_eco103400, w_eco103401, w_eco103402, w_eco103403, w_eco103404, w_eco103405, w_eco103406, w_eco103407, w_eco103408, w_eco103409, w_eco103410, w_eco103411, w_eco103412, w_eco103413, w_eco103414, w_eco103415, w_eco103416, w_eco103417, w_eco103418, w_eco103419, w_eco103420, w_eco103421, w_eco103422, w_eco103423, w_eco103424, w_eco103425, w_eco103426, w_eco103427, w_eco103428, w_eco103429, w_eco103430, w_eco103431, w_eco103432, w_eco103433, w_eco103434, w_eco103435, w_eco103436, w_eco103437, w_eco103438, w_eco103439, w_eco103440, w_eco103441, w_eco103442, w_eco103443, w_eco103444, w_eco103445, w_eco103446, w_eco103447, w_eco103448, w_eco103449, w_eco103450, w_eco103451, w_eco103452, w_eco103453, w_eco103454, w_eco103455, w_eco103456, w_eco103457, w_eco103458, w_eco103459, w_eco103460, w_eco103461, w_eco103462, w_eco103463, w_eco103464, w_eco103465, w_eco103466, w_eco103467, w_eco103468, w_eco103469, w_eco103470, w_eco103471, w_eco103472, w_eco103473, w_eco103474, w_eco103475, w_eco103476, w_eco103477, w_eco103478, w_eco103479, w_eco103480, w_eco103481, w_eco103482, w_eco103483, w_eco103484, w_eco103485, w_eco103486, w_eco103487, w_eco103488, w_eco103489, w_eco103490, w_eco103491, w_eco103492, w_eco103493, w_eco103494, w_eco103495, w_eco103496, w_eco103497, w_eco103498, w_eco103499, w_eco103500, w_eco103501, w_eco103502, w_eco103503, w_eco103504, w_eco103505, w_eco103506, w_eco103507, w_eco103508, w_eco103509, w_eco103510, w_eco103511, w_eco103512, w_eco103513, w_eco103514, w_eco103515, w_eco103516, w_eco103517, w_eco103518, w_eco103519, w_eco103520, w_eco103521, w_eco103522, w_eco103523, w_eco103524, w_eco103525, w_eco103526, w_eco103527, w_eco103528, w_eco103529, w_eco103530, w_eco103531, w_eco103532, w_eco103533, w_eco103534, w_eco103535, w_eco103536, w_eco103537, w_eco103538, w_eco103539, w_eco103540, w_eco103541, w_eco103542, w_eco103543, w_eco103544, w_eco103545, w_eco103546, w_eco103547, w_eco103548, w_eco103549, w_eco103550, w_eco103551, w_eco103552, w_eco103553, w_eco103554, w_eco103555, w_eco103556, w_eco103557, w_eco103558, w_eco103559, w_eco103560, w_eco103561, w_eco103562, w_eco103563, w_eco103564, w_eco103565, w_eco103566, w_eco103567, w_eco103568, w_eco103569, w_eco103570, w_eco103571, w_eco103572, w_eco103573, w_eco103574, w_eco103575, w_eco103576, w_eco103577, w_eco103578, w_eco103579, w_eco103580, w_eco103581, w_eco103582, w_eco103583, w_eco103584, w_eco103585, w_eco103586, w_eco103587, w_eco103588, w_eco103589, w_eco103590, w_eco103591, w_eco103592, w_eco103593, w_eco103594, w_eco103595, w_eco103596, w_eco103597, w_eco103598, w_eco103599, w_eco103600, w_eco103601, w_eco103602, w_eco103603, w_eco103604, w_eco103605, w_eco103606, w_eco103607, w_eco103608, w_eco103609, w_eco103610, w_eco103611, w_eco103612, w_eco103613, w_eco103614, w_eco103615, w_eco103616, w_eco103617, w_eco103618, w_eco103619, w_eco103620, w_eco103621, w_eco103622, w_eco103623, w_eco103624, w_eco103625, w_eco103626, w_eco103627, w_eco103628, w_eco103629, w_eco103630, w_eco103631, w_eco103632, w_eco103633, w_eco103634, w_eco103635, w_eco103636, w_eco103637, w_eco103638, w_eco103639, w_eco103640, w_eco103641, w_eco103642, w_eco103643, w_eco103644, w_eco103645, w_eco103646, w_eco103647, w_eco103648, w_eco103649, w_eco103650, w_eco103651, w_eco103652, w_eco103653, w_eco103654, w_eco103655, w_eco103656, w_eco103657, w_eco103658, w_eco103659, w_eco103660, w_eco103661, w_eco103662, w_eco103663, w_eco103664, w_eco103665, w_eco103666, w_eco103667, w_eco103668, w_eco103669, w_eco103670, w_eco103671, w_eco103672, w_eco103673, w_eco103674, w_eco103675, w_eco103676, w_eco103677, w_eco103678, w_eco103679, w_eco103680, w_eco103681, w_eco103682, w_eco103683, w_eco103684, w_eco103685, w_eco103686, w_eco103687, w_eco103688, w_eco103689, w_eco103690, w_eco103691, w_eco103692, w_eco103693, w_eco103694, w_eco103695, w_eco103696, w_eco103697, w_eco103698, w_eco103699, w_eco103700, w_eco103701, w_eco103702, w_eco103703, w_eco103704, w_eco103705, w_eco103706, w_eco103707, w_eco103708, w_eco103709, w_eco103710, w_eco103711, w_eco103712, w_eco103713, w_eco103714, w_eco103715, w_eco103716, w_eco103717, w_eco103718, w_eco103719, w_eco103720, w_eco103721, w_eco103722, w_eco103723, w_eco103724, w_eco103725, w_eco103726, w_eco103727, w_eco103728, w_eco103729, w_eco103730, w_eco103731, w_eco103732, w_eco103733, w_eco103734, w_eco103735, w_eco103736, w_eco103737, w_eco103738, w_eco103739, w_eco103740, w_eco103741, w_eco103742, w_eco103743, w_eco103744, w_eco103745, w_eco103746, w_eco103747, w_eco103748, w_eco103749, w_eco103750, w_eco103751, w_eco103752, w_eco103753, w_eco103754, w_eco103755, w_eco103756, w_eco103757, w_eco103758, w_eco103759, w_eco103760, w_eco103761, w_eco103762, w_eco103763, w_eco103764, w_eco103765, w_eco103766, w_eco103767, w_eco103768, w_eco103769, w_eco103770, w_eco103771, w_eco103772, w_eco103773, w_eco103774, w_eco103775, w_eco103776, w_eco103777, w_eco103778, w_eco103779, w_eco103780, w_eco103781, w_eco103782, w_eco103783, w_eco103784, w_eco103785, w_eco103786, w_eco103787, w_eco103788, w_eco103789, w_eco103790, w_eco103791, w_eco103792, w_eco103793, w_eco103794, w_eco103795, w_eco103796, w_eco103797, w_eco103798, w_eco103799, w_eco103800, w_eco103801, w_eco103802, w_eco103803, w_eco103804, w_eco103805, w_eco103806, w_eco103807, w_eco103808, w_eco103809, w_eco103810, w_eco103811, w_eco103812, w_eco103813, w_eco103814, w_eco103815, w_eco103816, w_eco103817, w_eco103818, w_eco103819, w_eco103820, w_eco103821, w_eco103822, w_eco103823, w_eco103824, w_eco103825, w_eco103826, w_eco103827, w_eco103828, w_eco103829, w_eco103830, w_eco103831, w_eco103832, w_eco103833, w_eco103834, w_eco103835, w_eco103836, w_eco103837, w_eco103838, w_eco103839, w_eco103840, w_eco103841, w_eco103842, w_eco103843, w_eco103844, w_eco103845, w_eco103846, w_eco103847, w_eco103848, w_eco103849, w_eco103850, w_eco103851, w_eco103852, w_eco103853, w_eco103854, w_eco103855, w_eco103856, w_eco103857, w_eco103858, w_eco103859, w_eco103860, w_eco103861, w_eco103862, w_eco103863, w_eco103864, w_eco103865, w_eco103866, w_eco103867, w_eco103868, w_eco103869, w_eco103870, w_eco103871, w_eco103872, w_eco103873, w_eco103874, w_eco103875, w_eco103876, w_eco103877, w_eco103878, w_eco103879, w_eco103880, w_eco103881, w_eco103882, w_eco103883, w_eco103884, w_eco103885, w_eco103886, w_eco103887, w_eco103888, w_eco103889, w_eco103890, w_eco103891, w_eco103892, w_eco103893, w_eco103894, w_eco103895, w_eco103896, w_eco103897, w_eco103898, w_eco103899, w_eco103900, w_eco103901, w_eco103902, w_eco103903, w_eco103904, w_eco103905, w_eco103906, w_eco103907, w_eco103908, w_eco103909, w_eco103910, w_eco103911, w_eco103912, w_eco103913, w_eco103914, w_eco103915, w_eco103916, w_eco103917, w_eco103918, w_eco103919, w_eco103920, w_eco103921, w_eco103922, w_eco103923, w_eco103924, w_eco103925, w_eco103926, w_eco103927, w_eco103928, w_eco103929, w_eco103930, w_eco103931, w_eco103932, w_eco103933, w_eco103934, w_eco103935, w_eco103936, w_eco103937, w_eco103938, w_eco103939, w_eco103940, w_eco103941, w_eco103942, w_eco103943, w_eco103944, w_eco103945, w_eco103946, w_eco103947, w_eco103948, w_eco103949, w_eco103950, w_eco103951, w_eco103952, w_eco103953, w_eco103954, w_eco103955, w_eco103956, w_eco103957, w_eco103958, w_eco103959, w_eco103960, w_eco103961, w_eco103962, w_eco103963, w_eco103964, w_eco103965, w_eco103966, w_eco103967, w_eco103968, w_eco103969, w_eco103970, w_eco103971, w_eco103972, w_eco103973, w_eco103974, w_eco103975, w_eco103976, w_eco103977, w_eco103978, w_eco103979, w_eco103980, w_eco103981, w_eco103982, w_eco103983, w_eco103984, w_eco103985, w_eco103986, w_eco103987, w_eco103988, w_eco103989, w_eco103990, w_eco103991, w_eco103992, w_eco103993, w_eco103994, w_eco103995, w_eco103996, w_eco103997, w_eco103998, w_eco103999, w_eco104000, w_eco104001, w_eco104002, w_eco104003, w_eco104004, w_eco104005, w_eco104006, w_eco104007, w_eco104008, w_eco104009, w_eco104010, w_eco104011, w_eco104012, w_eco104013, w_eco104014, w_eco104015, w_eco104016, w_eco104017, w_eco104018, w_eco104019, w_eco104020, w_eco104021, w_eco104022, w_eco104023, w_eco104024, w_eco104025, w_eco104026, w_eco104027, w_eco104028, w_eco104029, w_eco104030, w_eco104031, w_eco104032, w_eco104033, w_eco104034, w_eco104035, w_eco104036, w_eco104037, w_eco104038, w_eco104039, w_eco104040, w_eco104041, w_eco104042, w_eco104043, w_eco104044, w_eco104045, w_eco104046, w_eco104047, w_eco104048, w_eco104049, w_eco104050, w_eco104051, w_eco104052, w_eco104053, w_eco104054, w_eco104055, w_eco104056, w_eco104057, w_eco104058, w_eco104059, w_eco104060, w_eco104061, w_eco104062, w_eco104063, w_eco104064, w_eco104065, w_eco104066, w_eco104067, w_eco104068, w_eco104069, w_eco104070, w_eco104071, w_eco104072, w_eco104073, w_eco104074, w_eco104075, w_eco104076, w_eco104077, w_eco104078, w_eco104079, w_eco104080, w_eco104081, w_eco104082, w_eco104083, w_eco104084, w_eco104085, w_eco104086, w_eco104087, w_eco104088, w_eco104089, w_eco104090, w_eco104091, w_eco104092, w_eco104093, w_eco104094, w_eco104095, w_eco104096, w_eco104097, w_eco104098, w_eco104099, w_eco104100, w_eco104101, w_eco104102, w_eco104103, w_eco104104, w_eco104105, w_eco104106, w_eco104107, w_eco104108, w_eco104109, w_eco104110, w_eco104111, w_eco104112, w_eco104113, w_eco104114, w_eco104115, w_eco104116, w_eco104117, w_eco104118, w_eco104119, w_eco104120, w_eco104121, w_eco104122, w_eco104123, w_eco104124, w_eco104125, w_eco104126, w_eco104127, w_eco104128, w_eco104129, w_eco104130, w_eco104131, w_eco104132, w_eco104133, w_eco104134, w_eco104135, w_eco104136, w_eco104137, w_eco104138, w_eco104139, w_eco104140, w_eco104141, w_eco104142, w_eco104143, w_eco104144, w_eco104145, w_eco104146, w_eco104147, w_eco104148, w_eco104149, w_eco104150, w_eco104151, w_eco104152, w_eco104153, w_eco104154, w_eco104155, w_eco104156, w_eco104157, w_eco104158, w_eco104159, w_eco104160, w_eco104161, w_eco104162, w_eco104163, w_eco104164, w_eco104165, w_eco104166, w_eco104167, w_eco104168, w_eco104169, w_eco104170, w_eco104171, w_eco104172, w_eco104173, w_eco104174, w_eco104175, w_eco104176, w_eco104177, w_eco104178, w_eco104179, w_eco104180, w_eco104181, w_eco104182, w_eco104183, w_eco104184, w_eco104185, w_eco104186, w_eco104187, w_eco104188, w_eco104189, w_eco104190, w_eco104191, w_eco104192, w_eco104193, w_eco104194, w_eco104195, w_eco104196, w_eco104197, w_eco104198, w_eco104199, w_eco104200, w_eco104201, w_eco104202, w_eco104203, w_eco104204, w_eco104205, w_eco104206, w_eco104207, w_eco104208, w_eco104209, w_eco104210, w_eco104211, w_eco104212, w_eco104213, w_eco104214, w_eco104215, w_eco104216, w_eco104217, w_eco104218, w_eco104219, w_eco104220, w_eco104221, w_eco104222, w_eco104223, w_eco104224, w_eco104225, w_eco104226, w_eco104227, w_eco104228, w_eco104229, w_eco104230, w_eco104231, w_eco104232, w_eco104233, w_eco104234, w_eco104235, w_eco104236, w_eco104237, w_eco104238, w_eco104239, w_eco104240, w_eco104241, w_eco104242, w_eco104243, w_eco104244, w_eco104245, w_eco104246, w_eco104247, w_eco104248, w_eco104249, w_eco104250, w_eco104251, w_eco104252, w_eco104253, w_eco104254, w_eco104255, w_eco104256, w_eco104257, w_eco104258, w_eco104259, w_eco104260, w_eco104261, w_eco104262, w_eco104263, w_eco104264, w_eco104265, w_eco104266, w_eco104267, w_eco104268, w_eco104269, w_eco104270, w_eco104271, w_eco104272, w_eco104273, w_eco104274, w_eco104275, w_eco104276, w_eco104277, w_eco104278, w_eco104279, w_eco104280, w_eco104281, w_eco104282, w_eco104283, w_eco104284, w_eco104285, w_eco104286, w_eco104287, w_eco104288, w_eco104289, w_eco104290, w_eco104291, w_eco104292, w_eco104293, w_eco104294, w_eco104295, w_eco104296, w_eco104297, w_eco104298, w_eco104299, w_eco104300, w_eco104301, w_eco104302, w_eco104303, w_eco104304, w_eco104305, w_eco104306, w_eco104307, w_eco104308, w_eco104309, w_eco104310, w_eco104311, w_eco104312, w_eco104313, w_eco104314, w_eco104315, w_eco104316, w_eco104317, w_eco104318, w_eco104319, w_eco104320, w_eco104321, w_eco104322, w_eco104323, w_eco104324, w_eco104325, w_eco104326, w_eco104327, w_eco104328, w_eco104329, w_eco104330, w_eco104331, w_eco104332, w_eco104333, w_eco104334, w_eco104335, w_eco104336, w_eco104337, w_eco104338, w_eco104339, w_eco104340, w_eco104341, w_eco104342, w_eco104343, w_eco104344, w_eco104345, w_eco104346, w_eco104347, w_eco104348, w_eco104349, w_eco104350, w_eco104351, w_eco104352, w_eco104353, w_eco104354, w_eco104355, w_eco104356, w_eco104357, w_eco104358, w_eco104359, w_eco104360, w_eco104361, w_eco104362, w_eco104363, w_eco104364, w_eco104365, w_eco104366, w_eco104367, w_eco104368, w_eco104369, w_eco104370, w_eco104371, w_eco104372, w_eco104373, w_eco104374, w_eco104375, w_eco104376, w_eco104377, w_eco104378, w_eco104379, w_eco104380, w_eco104381, w_eco104382, w_eco104383, w_eco104384, w_eco104385, w_eco104386, w_eco104387, w_eco104388, w_eco104389, w_eco104390, w_eco104391, w_eco104392, w_eco104393, w_eco104394, w_eco104395, w_eco104396, w_eco104397, w_eco104398, w_eco104399, w_eco104400, w_eco104401, w_eco104402, w_eco104403, w_eco104404, w_eco104405, w_eco104406, w_eco104407, w_eco104408, w_eco104409, w_eco104410, w_eco104411, w_eco104412, w_eco104413, w_eco104414, w_eco104415, w_eco104416, w_eco104417, w_eco104418, w_eco104419, w_eco104420, w_eco104421, w_eco104422, w_eco104423, w_eco104424, w_eco104425, w_eco104426, w_eco104427, w_eco104428, w_eco104429, w_eco104430, w_eco104431, w_eco104432, w_eco104433, w_eco104434, w_eco104435, w_eco104436, w_eco104437, w_eco104438, w_eco104439, w_eco104440, w_eco104441, w_eco104442, w_eco104443, w_eco104444, w_eco104445, w_eco104446, w_eco104447, w_eco104448, w_eco104449, w_eco104450, w_eco104451, w_eco104452, w_eco104453, w_eco104454, w_eco104455, w_eco104456, w_eco104457, w_eco104458, w_eco104459, w_eco104460, w_eco104461, w_eco104462, w_eco104463, w_eco104464, w_eco104465, w_eco104466, w_eco104467, w_eco104468, w_eco104469, w_eco104470, w_eco104471, w_eco104472, w_eco104473, w_eco104474, w_eco104475, w_eco104476, w_eco104477, w_eco104478, w_eco104479, w_eco104480, w_eco104481, w_eco104482, w_eco104483, w_eco104484, w_eco104485, w_eco104486, w_eco104487, w_eco104488, w_eco104489, w_eco104490, w_eco104491, w_eco104492, w_eco104493, w_eco104494, w_eco104495, w_eco104496, w_eco104497, w_eco104498, w_eco104499, w_eco104500, w_eco104501, w_eco104502, w_eco104503, w_eco104504, w_eco104505, w_eco104506, w_eco104507, w_eco104508, w_eco104509, w_eco104510, w_eco104511, w_eco104512, w_eco104513, w_eco104514, w_eco104515, w_eco104516, w_eco104517, w_eco104518, w_eco104519, w_eco104520, w_eco104521, w_eco104522, w_eco104523, w_eco104524, w_eco104525, w_eco104526, w_eco104527, w_eco104528, w_eco104529, w_eco104530, w_eco104531, w_eco104532, w_eco104533, w_eco104534, w_eco104535, w_eco104536, w_eco104537, w_eco104538, w_eco104539, w_eco104540, w_eco104541, w_eco104542, w_eco104543, w_eco104544, w_eco104545, w_eco104546, w_eco104547, w_eco104548, w_eco104549, w_eco104550, w_eco104551, w_eco104552, w_eco104553, w_eco104554, w_eco104555, w_eco104556, w_eco104557, w_eco104558, w_eco104559, w_eco104560, w_eco104561, w_eco104562, w_eco104563, w_eco104564, w_eco104565, w_eco104566, w_eco104567, w_eco104568, w_eco104569, w_eco104570, w_eco104571, w_eco104572, w_eco104573, w_eco104574, w_eco104575, w_eco104576, w_eco104577, w_eco104578, w_eco104579, w_eco104580, w_eco104581, w_eco104582, w_eco104583, w_eco104584, w_eco104585, w_eco104586, w_eco104587, w_eco104588, w_eco104589, w_eco104590, w_eco104591, w_eco104592, w_eco104593, w_eco104594, w_eco104595, w_eco104596, w_eco104597, w_eco104598, w_eco104599, w_eco104600, w_eco104601, w_eco104602, w_eco104603, w_eco104604, w_eco104605, w_eco104606, w_eco104607, w_eco104608, w_eco104609, w_eco104610, w_eco104611, w_eco104612, w_eco104613, w_eco104614, w_eco104615, w_eco104616, w_eco104617, w_eco104618, w_eco104619, w_eco104620, w_eco104621, w_eco104622, w_eco104623, w_eco104624, w_eco104625, w_eco104626, w_eco104627, w_eco104628, w_eco104629, w_eco104630, w_eco104631, w_eco104632, w_eco104633, w_eco104634, w_eco104635, w_eco104636, w_eco104637, w_eco104638, w_eco104639, w_eco104640, w_eco104641, w_eco104642, w_eco104643, w_eco104644, w_eco104645, w_eco104646, w_eco104647, w_eco104648, w_eco104649, w_eco104650, w_eco104651, w_eco104652, w_eco104653, w_eco104654, w_eco104655, w_eco104656, w_eco104657, w_eco104658, w_eco104659, w_eco104660, w_eco104661, w_eco104662, w_eco104663, w_eco104664, w_eco104665, w_eco104666, w_eco104667, w_eco104668, w_eco104669, w_eco104670, w_eco104671, w_eco104672, w_eco104673, w_eco104674, w_eco104675, w_eco104676, w_eco104677, w_eco104678, w_eco104679, w_eco104680, w_eco104681, w_eco104682, w_eco104683, w_eco104684, w_eco104685, w_eco104686, w_eco104687, w_eco104688, w_eco104689, w_eco104690, w_eco104691, w_eco104692, w_eco104693, w_eco104694, w_eco104695, w_eco104696, w_eco104697, w_eco104698, w_eco104699, w_eco104700, w_eco104701, w_eco104702, w_eco104703, w_eco104704, w_eco104705, w_eco104706, w_eco104707, w_eco104708, w_eco104709, w_eco104710, w_eco104711, w_eco104712, w_eco104713, w_eco104714, w_eco104715, w_eco104716, w_eco104717, w_eco104718, w_eco104719, w_eco104720, w_eco104721, w_eco104722, w_eco104723, w_eco104724, w_eco104725, w_eco104726, w_eco104727, w_eco104728, w_eco104729, w_eco104730, w_eco104731, w_eco104732, w_eco104733, w_eco104734, w_eco104735, w_eco104736, w_eco104737, w_eco104738, w_eco104739, w_eco104740, w_eco104741, w_eco104742, w_eco104743, w_eco104744, w_eco104745, w_eco104746, w_eco104747, w_eco104748, w_eco104749, w_eco104750, w_eco104751, w_eco104752, w_eco104753, w_eco104754, w_eco104755, w_eco104756, w_eco104757, w_eco104758, w_eco104759, w_eco104760, w_eco104761, w_eco104762, w_eco104763, w_eco104764, w_eco104765, w_eco104766, w_eco104767, w_eco104768, w_eco104769, w_eco104770, w_eco104771, w_eco104772, w_eco104773, w_eco104774, w_eco104775, w_eco104776, w_eco104777, w_eco104778, w_eco104779, w_eco104780, w_eco104781, w_eco104782, w_eco104783, w_eco104784, w_eco104785, w_eco104786, w_eco104787, w_eco104788, w_eco104789, w_eco104790, w_eco104791, w_eco104792, w_eco104793, w_eco104794, w_eco104795, w_eco104796, w_eco104797, w_eco104798, w_eco104799, w_eco104800, w_eco104801, w_eco104802, w_eco104803, w_eco104804, w_eco104805, w_eco104806, w_eco104807, w_eco104808, w_eco104809, w_eco104810, w_eco104811, w_eco104812, w_eco104813, w_eco104814, w_eco104815, w_eco104816, w_eco104817, w_eco104818, w_eco104819, w_eco104820, w_eco104821, w_eco104822, w_eco104823, w_eco104824, w_eco104825, w_eco104826, w_eco104827, w_eco104828, w_eco104829, w_eco104830, w_eco104831, w_eco104832, w_eco104833, w_eco104834, w_eco104835, w_eco104836, w_eco104837, w_eco104838, w_eco104839, w_eco104840, w_eco104841, w_eco104842, w_eco104843, w_eco104844, w_eco104845, w_eco104846, w_eco104847, w_eco104848, w_eco104849, w_eco104850, w_eco104851, w_eco104852, w_eco104853, w_eco104854, w_eco104855, w_eco104856, w_eco104857, w_eco104858, w_eco104859, w_eco104860, w_eco104861, w_eco104862, w_eco104863, w_eco104864, w_eco104865, w_eco104866, w_eco104867, w_eco104868, w_eco104869, w_eco104870, w_eco104871, w_eco104872, w_eco104873, w_eco104874, w_eco104875, w_eco104876, w_eco104877, w_eco104878, w_eco104879, w_eco104880, w_eco104881, w_eco104882, w_eco104883, w_eco104884, w_eco104885, w_eco104886, w_eco104887, w_eco104888, w_eco104889, w_eco104890, w_eco104891, w_eco104892, w_eco104893, w_eco104894, w_eco104895, w_eco104896, w_eco104897, w_eco104898, w_eco104899, w_eco104900, w_eco104901, w_eco104902, w_eco104903, w_eco104904, w_eco104905, w_eco104906, w_eco104907, w_eco104908, w_eco104909, w_eco104910, w_eco104911, w_eco104912, w_eco104913, w_eco104914, w_eco104915, w_eco104916, w_eco104917, w_eco104918, w_eco104919, w_eco104920, w_eco104921, w_eco104922, w_eco104923, w_eco104924, w_eco104925, w_eco104926, w_eco104927, w_eco104928, w_eco104929, w_eco104930, w_eco104931, w_eco104932, w_eco104933, w_eco104934, w_eco104935, w_eco104936, w_eco104937, w_eco104938, w_eco104939, w_eco104940, w_eco104941, w_eco104942, w_eco104943, w_eco104944, w_eco104945, w_eco104946, w_eco104947, w_eco104948, w_eco104949, w_eco104950, w_eco104951, w_eco104952, w_eco104953, w_eco104954, w_eco104955, w_eco104956, w_eco104957, w_eco104958, w_eco104959, w_eco104960, w_eco104961, w_eco104962, w_eco104963, w_eco104964, w_eco104965, w_eco104966, w_eco104967, w_eco104968, w_eco104969, w_eco104970, w_eco104971, w_eco104972, w_eco104973, w_eco104974, w_eco104975, w_eco104976, w_eco104977, w_eco104978, w_eco104979, w_eco104980, w_eco104981, w_eco104982, w_eco104983, w_eco104984, w_eco104985, w_eco104986, w_eco104987, w_eco104988, w_eco104989, w_eco104990, w_eco104991, w_eco104992, w_eco104993, w_eco104994, w_eco104995, w_eco104996, w_eco104997, w_eco104998, w_eco104999, w_eco105000, w_eco105001, w_eco105002, w_eco105003, w_eco105004, w_eco105005, w_eco105006, w_eco105007, w_eco105008, w_eco105009, w_eco105010, w_eco105011, w_eco105012, w_eco105013, w_eco105014, w_eco105015, w_eco105016, w_eco105017, w_eco105018, w_eco105019, w_eco105020, w_eco105021, w_eco105022, w_eco105023, w_eco105024, w_eco105025, w_eco105026, w_eco105027, w_eco105028, w_eco105029, w_eco105030, w_eco105031, w_eco105032, w_eco105033, w_eco105034, w_eco105035, w_eco105036, w_eco105037, w_eco105038, w_eco105039, w_eco105040, w_eco105041, w_eco105042, w_eco105043, w_eco105044, w_eco105045, w_eco105046, w_eco105047, w_eco105048, w_eco105049, w_eco105050, w_eco105051, w_eco105052, w_eco105053, w_eco105054, w_eco105055, w_eco105056, w_eco105057, w_eco105058, w_eco105059, w_eco105060, w_eco105061, w_eco105062, w_eco105063, w_eco105064, w_eco105065, w_eco105066, w_eco105067, w_eco105068, w_eco105069, w_eco105070, w_eco105071, w_eco105072, w_eco105073, w_eco105074, w_eco105075, w_eco105076, w_eco105077, w_eco105078, w_eco105079, w_eco105080, w_eco105081, w_eco105082, w_eco105083, w_eco105084, w_eco105085, w_eco105086, w_eco105087, w_eco105088, w_eco105089, w_eco105090, w_eco105091, w_eco105092, w_eco105093, w_eco105094, w_eco105095, w_eco105096, w_eco105097, w_eco105098, w_eco105099, w_eco105100, w_eco105101, w_eco105102, w_eco105103, w_eco105104, w_eco105105, w_eco105106, w_eco105107, w_eco105108, w_eco105109, w_eco105110, w_eco105111, w_eco105112, w_eco105113, w_eco105114, w_eco105115, w_eco105116, w_eco105117, w_eco105118, w_eco105119, w_eco105120, w_eco105121, w_eco105122, w_eco105123, w_eco105124, w_eco105125, w_eco105126, w_eco105127, w_eco105128, w_eco105129, w_eco105130, w_eco105131, w_eco105132, w_eco105133, w_eco105134, w_eco105135, w_eco105136, w_eco105137, w_eco105138, w_eco105139, w_eco105140, w_eco105141, w_eco105142, w_eco105143, w_eco105144, w_eco105145, w_eco105146, w_eco105147, w_eco105148, w_eco105149, w_eco105150, w_eco105151, w_eco105152, w_eco105153, w_eco105154, w_eco105155, w_eco105156, w_eco105157, w_eco105158, w_eco105159, w_eco105160, w_eco105161, w_eco105162, w_eco105163, w_eco105164, w_eco105165, w_eco105166, w_eco105167, w_eco105168, w_eco105169, w_eco105170, w_eco105171, w_eco105172, w_eco105173, w_eco105174, w_eco105175, w_eco105176, w_eco105177, w_eco105178, w_eco105179, w_eco105180, w_eco105181, w_eco105182, w_eco105183, w_eco105184, w_eco105185, w_eco105186, w_eco105187, w_eco105188, w_eco105189, w_eco105190, w_eco105191, w_eco105192, w_eco105193, w_eco105194, w_eco105195, w_eco105196, w_eco105197, w_eco105198, w_eco105199, w_eco105200, w_eco105201, w_eco105202, w_eco105203, w_eco105204, w_eco105205, w_eco105206, w_eco105207, w_eco105208, w_eco105209, w_eco105210, w_eco105211, w_eco105212, w_eco105213, w_eco105214, w_eco105215, w_eco105216, w_eco105217, w_eco105218, w_eco105219, w_eco105220, w_eco105221, w_eco105222, w_eco105223, w_eco105224, w_eco105225, w_eco105226, w_eco105227, w_eco105228, w_eco105229, w_eco105230, w_eco105231, w_eco105232, w_eco105233, w_eco105234, w_eco105235, w_eco105236, w_eco105237, w_eco105238, w_eco105239, w_eco105240, w_eco105241, w_eco105242, w_eco105243, w_eco105244, w_eco105245, w_eco105246, w_eco105247, w_eco105248, w_eco105249, w_eco105250, w_eco105251, w_eco105252, w_eco105253, w_eco105254, w_eco105255, w_eco105256, w_eco105257, w_eco105258, w_eco105259, w_eco105260, w_eco105261, w_eco105262, w_eco105263, w_eco105264, w_eco105265, w_eco105266, w_eco105267, w_eco105268, w_eco105269, w_eco105270, w_eco105271, w_eco105272, w_eco105273, w_eco105274, w_eco105275, w_eco105276, w_eco105277, w_eco105278, w_eco105279, w_eco105280, w_eco105281, w_eco105282, w_eco105283, w_eco105284, w_eco105285, w_eco105286, w_eco105287, w_eco105288, w_eco105289, w_eco105290, w_eco105291, w_eco105292, w_eco105293, w_eco105294, w_eco105295, w_eco105296, w_eco105297, w_eco105298, w_eco105299, w_eco105300, w_eco105301, w_eco105302, w_eco105303, w_eco105304, w_eco105305, w_eco105306, w_eco105307, w_eco105308, w_eco105309, w_eco105310, w_eco105311, w_eco105312, w_eco105313, w_eco105314, w_eco105315, w_eco105316, w_eco105317, w_eco105318, w_eco105319, w_eco105320, w_eco105321, w_eco105322, w_eco105323, w_eco105324, w_eco105325, w_eco105326, w_eco105327, w_eco105328, w_eco105329, w_eco105330, w_eco105331, w_eco105332, w_eco105333, w_eco105334, w_eco105335, w_eco105336, w_eco105337, w_eco105338, w_eco105339, w_eco105340, w_eco105341, w_eco105342, w_eco105343, w_eco105344, w_eco105345, w_eco105346, w_eco105347, w_eco105348, w_eco105349, w_eco105350, w_eco105351, w_eco105352, w_eco105353, w_eco105354, w_eco105355, w_eco105356, w_eco105357, w_eco105358, w_eco105359, w_eco105360, w_eco105361, w_eco105362, w_eco105363, w_eco105364, w_eco105365, w_eco105366, w_eco105367, w_eco105368, w_eco105369, w_eco105370, w_eco105371, w_eco105372, w_eco105373, w_eco105374, w_eco105375, w_eco105376, w_eco105377, w_eco105378, w_eco105379, w_eco105380, w_eco105381, w_eco105382, w_eco105383, w_eco105384, w_eco105385, w_eco105386, w_eco105387, w_eco105388, w_eco105389, w_eco105390, w_eco105391, w_eco105392, w_eco105393, w_eco105394, w_eco105395, w_eco105396, w_eco105397, w_eco105398, w_eco105399, w_eco105400, w_eco105401, w_eco105402, w_eco105403, w_eco105404, w_eco105405, w_eco105406, w_eco105407, w_eco105408, w_eco105409, w_eco105410, w_eco105411, w_eco105412, w_eco105413, w_eco105414, w_eco105415, w_eco105416, w_eco105417, w_eco105418, w_eco105419, w_eco105420, w_eco105421, w_eco105422, w_eco105423, w_eco105424, w_eco105425, w_eco105426, w_eco105427, w_eco105428, w_eco105429, w_eco105430, w_eco105431, w_eco105432, w_eco105433, w_eco105434, w_eco105435, w_eco105436, w_eco105437, w_eco105438, w_eco105439, w_eco105440, w_eco105441, w_eco105442, w_eco105443, w_eco105444, w_eco105445, w_eco105446, w_eco105447, w_eco105448, w_eco105449, w_eco105450, w_eco105451, w_eco105452, w_eco105453, w_eco105454, w_eco105455, w_eco105456, w_eco105457, w_eco105458, w_eco105459, w_eco105460, w_eco105461, w_eco105462, w_eco105463, w_eco105464, w_eco105465, w_eco105466, w_eco105467, w_eco105468, w_eco105469, w_eco105470, w_eco105471, w_eco105472, w_eco105473, w_eco105474, w_eco105475, w_eco105476, w_eco105477, w_eco105478, w_eco105479, w_eco105480, w_eco105481, w_eco105482, w_eco105483, w_eco105484, w_eco105485, w_eco105486, w_eco105487, w_eco105488, w_eco105489, w_eco105490, w_eco105491, w_eco105492, w_eco105493, w_eco105494, w_eco105495, w_eco105496, w_eco105497, w_eco105498, w_eco105499, w_eco105500, w_eco105501, w_eco105502, w_eco105503, w_eco105504, w_eco105505, w_eco105506, w_eco105507, w_eco105508, w_eco105509, w_eco105510, w_eco105511, w_eco105512, w_eco105513, w_eco105514, w_eco105515, w_eco105516, w_eco105517, w_eco105518, w_eco105519, w_eco105520, w_eco105521, w_eco105522, w_eco105523, w_eco105524, w_eco105525, w_eco105526, w_eco105527, w_eco105528, w_eco105529, w_eco105530, w_eco105531, w_eco105532, w_eco105533, w_eco105534, w_eco105535, w_eco105536, w_eco105537, w_eco105538, w_eco105539, w_eco105540, w_eco105541, w_eco105542, w_eco105543, w_eco105544, w_eco105545, w_eco105546, w_eco105547, w_eco105548, w_eco105549, w_eco105550, w_eco105551, w_eco105552, w_eco105553, w_eco105554, w_eco105555, w_eco105556, w_eco105557, w_eco105558, w_eco105559, w_eco105560, w_eco105561, w_eco105562, w_eco105563, w_eco105564, w_eco105565, w_eco105566, w_eco105567, w_eco105568, w_eco105569, w_eco105570, w_eco105571, w_eco105572, w_eco105573, w_eco105574, w_eco105575, w_eco105576, w_eco105577, w_eco105578, w_eco105579, w_eco105580, w_eco105581, w_eco105582, w_eco105583, w_eco105584, w_eco105585, w_eco105586, w_eco105587, w_eco105588, w_eco105589, w_eco105590, w_eco105591, w_eco105592, w_eco105593, w_eco105594, w_eco105595, w_eco105596, w_eco105597, w_eco105598, w_eco105599, w_eco105600, w_eco105601, w_eco105602, w_eco105603, w_eco105604, w_eco105605, w_eco105606, w_eco105607, w_eco105608, w_eco105609, w_eco105610, w_eco105611, w_eco105612, w_eco105613, w_eco105614, w_eco105615, w_eco105616, w_eco105617, w_eco105618, w_eco105619, w_eco105620, w_eco105621, w_eco105622, w_eco105623, w_eco105624, w_eco105625, w_eco105626, w_eco105627, w_eco105628, w_eco105629, w_eco105630, w_eco105631, w_eco105632, w_eco105633, w_eco105634, w_eco105635, w_eco105636, w_eco105637, w_eco105638, w_eco105639, w_eco105640, w_eco105641, w_eco105642, w_eco105643, w_eco105644, w_eco105645, w_eco105646, w_eco105647, w_eco105648, w_eco105649, w_eco105650, w_eco105651, w_eco105652, w_eco105653, w_eco105654, w_eco105655, w_eco105656, w_eco105657, w_eco105658, w_eco105659, w_eco105660, w_eco105661, w_eco105662, w_eco105663, w_eco105664, w_eco105665, w_eco105666, w_eco105667, w_eco105668, w_eco105669, w_eco105670, w_eco105671, w_eco105672, w_eco105673, w_eco105674, w_eco105675, w_eco105676, w_eco105677, w_eco105678, w_eco105679, w_eco105680, w_eco105681, w_eco105682, w_eco105683, w_eco105684, w_eco105685, w_eco105686, w_eco105687, w_eco105688, w_eco105689, w_eco105690, w_eco105691, w_eco105692, w_eco105693, w_eco105694, w_eco105695, w_eco105696, w_eco105697, w_eco105698, w_eco105699, w_eco105700, w_eco105701, w_eco105702, w_eco105703, w_eco105704, w_eco105705, w_eco105706, w_eco105707, w_eco105708, w_eco105709, w_eco105710, w_eco105711, w_eco105712, w_eco105713, w_eco105714, w_eco105715, w_eco105716, w_eco105717, w_eco105718, w_eco105719, w_eco105720, w_eco105721, w_eco105722, w_eco105723, w_eco105724, w_eco105725, w_eco105726, w_eco105727, w_eco105728, w_eco105729, w_eco105730, w_eco105731, w_eco105732, w_eco105733, w_eco105734, w_eco105735, w_eco105736, w_eco105737, w_eco105738, w_eco105739, w_eco105740, w_eco105741, w_eco105742, w_eco105743, w_eco105744, w_eco105745, w_eco105746, w_eco105747, w_eco105748, w_eco105749, w_eco105750, w_eco105751, w_eco105752, w_eco105753, w_eco105754, w_eco105755, w_eco105756, w_eco105757, w_eco105758, w_eco105759, w_eco105760, w_eco105761, w_eco105762, w_eco105763, w_eco105764, w_eco105765, w_eco105766, w_eco105767, w_eco105768, w_eco105769, w_eco105770, w_eco105771, w_eco105772, w_eco105773, w_eco105774, w_eco105775, w_eco105776, w_eco105777, w_eco105778, w_eco105779, w_eco105780, w_eco105781, w_eco105782, w_eco105783, w_eco105784, w_eco105785, w_eco105786, w_eco105787, w_eco105788, w_eco105789, w_eco105790, w_eco105791, w_eco105792, w_eco105793, w_eco105794, w_eco105795, w_eco105796, w_eco105797, w_eco105798, w_eco105799, w_eco105800, w_eco105801, w_eco105802, w_eco105803, w_eco105804, w_eco105805, w_eco105806, w_eco105807, w_eco105808, w_eco105809, w_eco105810, w_eco105811, w_eco105812, w_eco105813, w_eco105814, w_eco105815, w_eco105816, w_eco105817, w_eco105818, w_eco105819, w_eco105820, w_eco105821, w_eco105822, w_eco105823, w_eco105824, w_eco105825, w_eco105826, w_eco105827, w_eco105828, w_eco105829, w_eco105830, w_eco105831, w_eco105832, w_eco105833, w_eco105834, w_eco105835, w_eco105836, w_eco105837, w_eco105838, w_eco105839, w_eco105840, w_eco105841, w_eco105842, w_eco105843, w_eco105844, w_eco105845, w_eco105846, w_eco105847, w_eco105848, w_eco105849, w_eco105850, w_eco105851, w_eco105852, w_eco105853, w_eco105854, w_eco105855, w_eco105856, w_eco105857, w_eco105858, w_eco105859, w_eco105860, w_eco105861, w_eco105862, w_eco105863, w_eco105864, w_eco105865, w_eco105866, w_eco105867, w_eco105868, w_eco105869, w_eco105870, w_eco105871, w_eco105872, w_eco105873, w_eco105874, w_eco105875, w_eco105876, w_eco105877, w_eco105878, w_eco105879, w_eco105880, w_eco105881, w_eco105882, w_eco105883, w_eco105884, w_eco105885, w_eco105886, w_eco105887, w_eco105888, w_eco105889, w_eco105890, w_eco105891, w_eco105892, w_eco105893, w_eco105894, w_eco105895, w_eco105896, w_eco105897, w_eco105898, w_eco105899, w_eco105900, w_eco105901, w_eco105902, w_eco105903, w_eco105904, w_eco105905, w_eco105906, w_eco105907, w_eco105908, w_eco105909, w_eco105910, w_eco105911, w_eco105912, w_eco105913, w_eco105914, w_eco105915, w_eco105916, w_eco105917, w_eco105918, w_eco105919, w_eco105920, w_eco105921, w_eco105922, w_eco105923, w_eco105924, w_eco105925, w_eco105926, w_eco105927, w_eco105928, w_eco105929, w_eco105930, w_eco105931, w_eco105932, w_eco105933, w_eco105934, w_eco105935, w_eco105936, w_eco105937, w_eco105938, w_eco105939, w_eco105940, w_eco105941, w_eco105942, w_eco105943, w_eco105944, w_eco105945, w_eco105946, w_eco105947, w_eco105948, w_eco105949, w_eco105950, w_eco105951, w_eco105952, w_eco105953, w_eco105954, w_eco105955, w_eco105956, w_eco105957, w_eco105958, w_eco105959, w_eco105960, w_eco105961, w_eco105962, w_eco105963, w_eco105964, w_eco105965, w_eco105966, w_eco105967, w_eco105968, w_eco105969, w_eco105970, w_eco105971, w_eco105972, w_eco105973, w_eco105974, w_eco105975, w_eco105976, w_eco105977, w_eco105978, w_eco105979, w_eco105980, w_eco105981, w_eco105982, w_eco105983, w_eco105984, w_eco105985, w_eco105986, w_eco105987, w_eco105988, w_eco105989, w_eco105990, w_eco105991, w_eco105992, w_eco105993, w_eco105994, w_eco105995, w_eco105996, w_eco105997, w_eco105998, w_eco105999, w_eco106000, w_eco106001, w_eco106002, w_eco106003, w_eco106004, w_eco106005, w_eco106006, w_eco106007, w_eco106008, w_eco106009, w_eco106010, w_eco106011, w_eco106012, w_eco106013, w_eco106014, w_eco106015, w_eco106016, w_eco106017, w_eco106018, w_eco106019, w_eco106020, w_eco106021, w_eco106022, w_eco106023, w_eco106024, w_eco106025, w_eco106026, w_eco106027, w_eco106028, w_eco106029, w_eco106030, w_eco106031, w_eco106032, w_eco106033, w_eco106034, w_eco106035, w_eco106036, w_eco106037, w_eco106038, w_eco106039, w_eco106040, w_eco106041, w_eco106042, w_eco106043, w_eco106044, w_eco106045, w_eco106046, w_eco106047, w_eco106048, w_eco106049, w_eco106050, w_eco106051, w_eco106052, w_eco106053, w_eco106054, w_eco106055, w_eco106056, w_eco106057, w_eco106058, w_eco106059, w_eco106060, w_eco106061, w_eco106062, w_eco106063, w_eco106064, w_eco106065, w_eco106066, w_eco106067, w_eco106068, w_eco106069, w_eco106070, w_eco106071, w_eco106072, w_eco106073, w_eco106074, w_eco106075, w_eco106076, w_eco106077, w_eco106078, w_eco106079, w_eco106080, w_eco106081, w_eco106082, w_eco106083, w_eco106084, w_eco106085, w_eco106086, w_eco106087, w_eco106088, w_eco106089, w_eco106090, w_eco106091, w_eco106092, w_eco106093, w_eco106094, w_eco106095, w_eco106096, w_eco106097, w_eco106098, w_eco106099, w_eco106100, w_eco106101, w_eco106102, w_eco106103, w_eco106104, w_eco106105, w_eco106106, w_eco106107, w_eco106108, w_eco106109, w_eco106110, w_eco106111, w_eco106112, w_eco106113, w_eco106114, w_eco106115, w_eco106116, w_eco106117, w_eco106118, w_eco106119, w_eco106120, w_eco106121, w_eco106122, w_eco106123, w_eco106124, w_eco106125, w_eco106126, w_eco106127, w_eco106128, w_eco106129, w_eco106130, w_eco106131, w_eco106132, w_eco106133, w_eco106134, w_eco106135, w_eco106136, w_eco106137, w_eco106138, w_eco106139, w_eco106140, w_eco106141, w_eco106142, w_eco106143, w_eco106144, w_eco106145, w_eco106146, w_eco106147, w_eco106148, w_eco106149, w_eco106150, w_eco106151, w_eco106152, w_eco106153, w_eco106154, w_eco106155, w_eco106156, w_eco106157, w_eco106158, w_eco106159, w_eco106160, w_eco106161, w_eco106162, w_eco106163, w_eco106164, w_eco106165, w_eco106166, w_eco106167, w_eco106168, w_eco106169, w_eco106170, w_eco106171, w_eco106172, w_eco106173, w_eco106174, w_eco106175, w_eco106176, w_eco106177, w_eco106178, w_eco106179, w_eco106180, w_eco106181, w_eco106182, w_eco106183, w_eco106184, w_eco106185, w_eco106186, w_eco106187, w_eco106188, w_eco106189, w_eco106190, w_eco106191, w_eco106192, w_eco106193, w_eco106194, w_eco106195, w_eco106196, w_eco106197, w_eco106198, w_eco106199, w_eco106200, w_eco106201, w_eco106202, w_eco106203, w_eco106204, w_eco106205, w_eco106206, w_eco106207, w_eco106208, w_eco106209, w_eco106210, w_eco106211, w_eco106212, w_eco106213, w_eco106214, w_eco106215, w_eco106216, w_eco106217, w_eco106218, w_eco106219, w_eco106220, w_eco106221, w_eco106222, w_eco106223, w_eco106224, w_eco106225, w_eco106226, w_eco106227, w_eco106228, w_eco106229, w_eco106230, w_eco106231, w_eco106232, w_eco106233, w_eco106234, w_eco106235, w_eco106236, w_eco106237, w_eco106238, w_eco106239, w_eco106240, w_eco106241, w_eco106242, w_eco106243, w_eco106244, w_eco106245, w_eco106246, w_eco106247, w_eco106248, w_eco106249, w_eco106250, w_eco106251, w_eco106252, w_eco106253, w_eco106254, w_eco106255, w_eco106256, w_eco106257, w_eco106258, w_eco106259, w_eco106260, w_eco106261, w_eco106262, w_eco106263, w_eco106264, w_eco106265, w_eco106266, w_eco106267, w_eco106268, w_eco106269, w_eco106270, w_eco106271, w_eco106272, w_eco106273, w_eco106274, w_eco106275, w_eco106276, w_eco106277, w_eco106278, w_eco106279, w_eco106280, w_eco106281, w_eco106282, w_eco106283, w_eco106284, w_eco106285, w_eco106286, w_eco106287, w_eco106288, w_eco106289, w_eco106290, w_eco106291, w_eco106292, w_eco106293, w_eco106294, w_eco106295, w_eco106296, w_eco106297, w_eco106298, w_eco106299, w_eco106300, w_eco106301, w_eco106302, w_eco106303, w_eco106304, w_eco106305, w_eco106306, w_eco106307, w_eco106308, w_eco106309, w_eco106310, w_eco106311, w_eco106312, w_eco106313, w_eco106314, w_eco106315, w_eco106316, w_eco106317, w_eco106318, w_eco106319, w_eco106320, w_eco106321, w_eco106322, w_eco106323, w_eco106324, w_eco106325, w_eco106326, w_eco106327, w_eco106328, w_eco106329, w_eco106330, w_eco106331, w_eco106332, w_eco106333, w_eco106334, w_eco106335, w_eco106336, w_eco106337, w_eco106338, w_eco106339, w_eco106340, w_eco106341, w_eco106342, w_eco106343, w_eco106344, w_eco106345, w_eco106346, w_eco106347, w_eco106348, w_eco106349, w_eco106350, w_eco106351, w_eco106352, w_eco106353, w_eco106354, w_eco106355, w_eco106356, w_eco106357, w_eco106358, w_eco106359, w_eco106360, w_eco106361, w_eco106362, w_eco106363, w_eco106364, w_eco106365, w_eco106366, w_eco106367, w_eco106368, w_eco106369, w_eco106370, w_eco106371, w_eco106372, w_eco106373, w_eco106374, w_eco106375, w_eco106376, w_eco106377, w_eco106378, w_eco106379, w_eco106380, w_eco106381, w_eco106382, w_eco106383, w_eco106384, w_eco106385, w_eco106386, w_eco106387, w_eco106388, w_eco106389, w_eco106390, w_eco106391, w_eco106392, w_eco106393, w_eco106394, w_eco106395, w_eco106396, w_eco106397, w_eco106398, w_eco106399, w_eco106400, w_eco106401, w_eco106402, w_eco106403, w_eco106404, w_eco106405, w_eco106406, w_eco106407, w_eco106408, w_eco106409, w_eco106410, w_eco106411, w_eco106412, w_eco106413, w_eco106414, w_eco106415, w_eco106416, w_eco106417, w_eco106418, w_eco106419, w_eco106420, w_eco106421, w_eco106422, w_eco106423, w_eco106424, w_eco106425, w_eco106426, w_eco106427, w_eco106428, w_eco106429, w_eco106430, w_eco106431, w_eco106432, w_eco106433, w_eco106434, w_eco106435, w_eco106436, w_eco106437, w_eco106438, w_eco106439, w_eco106440, w_eco106441, w_eco106442, w_eco106443, w_eco106444, w_eco106445, w_eco106446, w_eco106447, w_eco106448, w_eco106449, w_eco106450, w_eco106451, w_eco106452, w_eco106453, w_eco106454, w_eco106455, w_eco106456, w_eco106457, w_eco106458, w_eco106459, w_eco106460, w_eco106461, w_eco106462, w_eco106463, w_eco106464, w_eco106465, w_eco106466, w_eco106467, w_eco106468, w_eco106469, w_eco106470, w_eco106471, w_eco106472, w_eco106473, w_eco106474, w_eco106475, w_eco106476, w_eco106477, w_eco106478, w_eco106479, w_eco106480, w_eco106481, w_eco106482, w_eco106483, w_eco106484, w_eco106485, w_eco106486, w_eco106487, w_eco106488, w_eco106489, w_eco106490, w_eco106491, w_eco106492, w_eco106493, w_eco106494, w_eco106495, w_eco106496, w_eco106497, w_eco106498, w_eco106499, w_eco106500, w_eco106501, w_eco106502, w_eco106503, w_eco106504, w_eco106505, w_eco106506, w_eco106507, w_eco106508, w_eco106509, w_eco106510, w_eco106511, w_eco106512, w_eco106513, w_eco106514, w_eco106515, w_eco106516, w_eco106517, w_eco106518, w_eco106519, w_eco106520, w_eco106521, w_eco106522, w_eco106523, w_eco106524, w_eco106525, w_eco106526, w_eco106527, w_eco106528, w_eco106529, w_eco106530, w_eco106531, w_eco106532, w_eco106533, w_eco106534, w_eco106535, w_eco106536, w_eco106537, w_eco106538, w_eco106539, w_eco106540, w_eco106541, w_eco106542, w_eco106543, w_eco106544, w_eco106545, w_eco106546, w_eco106547, w_eco106548, w_eco106549, w_eco106550, w_eco106551, w_eco106552, w_eco106553, w_eco106554, w_eco106555, w_eco106556, w_eco106557, w_eco106558, w_eco106559, w_eco106560, w_eco106561, w_eco106562, w_eco106563, w_eco106564, w_eco106565, w_eco106566, w_eco106567, w_eco106568, w_eco106569, w_eco106570, w_eco106571, w_eco106572, w_eco106573, w_eco106574, w_eco106575, w_eco106576, w_eco106577, w_eco106578, w_eco106579, w_eco106580, w_eco106581, w_eco106582, w_eco106583, w_eco106584, w_eco106585, w_eco106586, w_eco106587, w_eco106588, w_eco106589, w_eco106590, w_eco106591, w_eco106592, w_eco106593, w_eco106594, w_eco106595, w_eco106596, w_eco106597, w_eco106598, w_eco106599, w_eco106600, w_eco106601, w_eco106602, w_eco106603, w_eco106604, w_eco106605, w_eco106606, w_eco106607, w_eco106608, w_eco106609, w_eco106610, w_eco106611, w_eco106612, w_eco106613, w_eco106614, w_eco106615, w_eco106616, w_eco106617, w_eco106618, w_eco106619, w_eco106620, w_eco106621, w_eco106622, w_eco106623, w_eco106624, w_eco106625, w_eco106626, w_eco106627, w_eco106628, w_eco106629, w_eco106630, w_eco106631, w_eco106632, w_eco106633, w_eco106634, w_eco106635, w_eco106636, w_eco106637, w_eco106638, w_eco106639, w_eco106640, w_eco106641, w_eco106642, w_eco106643, w_eco106644, w_eco106645, w_eco106646, w_eco106647, w_eco106648, w_eco106649, w_eco106650, w_eco106651, w_eco106652, w_eco106653, w_eco106654, w_eco106655, w_eco106656, w_eco106657, w_eco106658, w_eco106659, w_eco106660, w_eco106661, w_eco106662, w_eco106663, w_eco106664, w_eco106665, w_eco106666, w_eco106667, w_eco106668, w_eco106669, w_eco106670, w_eco106671, w_eco106672, w_eco106673, w_eco106674, w_eco106675, w_eco106676, w_eco106677, w_eco106678, w_eco106679, w_eco106680, w_eco106681, w_eco106682, w_eco106683, w_eco106684, w_eco106685, w_eco106686, w_eco106687, w_eco106688, w_eco106689, w_eco106690, w_eco106691, w_eco106692, w_eco106693, w_eco106694, w_eco106695, w_eco106696, w_eco106697, w_eco106698, w_eco106699, w_eco106700, w_eco106701, w_eco106702, w_eco106703, w_eco106704, w_eco106705, w_eco106706, w_eco106707, w_eco106708, w_eco106709, w_eco106710, w_eco106711, w_eco106712, w_eco106713, w_eco106714, w_eco106715, w_eco106716, w_eco106717, w_eco106718, w_eco106719, w_eco106720, w_eco106721, w_eco106722, w_eco106723, w_eco106724, w_eco106725, w_eco106726, w_eco106727, w_eco106728, w_eco106729, w_eco106730, w_eco106731, w_eco106732, w_eco106733, w_eco106734, w_eco106735, w_eco106736, w_eco106737, w_eco106738, w_eco106739, w_eco106740, w_eco106741, w_eco106742, w_eco106743, w_eco106744, w_eco106745, w_eco106746, w_eco106747, w_eco106748, w_eco106749, w_eco106750, w_eco106751, w_eco106752, w_eco106753, w_eco106754, w_eco106755, w_eco106756, w_eco106757, w_eco106758, w_eco106759, w_eco106760, w_eco106761, w_eco106762, w_eco106763, w_eco106764, w_eco106765, w_eco106766, w_eco106767, w_eco106768, w_eco106769, w_eco106770, w_eco106771, w_eco106772, w_eco106773, w_eco106774, w_eco106775, w_eco106776, w_eco106777, w_eco106778, w_eco106779, w_eco106780, w_eco106781, w_eco106782, w_eco106783, w_eco106784, w_eco106785, w_eco106786, w_eco106787, w_eco106788, w_eco106789, w_eco106790, w_eco106791, w_eco106792, w_eco106793, w_eco106794, w_eco106795, w_eco106796, w_eco106797, w_eco106798, w_eco106799, w_eco106800, w_eco106801, w_eco106802, w_eco106803, w_eco106804, w_eco106805, w_eco106806, w_eco106807, w_eco106808, w_eco106809, w_eco106810, w_eco106811, w_eco106812, w_eco106813, w_eco106814, w_eco106815, w_eco106816, w_eco106817, w_eco106818, w_eco106819, w_eco106820, w_eco106821, w_eco106822, w_eco106823, w_eco106824, w_eco106825, w_eco106826, w_eco106827, w_eco106828, w_eco106829, w_eco106830, w_eco106831, w_eco106832, w_eco106833, w_eco106834, w_eco106835, w_eco106836, w_eco106837, w_eco106838, w_eco106839, w_eco106840, w_eco106841, w_eco106842, w_eco106843, w_eco106844, w_eco106845, w_eco106846, w_eco106847, w_eco106848, w_eco106849, w_eco106850, w_eco106851, w_eco106852, w_eco106853, w_eco106854, w_eco106855, w_eco106856, w_eco106857, w_eco106858, w_eco106859, w_eco106860, w_eco106861, w_eco106862, w_eco106863, w_eco106864, w_eco106865, w_eco106866, w_eco106867, w_eco106868, w_eco106869, w_eco106870, w_eco106871, w_eco106872, w_eco106873, w_eco106874, w_eco106875, w_eco106876, w_eco106877, w_eco106878, w_eco106879, w_eco106880, w_eco106881, w_eco106882, w_eco106883, w_eco106884, w_eco106885, w_eco106886, w_eco106887, w_eco106888, w_eco106889, w_eco106890, w_eco106891, w_eco106892, w_eco106893, w_eco106894, w_eco106895, w_eco106896, w_eco106897, w_eco106898, w_eco106899, w_eco106900, w_eco106901, w_eco106902, w_eco106903, w_eco106904, w_eco106905, w_eco106906, w_eco106907, w_eco106908, w_eco106909, w_eco106910, w_eco106911, w_eco106912, w_eco106913, w_eco106914, w_eco106915, w_eco106916, w_eco106917, w_eco106918, w_eco106919, w_eco106920, w_eco106921, w_eco106922, w_eco106923, w_eco106924, w_eco106925, w_eco106926, w_eco106927, w_eco106928, w_eco106929, w_eco106930, w_eco106931, w_eco106932, w_eco106933, w_eco106934, w_eco106935, w_eco106936, w_eco106937, w_eco106938, w_eco106939, w_eco106940, w_eco106941, w_eco106942, w_eco106943, w_eco106944, w_eco106945, w_eco106946, w_eco106947, w_eco106948, w_eco106949, w_eco106950, w_eco106951, w_eco106952, w_eco106953, w_eco106954, w_eco106955, w_eco106956, w_eco106957, w_eco106958, w_eco106959, w_eco106960, w_eco106961, w_eco106962, w_eco106963, w_eco106964, w_eco106965, w_eco106966, w_eco106967, w_eco106968, w_eco106969, w_eco106970, w_eco106971, w_eco106972, w_eco106973, w_eco106974, w_eco106975, w_eco106976, w_eco106977, w_eco106978, w_eco106979, w_eco106980, w_eco106981, w_eco106982, w_eco106983, w_eco106984, w_eco106985, w_eco106986, w_eco106987, w_eco106988, w_eco106989, w_eco106990, w_eco106991, w_eco106992, w_eco106993, w_eco106994, w_eco106995, w_eco106996, w_eco106997, w_eco106998, w_eco106999, w_eco107000, w_eco107001, w_eco107002, w_eco107003, w_eco107004, w_eco107005, w_eco107006, w_eco107007, w_eco107008, w_eco107009, w_eco107010, w_eco107011, w_eco107012, w_eco107013, w_eco107014, w_eco107015, w_eco107016, w_eco107017, w_eco107018, w_eco107019, w_eco107020, w_eco107021, w_eco107022, w_eco107023, w_eco107024, w_eco107025, w_eco107026, w_eco107027, w_eco107028, w_eco107029, w_eco107030, w_eco107031, w_eco107032, w_eco107033, w_eco107034, w_eco107035, w_eco107036, w_eco107037, w_eco107038, w_eco107039, w_eco107040, w_eco107041, w_eco107042, w_eco107043, w_eco107044, w_eco107045, w_eco107046, w_eco107047, w_eco107048, w_eco107049, w_eco107050, w_eco107051, w_eco107052, w_eco107053, w_eco107054, w_eco107055, w_eco107056, w_eco107057, w_eco107058, w_eco107059, w_eco107060, w_eco107061, w_eco107062, w_eco107063, w_eco107064, w_eco107065, w_eco107066, w_eco107067, w_eco107068, w_eco107069, w_eco107070, w_eco107071, w_eco107072, w_eco107073, w_eco107074, w_eco107075, w_eco107076, w_eco107077, w_eco107078, w_eco107079, w_eco107080, w_eco107081, w_eco107082, w_eco107083, w_eco107084, w_eco107085, w_eco107086, w_eco107087, w_eco107088, w_eco107089, w_eco107090, w_eco107091, w_eco107092, w_eco107093, w_eco107094, w_eco107095, w_eco107096, w_eco107097, w_eco107098, w_eco107099, w_eco107100, w_eco107101, w_eco107102, w_eco107103, w_eco107104, w_eco107105, w_eco107106, w_eco107107, w_eco107108, w_eco107109, w_eco107110, w_eco107111, w_eco107112, w_eco107113, w_eco107114, w_eco107115, w_eco107116, w_eco107117, w_eco107118, w_eco107119, w_eco107120, w_eco107121, w_eco107122, w_eco107123, w_eco107124, w_eco107125, w_eco107126, w_eco107127, w_eco107128, w_eco107129, w_eco107130, w_eco107131, w_eco107132, w_eco107133, w_eco107134, w_eco107135, w_eco107136, w_eco107137, w_eco107138, w_eco107139, w_eco107140, w_eco107141, w_eco107142, w_eco107143, w_eco107144, w_eco107145, w_eco107146, w_eco107147, w_eco107148, w_eco107149, w_eco107150, w_eco107151, w_eco107152, w_eco107153, w_eco107154, w_eco107155, w_eco107156, w_eco107157, w_eco107158, w_eco107159, w_eco107160, w_eco107161, w_eco107162, w_eco107163, w_eco107164, w_eco107165, w_eco107166, w_eco107167, w_eco107168, w_eco107169, w_eco107170, w_eco107171, w_eco107172, w_eco107173, w_eco107174, w_eco107175, w_eco107176, w_eco107177, w_eco107178, w_eco107179, w_eco107180, w_eco107181, w_eco107182, w_eco107183, w_eco107184, w_eco107185, w_eco107186, w_eco107187, w_eco107188, w_eco107189, w_eco107190, w_eco107191, w_eco107192, w_eco107193, w_eco107194, w_eco107195, w_eco107196, w_eco107197, w_eco107198, w_eco107199, w_eco107200, w_eco107201, w_eco107202, w_eco107203, w_eco107204, w_eco107205, w_eco107206, w_eco107207, w_eco107208, w_eco107209, w_eco107210, w_eco107211, w_eco107212, w_eco107213, w_eco107214, w_eco107215, w_eco107216, w_eco107217, w_eco107218, w_eco107219, w_eco107220, w_eco107221, w_eco107222, w_eco107223, w_eco107224, w_eco107225, w_eco107226, w_eco107227, w_eco107228, w_eco107229, w_eco107230, w_eco107231, w_eco107232, w_eco107233, w_eco107234, w_eco107235, w_eco107236, w_eco107237, w_eco107238, w_eco107239, w_eco107240, w_eco107241, w_eco107242, w_eco107243, w_eco107244, w_eco107245, w_eco107246, w_eco107247, w_eco107248, w_eco107249, w_eco107250, w_eco107251, w_eco107252, w_eco107253, w_eco107254, w_eco107255, w_eco107256, w_eco107257, w_eco107258, w_eco107259, w_eco107260, w_eco107261, w_eco107262, w_eco107263, w_eco107264, w_eco107265, w_eco107266, w_eco107267, w_eco107268, w_eco107269, w_eco107270, w_eco107271, w_eco107272, w_eco107273, w_eco107274, w_eco107275, w_eco107276, w_eco107277, w_eco107278, w_eco107279, w_eco107280, w_eco107281, w_eco107282, w_eco107283, w_eco107284, w_eco107285, w_eco107286, w_eco107287, w_eco107288, w_eco107289, w_eco107290, w_eco107291, w_eco107292, w_eco107293, w_eco107294, w_eco107295, w_eco107296, w_eco107297, w_eco107298, w_eco107299, w_eco107300, w_eco107301, w_eco107302, w_eco107303, w_eco107304, w_eco107305, w_eco107306, w_eco107307, w_eco107308, w_eco107309, w_eco107310, w_eco107311, w_eco107312, w_eco107313, w_eco107314, w_eco107315, w_eco107316, w_eco107317, w_eco107318, w_eco107319, w_eco107320, w_eco107321, w_eco107322, w_eco107323, w_eco107324, w_eco107325, w_eco107326, w_eco107327, w_eco107328, w_eco107329, w_eco107330, w_eco107331, w_eco107332, w_eco107333, w_eco107334, w_eco107335, w_eco107336, w_eco107337, w_eco107338, w_eco107339, w_eco107340, w_eco107341, w_eco107342, w_eco107343, w_eco107344, w_eco107345, w_eco107346, w_eco107347, w_eco107348, w_eco107349, w_eco107350, w_eco107351, w_eco107352, w_eco107353, w_eco107354, w_eco107355, w_eco107356, w_eco107357, w_eco107358, w_eco107359, w_eco107360, w_eco107361, w_eco107362, w_eco107363, w_eco107364, w_eco107365, w_eco107366, w_eco107367, w_eco107368, w_eco107369, w_eco107370, w_eco107371, w_eco107372, w_eco107373, w_eco107374, w_eco107375, w_eco107376, w_eco107377, w_eco107378, w_eco107379, w_eco107380, w_eco107381, w_eco107382, w_eco107383, w_eco107384, w_eco107385, w_eco107386, w_eco107387, w_eco107388, w_eco107389, w_eco107390, w_eco107391, w_eco107392, w_eco107393, w_eco107394, w_eco107395, w_eco107396, w_eco107397, w_eco107398, w_eco107399, w_eco107400, w_eco107401, w_eco107402, w_eco107403, w_eco107404, w_eco107405, w_eco107406, w_eco107407, w_eco107408, w_eco107409, w_eco107410, w_eco107411, w_eco107412, w_eco107413, w_eco107414, w_eco107415, w_eco107416, w_eco107417, w_eco107418, w_eco107419, w_eco107420, w_eco107421, w_eco107422, w_eco107423, w_eco107424, w_eco107425, w_eco107426, w_eco107427, w_eco107428, w_eco107429, w_eco107430, w_eco107431, w_eco107432, w_eco107433, w_eco107434, w_eco107435, w_eco107436, w_eco107437, w_eco107438, w_eco107439, w_eco107440, w_eco107441, w_eco107442, w_eco107443, w_eco107444, w_eco107445, w_eco107446, w_eco107447, w_eco107448, w_eco107449, w_eco107450, w_eco107451, w_eco107452, w_eco107453, w_eco107454, w_eco107455, w_eco107456, w_eco107457, w_eco107458, w_eco107459, w_eco107460, w_eco107461, w_eco107462, w_eco107463, w_eco107464, w_eco107465, w_eco107466, w_eco107467, w_eco107468, w_eco107469, w_eco107470, w_eco107471, w_eco107472, w_eco107473, w_eco107474, w_eco107475, w_eco107476, w_eco107477, w_eco107478, w_eco107479, w_eco107480, w_eco107481, w_eco107482, w_eco107483, w_eco107484, w_eco107485, w_eco107486, w_eco107487, w_eco107488, w_eco107489, w_eco107490, w_eco107491, w_eco107492, w_eco107493, w_eco107494, w_eco107495, w_eco107496, w_eco107497, w_eco107498, w_eco107499, w_eco107500, w_eco107501, w_eco107502, w_eco107503, w_eco107504, w_eco107505, w_eco107506, w_eco107507, w_eco107508, w_eco107509, w_eco107510, w_eco107511, w_eco107512, w_eco107513, w_eco107514, w_eco107515, w_eco107516, w_eco107517, w_eco107518, w_eco107519, w_eco107520, w_eco107521, w_eco107522, w_eco107523, w_eco107524, w_eco107525, w_eco107526, w_eco107527, w_eco107528, w_eco107529, w_eco107530, w_eco107531, w_eco107532, w_eco107533, w_eco107534, w_eco107535, w_eco107536, w_eco107537, w_eco107538, w_eco107539, w_eco107540, w_eco107541, w_eco107542, w_eco107543, w_eco107544, w_eco107545, w_eco107546, w_eco107547, w_eco107548, w_eco107549, w_eco107550, w_eco107551, w_eco107552, w_eco107553, w_eco107554, w_eco107555, w_eco107556, w_eco107557, w_eco107558, w_eco107559, w_eco107560, w_eco107561, w_eco107562, w_eco107563, w_eco107564, w_eco107565, w_eco107566, w_eco107567, w_eco107568, w_eco107569, w_eco107570, w_eco107571, w_eco107572, w_eco107573, w_eco107574, w_eco107575, w_eco107576, w_eco107577, w_eco107578, w_eco107579, w_eco107580, w_eco107581, w_eco107582, w_eco107583, w_eco107584, w_eco107585, w_eco107586, w_eco107587, w_eco107588, w_eco107589, w_eco107590, w_eco107591, w_eco107592, w_eco107593, w_eco107594, w_eco107595, w_eco107596, w_eco107597, w_eco107598, w_eco107599, w_eco107600, w_eco107601, w_eco107602, w_eco107603, w_eco107604, w_eco107605, w_eco107606, w_eco107607, w_eco107608, w_eco107609, w_eco107610, w_eco107611, w_eco107612, w_eco107613, w_eco107614, w_eco107615, w_eco107616, w_eco107617, w_eco107618, w_eco107619, w_eco107620, w_eco107621, w_eco107622, w_eco107623, w_eco107624, w_eco107625, w_eco107626, w_eco107627, w_eco107628, w_eco107629, w_eco107630, w_eco107631, w_eco107632, w_eco107633, w_eco107634, w_eco107635, w_eco107636, w_eco107637, w_eco107638, w_eco107639, w_eco107640, w_eco107641, w_eco107642, w_eco107643, w_eco107644, w_eco107645, w_eco107646, w_eco107647, w_eco107648, w_eco107649, w_eco107650, w_eco107651, w_eco107652, w_eco107653, w_eco107654, w_eco107655, w_eco107656, w_eco107657, w_eco107658, w_eco107659, w_eco107660, w_eco107661, w_eco107662, w_eco107663, w_eco107664, w_eco107665, w_eco107666, w_eco107667, w_eco107668, w_eco107669, w_eco107670, w_eco107671, w_eco107672, w_eco107673, w_eco107674, w_eco107675, w_eco107676, w_eco107677, w_eco107678, w_eco107679, w_eco107680, w_eco107681, w_eco107682, w_eco107683, w_eco107684, w_eco107685, w_eco107686, w_eco107687, w_eco107688, w_eco107689, w_eco107690, w_eco107691, w_eco107692, w_eco107693, w_eco107694, w_eco107695, w_eco107696, w_eco107697, w_eco107698, w_eco107699, w_eco107700, w_eco107701, w_eco107702, w_eco107703, w_eco107704, w_eco107705, w_eco107706, w_eco107707, w_eco107708, w_eco107709, w_eco107710, w_eco107711, w_eco107712, w_eco107713, w_eco107714, w_eco107715, w_eco107716, w_eco107717, w_eco107718, w_eco107719, w_eco107720, w_eco107721, w_eco107722, w_eco107723, w_eco107724, w_eco107725, w_eco107726, w_eco107727, w_eco107728, w_eco107729, w_eco107730, w_eco107731, w_eco107732, w_eco107733, w_eco107734, w_eco107735, w_eco107736, w_eco107737, w_eco107738, w_eco107739, w_eco107740, w_eco107741, w_eco107742, w_eco107743, w_eco107744, w_eco107745, w_eco107746, w_eco107747, w_eco107748, w_eco107749, w_eco107750, w_eco107751, w_eco107752, w_eco107753, w_eco107754, w_eco107755, w_eco107756, w_eco107757, w_eco107758, w_eco107759, w_eco107760, w_eco107761, w_eco107762, w_eco107763, w_eco107764, w_eco107765, w_eco107766, w_eco107767, w_eco107768, w_eco107769, w_eco107770, w_eco107771, w_eco107772, w_eco107773, w_eco107774, w_eco107775, w_eco107776, w_eco107777, w_eco107778, w_eco107779, w_eco107780, w_eco107781, w_eco107782, w_eco107783, w_eco107784, w_eco107785, w_eco107786, w_eco107787, w_eco107788, w_eco107789, w_eco107790, w_eco107791, w_eco107792, w_eco107793, w_eco107794, w_eco107795, w_eco107796, w_eco107797, w_eco107798, w_eco107799, w_eco107800, w_eco107801, w_eco107802, w_eco107803, w_eco107804, w_eco107805, w_eco107806, w_eco107807, w_eco107808, w_eco107809, w_eco107810, w_eco107811, w_eco107812, w_eco107813, w_eco107814, w_eco107815, w_eco107816, w_eco107817, w_eco107818, w_eco107819, w_eco107820, w_eco107821, w_eco107822, w_eco107823, w_eco107824, w_eco107825, w_eco107826, w_eco107827, w_eco107828, w_eco107829, w_eco107830, w_eco107831, w_eco107832, w_eco107833, w_eco107834, w_eco107835, w_eco107836, w_eco107837, w_eco107838, w_eco107839, w_eco107840, w_eco107841, w_eco107842, w_eco107843, w_eco107844, w_eco107845, w_eco107846, w_eco107847, w_eco107848, w_eco107849, w_eco107850, w_eco107851, w_eco107852, w_eco107853, w_eco107854, w_eco107855, w_eco107856, w_eco107857, w_eco107858, w_eco107859, w_eco107860, w_eco107861, w_eco107862, w_eco107863, w_eco107864, w_eco107865, w_eco107866, w_eco107867, w_eco107868, w_eco107869, w_eco107870, w_eco107871, w_eco107872, w_eco107873, w_eco107874, w_eco107875, w_eco107876, w_eco107877, w_eco107878, w_eco107879, w_eco107880, w_eco107881, w_eco107882, w_eco107883, w_eco107884, w_eco107885, w_eco107886, w_eco107887, w_eco107888, w_eco107889, w_eco107890, w_eco107891, w_eco107892, w_eco107893, w_eco107894, w_eco107895, w_eco107896, w_eco107897, w_eco107898, w_eco107899, w_eco107900, w_eco107901, w_eco107902, w_eco107903, w_eco107904, w_eco107905, w_eco107906, w_eco107907, w_eco107908, w_eco107909, w_eco107910, w_eco107911, w_eco107912, w_eco107913, w_eco107914, w_eco107915, w_eco107916, w_eco107917, w_eco107918, w_eco107919, w_eco107920, w_eco107921, w_eco107922, w_eco107923, w_eco107924, w_eco107925, w_eco107926, w_eco107927, w_eco107928, w_eco107929, w_eco107930, w_eco107931, w_eco107932, w_eco107933, w_eco107934, w_eco107935, w_eco107936, w_eco107937, w_eco107938, w_eco107939, w_eco107940, w_eco107941, w_eco107942, w_eco107943, w_eco107944, w_eco107945, w_eco107946, w_eco107947, w_eco107948, w_eco107949, w_eco107950, w_eco107951, w_eco107952, w_eco107953, w_eco107954, w_eco107955, w_eco107956, w_eco107957, w_eco107958, w_eco107959, w_eco107960, w_eco107961, w_eco107962, w_eco107963, w_eco107964, w_eco107965, w_eco107966, w_eco107967, w_eco107968, w_eco107969, w_eco107970, w_eco107971, w_eco107972, w_eco107973, w_eco107974, w_eco107975, w_eco107976, w_eco107977, w_eco107978, w_eco107979, w_eco107980, w_eco107981, w_eco107982, w_eco107983, w_eco107984, w_eco107985, w_eco107986, w_eco107987, w_eco107988, w_eco107989, w_eco107990, w_eco107991, w_eco107992, w_eco107993, w_eco107994, w_eco107995, w_eco107996, w_eco107997, w_eco107998, w_eco107999, w_eco108000, w_eco108001, w_eco108002, w_eco108003, w_eco108004, w_eco108005, w_eco108006, w_eco108007, w_eco108008, w_eco108009, w_eco108010, w_eco108011, w_eco108012, w_eco108013, w_eco108014, w_eco108015, w_eco108016, w_eco108017, w_eco108018, w_eco108019, w_eco108020, w_eco108021, w_eco108022, w_eco108023, w_eco108024, w_eco108025, w_eco108026, w_eco108027, w_eco108028, w_eco108029, w_eco108030, w_eco108031, w_eco108032, w_eco108033, w_eco108034, w_eco108035, w_eco108036, w_eco108037, w_eco108038, w_eco108039, w_eco108040, w_eco108041, w_eco108042, w_eco108043, w_eco108044, w_eco108045, w_eco108046, w_eco108047, w_eco108048, w_eco108049, w_eco108050, w_eco108051, w_eco108052, w_eco108053, w_eco108054, w_eco108055, w_eco108056, w_eco108057, w_eco108058, w_eco108059, w_eco108060, w_eco108061, w_eco108062, w_eco108063, w_eco108064, w_eco108065, w_eco108066, w_eco108067, w_eco108068, w_eco108069, w_eco108070, w_eco108071, w_eco108072, w_eco108073, w_eco108074, w_eco108075, w_eco108076, w_eco108077, w_eco108078, w_eco108079, w_eco108080, w_eco108081, w_eco108082, w_eco108083, w_eco108084, w_eco108085, w_eco108086, w_eco108087, w_eco108088, w_eco108089, w_eco108090, w_eco108091, w_eco108092, w_eco108093, w_eco108094, w_eco108095, w_eco108096, w_eco108097, w_eco108098, w_eco108099, w_eco108100, w_eco108101, w_eco108102, w_eco108103, w_eco108104, w_eco108105, w_eco108106, w_eco108107, w_eco108108, w_eco108109, w_eco108110, w_eco108111, w_eco108112, w_eco108113, w_eco108114, w_eco108115, w_eco108116, w_eco108117, w_eco108118, w_eco108119, w_eco108120, w_eco108121, w_eco108122, w_eco108123, w_eco108124, w_eco108125, w_eco108126, w_eco108127, w_eco108128, w_eco108129, w_eco108130, w_eco108131, w_eco108132, w_eco108133, w_eco108134, w_eco108135, w_eco108136, w_eco108137, w_eco108138, w_eco108139, w_eco108140, w_eco108141, w_eco108142, w_eco108143, w_eco108144, w_eco108145, w_eco108146, w_eco108147, w_eco108148, w_eco108149, w_eco108150, w_eco108151, w_eco108152, w_eco108153, w_eco108154, w_eco108155, w_eco108156, w_eco108157, w_eco108158, w_eco108159, w_eco108160, w_eco108161, w_eco108162, w_eco108163, w_eco108164, w_eco108165, w_eco108166, w_eco108167, w_eco108168, w_eco108169, w_eco108170, w_eco108171, w_eco108172, w_eco108173, w_eco108174, w_eco108175, w_eco108176, w_eco108177, w_eco108178, w_eco108179, w_eco108180, w_eco108181, w_eco108182, w_eco108183, w_eco108184, w_eco108185, w_eco108186, w_eco108187, w_eco108188, w_eco108189, w_eco108190, w_eco108191, w_eco108192, w_eco108193, w_eco108194, w_eco108195, w_eco108196, w_eco108197, w_eco108198, w_eco108199, w_eco108200, w_eco108201, w_eco108202, w_eco108203, w_eco108204, w_eco108205, w_eco108206, w_eco108207, w_eco108208, w_eco108209, w_eco108210, w_eco108211, w_eco108212, w_eco108213, w_eco108214, w_eco108215, w_eco108216, w_eco108217, w_eco108218, w_eco108219, w_eco108220, w_eco108221, w_eco108222, w_eco108223, w_eco108224, w_eco108225, w_eco108226, w_eco108227, w_eco108228, w_eco108229, w_eco108230, w_eco108231, w_eco108232, w_eco108233, w_eco108234, w_eco108235, w_eco108236, w_eco108237, w_eco108238, w_eco108239, w_eco108240, w_eco108241, w_eco108242, w_eco108243, w_eco108244, w_eco108245, w_eco108246, w_eco108247, w_eco108248, w_eco108249, w_eco108250, w_eco108251, w_eco108252, w_eco108253, w_eco108254, w_eco108255, w_eco108256, w_eco108257, w_eco108258, w_eco108259, w_eco108260, w_eco108261, w_eco108262, w_eco108263, w_eco108264, w_eco108265, w_eco108266, w_eco108267, w_eco108268, w_eco108269, w_eco108270, w_eco108271, w_eco108272, w_eco108273, w_eco108274, w_eco108275, w_eco108276, w_eco108277, w_eco108278, w_eco108279, w_eco108280, w_eco108281, w_eco108282, w_eco108283, w_eco108284, w_eco108285, w_eco108286, w_eco108287, w_eco108288, w_eco108289, w_eco108290, w_eco108291, w_eco108292, w_eco108293, w_eco108294, w_eco108295, w_eco108296, w_eco108297, w_eco108298, w_eco108299, w_eco108300, w_eco108301, w_eco108302, w_eco108303, w_eco108304, w_eco108305, w_eco108306, w_eco108307, w_eco108308, w_eco108309, w_eco108310, w_eco108311, w_eco108312, w_eco108313, w_eco108314, w_eco108315, w_eco108316, w_eco108317, w_eco108318, w_eco108319, w_eco108320, w_eco108321, w_eco108322, w_eco108323, w_eco108324, w_eco108325, w_eco108326, w_eco108327, w_eco108328, w_eco108329, w_eco108330, w_eco108331, w_eco108332, w_eco108333, w_eco108334, w_eco108335, w_eco108336, w_eco108337, w_eco108338, w_eco108339, w_eco108340, w_eco108341, w_eco108342, w_eco108343, w_eco108344, w_eco108345, w_eco108346, w_eco108347, w_eco108348, w_eco108349, w_eco108350, w_eco108351, w_eco108352, w_eco108353, w_eco108354, w_eco108355, w_eco108356, w_eco108357, w_eco108358, w_eco108359, w_eco108360, w_eco108361, w_eco108362, w_eco108363, w_eco108364, w_eco108365, w_eco108366, w_eco108367, w_eco108368, w_eco108369, w_eco108370, w_eco108371, w_eco108372, w_eco108373, w_eco108374, w_eco108375, w_eco108376, w_eco108377, w_eco108378, w_eco108379, w_eco108380, w_eco108381, w_eco108382, w_eco108383, w_eco108384, w_eco108385, w_eco108386, w_eco108387, w_eco108388, w_eco108389, w_eco108390, w_eco108391, w_eco108392, w_eco108393, w_eco108394, w_eco108395, w_eco108396, w_eco108397, w_eco108398, w_eco108399, w_eco108400, w_eco108401, w_eco108402, w_eco108403, w_eco108404, w_eco108405, w_eco108406, w_eco108407, w_eco108408, w_eco108409, w_eco108410, w_eco108411, w_eco108412, w_eco108413, w_eco108414, w_eco108415, w_eco108416, w_eco108417, w_eco108418, w_eco108419, w_eco108420, w_eco108421, w_eco108422, w_eco108423, w_eco108424, w_eco108425, w_eco108426, w_eco108427, w_eco108428, w_eco108429, w_eco108430, w_eco108431, w_eco108432, w_eco108433, w_eco108434, w_eco108435, w_eco108436, w_eco108437, w_eco108438, w_eco108439, w_eco108440, w_eco108441, w_eco108442, w_eco108443, w_eco108444, w_eco108445, w_eco108446, w_eco108447, w_eco108448, w_eco108449, w_eco108450, w_eco108451, w_eco108452, w_eco108453, w_eco108454, w_eco108455, w_eco108456, w_eco108457, w_eco108458, w_eco108459, w_eco108460, w_eco108461, w_eco108462, w_eco108463, w_eco108464, w_eco108465, w_eco108466, w_eco108467, w_eco108468, w_eco108469, w_eco108470, w_eco108471, w_eco108472, w_eco108473, w_eco108474, w_eco108475, w_eco108476, w_eco108477, w_eco108478, w_eco108479, w_eco108480, w_eco108481, w_eco108482, w_eco108483, w_eco108484, w_eco108485, w_eco108486, w_eco108487, w_eco108488, w_eco108489, w_eco108490, w_eco108491, w_eco108492, w_eco108493, w_eco108494, w_eco108495, w_eco108496, w_eco108497, w_eco108498, w_eco108499, w_eco108500, w_eco108501, w_eco108502, w_eco108503, w_eco108504, w_eco108505, w_eco108506, w_eco108507, w_eco108508, w_eco108509, w_eco108510, w_eco108511, w_eco108512, w_eco108513, w_eco108514, w_eco108515, w_eco108516, w_eco108517, w_eco108518, w_eco108519, w_eco108520, w_eco108521, w_eco108522, w_eco108523, w_eco108524, w_eco108525, w_eco108526, w_eco108527, w_eco108528, w_eco108529, w_eco108530, w_eco108531, w_eco108532, w_eco108533, w_eco108534, w_eco108535, w_eco108536, w_eco108537, w_eco108538, w_eco108539, w_eco108540, w_eco108541, w_eco108542, w_eco108543, w_eco108544, w_eco108545, w_eco108546, w_eco108547, w_eco108548, w_eco108549, w_eco108550, w_eco108551, w_eco108552, w_eco108553, w_eco108554, w_eco108555, w_eco108556, w_eco108557, w_eco108558, w_eco108559, w_eco108560, w_eco108561, w_eco108562, w_eco108563, w_eco108564, w_eco108565, w_eco108566, w_eco108567, w_eco108568, w_eco108569, w_eco108570, w_eco108571, w_eco108572, w_eco108573, w_eco108574, w_eco108575, w_eco108576, w_eco108577, w_eco108578, w_eco108579, w_eco108580, w_eco108581, w_eco108582, w_eco108583, w_eco108584, w_eco108585, w_eco108586, w_eco108587, w_eco108588, w_eco108589, w_eco108590, w_eco108591, w_eco108592, w_eco108593, w_eco108594, w_eco108595, w_eco108596, w_eco108597, w_eco108598, w_eco108599, w_eco108600, w_eco108601, w_eco108602, w_eco108603, w_eco108604, w_eco108605, w_eco108606, w_eco108607, w_eco108608, w_eco108609, w_eco108610, w_eco108611, w_eco108612, w_eco108613, w_eco108614, w_eco108615, w_eco108616, w_eco108617, w_eco108618, w_eco108619, w_eco108620, w_eco108621, w_eco108622, w_eco108623, w_eco108624, w_eco108625, w_eco108626, w_eco108627, w_eco108628, w_eco108629, w_eco108630, w_eco108631, w_eco108632, w_eco108633, w_eco108634, w_eco108635, w_eco108636, w_eco108637, w_eco108638, w_eco108639, w_eco108640, w_eco108641, w_eco108642, w_eco108643, w_eco108644, w_eco108645, w_eco108646, w_eco108647, w_eco108648, w_eco108649, w_eco108650, w_eco108651, w_eco108652, w_eco108653, w_eco108654, w_eco108655, w_eco108656, w_eco108657, w_eco108658, w_eco108659, w_eco108660, w_eco108661, w_eco108662, w_eco108663, w_eco108664, w_eco108665, w_eco108666, w_eco108667, w_eco108668, w_eco108669, w_eco108670, w_eco108671, w_eco108672, w_eco108673, w_eco108674, w_eco108675, w_eco108676, w_eco108677, w_eco108678, w_eco108679, w_eco108680, w_eco108681, w_eco108682, w_eco108683, w_eco108684, w_eco108685, w_eco108686, w_eco108687, w_eco108688, w_eco108689, w_eco108690, w_eco108691, w_eco108692, w_eco108693, w_eco108694, w_eco108695, w_eco108696, w_eco108697, w_eco108698, w_eco108699, w_eco108700, w_eco108701, w_eco108702, w_eco108703, w_eco108704, w_eco108705, w_eco108706, w_eco108707, w_eco108708, w_eco108709, w_eco108710, w_eco108711, w_eco108712, w_eco108713, w_eco108714, w_eco108715, w_eco108716, w_eco108717, w_eco108718, w_eco108719, w_eco108720, w_eco108721, w_eco108722, w_eco108723, w_eco108724, w_eco108725, w_eco108726, w_eco108727, w_eco108728, w_eco108729, w_eco108730, w_eco108731, w_eco108732, w_eco108733, w_eco108734, w_eco108735, w_eco108736, w_eco108737, w_eco108738, w_eco108739, w_eco108740, w_eco108741, w_eco108742, w_eco108743, w_eco108744, w_eco108745, w_eco108746, w_eco108747, w_eco108748, w_eco108749, w_eco108750, w_eco108751, w_eco108752, w_eco108753, w_eco108754, w_eco108755, w_eco108756, w_eco108757, w_eco108758, w_eco108759, w_eco108760, w_eco108761, w_eco108762, w_eco108763, w_eco108764, w_eco108765, w_eco108766, w_eco108767, w_eco108768, w_eco108769, w_eco108770, w_eco108771, w_eco108772, w_eco108773, w_eco108774, w_eco108775, w_eco108776, w_eco108777, w_eco108778, w_eco108779, w_eco108780, w_eco108781, w_eco108782, w_eco108783, w_eco108784, w_eco108785, w_eco108786, w_eco108787, w_eco108788, w_eco108789, w_eco108790, w_eco108791, w_eco108792, w_eco108793, w_eco108794, w_eco108795, w_eco108796, w_eco108797, w_eco108798, w_eco108799, w_eco108800, w_eco108801, w_eco108802, w_eco108803, w_eco108804, w_eco108805, w_eco108806, w_eco108807, w_eco108808, w_eco108809, w_eco108810, w_eco108811, w_eco108812, w_eco108813, w_eco108814, w_eco108815, w_eco108816, w_eco108817, w_eco108818, w_eco108819, w_eco108820, w_eco108821, w_eco108822, w_eco108823, w_eco108824, w_eco108825, w_eco108826, w_eco108827, w_eco108828, w_eco108829, w_eco108830, w_eco108831, w_eco108832, w_eco108833, w_eco108834, w_eco108835, w_eco108836, w_eco108837, w_eco108838, w_eco108839, w_eco108840, w_eco108841, w_eco108842, w_eco108843, w_eco108844, w_eco108845, w_eco108846, w_eco108847, w_eco108848, w_eco108849, w_eco108850, w_eco108851, w_eco108852, w_eco108853, w_eco108854, w_eco108855, w_eco108856, w_eco108857, w_eco108858, w_eco108859, w_eco108860, w_eco108861, w_eco108862, w_eco108863, w_eco108864, w_eco108865, w_eco108866, w_eco108867, w_eco108868, w_eco108869, w_eco108870, w_eco108871, w_eco108872, w_eco108873, w_eco108874, w_eco108875, w_eco108876, w_eco108877, w_eco108878, w_eco108879, w_eco108880, w_eco108881, w_eco108882, w_eco108883, w_eco108884, w_eco108885, w_eco108886, w_eco108887, w_eco108888, w_eco108889, w_eco108890, w_eco108891, w_eco108892, w_eco108893, w_eco108894, w_eco108895, w_eco108896, w_eco108897, w_eco108898, w_eco108899, w_eco108900, w_eco108901, w_eco108902, w_eco108903, w_eco108904, w_eco108905, w_eco108906, w_eco108907, w_eco108908, w_eco108909, w_eco108910, w_eco108911, w_eco108912, w_eco108913, w_eco108914, w_eco108915, w_eco108916, w_eco108917, w_eco108918, w_eco108919, w_eco108920, w_eco108921, w_eco108922, w_eco108923, w_eco108924, w_eco108925, w_eco108926, w_eco108927, w_eco108928, w_eco108929, w_eco108930, w_eco108931, w_eco108932, w_eco108933, w_eco108934, w_eco108935, w_eco108936, w_eco108937, w_eco108938, w_eco108939, w_eco108940, w_eco108941, w_eco108942, w_eco108943, w_eco108944, w_eco108945, w_eco108946, w_eco108947, w_eco108948, w_eco108949, w_eco108950, w_eco108951, w_eco108952, w_eco108953, w_eco108954, w_eco108955, w_eco108956, w_eco108957, w_eco108958, w_eco108959, w_eco108960, w_eco108961, w_eco108962, w_eco108963, w_eco108964, w_eco108965, w_eco108966, w_eco108967, w_eco108968, w_eco108969, w_eco108970, w_eco108971, w_eco108972, w_eco108973, w_eco108974, w_eco108975, w_eco108976, w_eco108977, w_eco108978, w_eco108979, w_eco108980, w_eco108981, w_eco108982, w_eco108983, w_eco108984, w_eco108985, w_eco108986, w_eco108987, w_eco108988, w_eco108989, w_eco108990, w_eco108991, w_eco108992, w_eco108993, w_eco108994, w_eco108995, w_eco108996, w_eco108997, w_eco108998, w_eco108999, w_eco109000, w_eco109001, w_eco109002, w_eco109003, w_eco109004, w_eco109005, w_eco109006, w_eco109007, w_eco109008, w_eco109009, w_eco109010, w_eco109011, w_eco109012, w_eco109013, w_eco109014, w_eco109015, w_eco109016, w_eco109017, w_eco109018, w_eco109019, w_eco109020, w_eco109021, w_eco109022, w_eco109023, w_eco109024, w_eco109025, w_eco109026, w_eco109027, w_eco109028, w_eco109029, w_eco109030, w_eco109031, w_eco109032, w_eco109033, w_eco109034, w_eco109035, w_eco109036, w_eco109037, w_eco109038, w_eco109039, w_eco109040, w_eco109041, w_eco109042, w_eco109043, w_eco109044, w_eco109045, w_eco109046, w_eco109047, w_eco109048, w_eco109049, w_eco109050, w_eco109051, w_eco109052, w_eco109053, w_eco109054, w_eco109055, w_eco109056, w_eco109057, w_eco109058, w_eco109059, w_eco109060, w_eco109061, w_eco109062, w_eco109063, w_eco109064, w_eco109065, w_eco109066, w_eco109067, w_eco109068, w_eco109069, w_eco109070, w_eco109071, w_eco109072, w_eco109073, w_eco109074, w_eco109075, w_eco109076, w_eco109077, w_eco109078, w_eco109079, w_eco109080, w_eco109081, w_eco109082, w_eco109083, w_eco109084, w_eco109085, w_eco109086, w_eco109087, w_eco109088, w_eco109089, w_eco109090, w_eco109091, w_eco109092, w_eco109093, w_eco109094, w_eco109095, w_eco109096, w_eco109097, w_eco109098, w_eco109099, w_eco109100, w_eco109101, w_eco109102, w_eco109103, w_eco109104, w_eco109105, w_eco109106, w_eco109107, w_eco109108, w_eco109109, w_eco109110, w_eco109111, w_eco109112, w_eco109113, w_eco109114, w_eco109115, w_eco109116, w_eco109117, w_eco109118, w_eco109119, w_eco109120, w_eco109121, w_eco109122, w_eco109123, w_eco109124, w_eco109125, w_eco109126, w_eco109127, w_eco109128, w_eco109129, w_eco109130, w_eco109131, w_eco109132, w_eco109133, w_eco109134, w_eco109135, w_eco109136, w_eco109137, w_eco109138, w_eco109139, w_eco109140, w_eco109141, w_eco109142, w_eco109143, w_eco109144, w_eco109145, w_eco109146, w_eco109147, w_eco109148, w_eco109149, w_eco109150, w_eco109151, w_eco109152, w_eco109153, w_eco109154, w_eco109155, w_eco109156, w_eco109157, w_eco109158, w_eco109159, w_eco109160, w_eco109161, w_eco109162, w_eco109163, w_eco109164, w_eco109165, w_eco109166, w_eco109167, w_eco109168, w_eco109169, w_eco109170, w_eco109171, w_eco109172, w_eco109173, w_eco109174, w_eco109175, w_eco109176, w_eco109177, w_eco109178, w_eco109179, w_eco109180, w_eco109181, w_eco109182, w_eco109183, w_eco109184, w_eco109185, w_eco109186, w_eco109187, w_eco109188, w_eco109189, w_eco109190, w_eco109191, w_eco109192, w_eco109193, w_eco109194, w_eco109195, w_eco109196, w_eco109197, w_eco109198, w_eco109199, w_eco109200, w_eco109201, w_eco109202, w_eco109203, w_eco109204, w_eco109205, w_eco109206, w_eco109207, w_eco109208, w_eco109209, w_eco109210, w_eco109211, w_eco109212, w_eco109213, w_eco109214, w_eco109215, w_eco109216, w_eco109217, w_eco109218, w_eco109219, w_eco109220, w_eco109221, w_eco109222, w_eco109223, w_eco109224, w_eco109225, w_eco109226, w_eco109227, w_eco109228, w_eco109229, w_eco109230, w_eco109231, w_eco109232, w_eco109233, w_eco109234, w_eco109235, w_eco109236, w_eco109237, w_eco109238, w_eco109239, w_eco109240, w_eco109241, w_eco109242, w_eco109243, w_eco109244, w_eco109245, w_eco109246, w_eco109247, w_eco109248, w_eco109249, w_eco109250, w_eco109251, w_eco109252, w_eco109253, w_eco109254, w_eco109255, w_eco109256, w_eco109257, w_eco109258, w_eco109259, w_eco109260, w_eco109261, w_eco109262, w_eco109263, w_eco109264, w_eco109265, w_eco109266, w_eco109267, w_eco109268, w_eco109269, w_eco109270, w_eco109271, w_eco109272, w_eco109273, w_eco109274, w_eco109275, w_eco109276, w_eco109277, w_eco109278, w_eco109279, w_eco109280, w_eco109281, w_eco109282, w_eco109283, w_eco109284, w_eco109285, w_eco109286, w_eco109287, w_eco109288, w_eco109289, w_eco109290, w_eco109291, w_eco109292, w_eco109293, w_eco109294, w_eco109295, w_eco109296, w_eco109297, w_eco109298, w_eco109299, w_eco109300, w_eco109301, w_eco109302, w_eco109303, w_eco109304, w_eco109305, w_eco109306, w_eco109307, w_eco109308, w_eco109309, w_eco109310, w_eco109311, w_eco109312, w_eco109313, w_eco109314, w_eco109315, w_eco109316, w_eco109317, w_eco109318, w_eco109319, w_eco109320, w_eco109321, w_eco109322, w_eco109323, w_eco109324, w_eco109325, w_eco109326, w_eco109327, w_eco109328, w_eco109329, w_eco109330, w_eco109331, w_eco109332, w_eco109333, w_eco109334, w_eco109335, w_eco109336, w_eco109337, w_eco109338, w_eco109339, w_eco109340, w_eco109341, w_eco109342, w_eco109343, w_eco109344, w_eco109345, w_eco109346, w_eco109347, w_eco109348, w_eco109349, w_eco109350, w_eco109351, w_eco109352, w_eco109353, w_eco109354, w_eco109355, w_eco109356, w_eco109357, w_eco109358, w_eco109359, w_eco109360, w_eco109361, w_eco109362, w_eco109363, w_eco109364, w_eco109365, w_eco109366, w_eco109367, w_eco109368, w_eco109369, w_eco109370, w_eco109371, w_eco109372, w_eco109373, w_eco109374, w_eco109375, w_eco109376, w_eco109377, w_eco109378, w_eco109379, w_eco109380, w_eco109381, w_eco109382, w_eco109383, w_eco109384, w_eco109385, w_eco109386, w_eco109387, w_eco109388, w_eco109389, w_eco109390, w_eco109391, w_eco109392, w_eco109393, w_eco109394, w_eco109395, w_eco109396, w_eco109397, w_eco109398, w_eco109399, w_eco109400, w_eco109401, w_eco109402, w_eco109403, w_eco109404, w_eco109405, w_eco109406, w_eco109407, w_eco109408, w_eco109409, w_eco109410, w_eco109411, w_eco109412, w_eco109413, w_eco109414, w_eco109415, w_eco109416, w_eco109417, w_eco109418, w_eco109419, w_eco109420, w_eco109421, w_eco109422, w_eco109423, w_eco109424, w_eco109425, w_eco109426, w_eco109427, w_eco109428, w_eco109429, w_eco109430, w_eco109431, w_eco109432, w_eco109433, w_eco109434, w_eco109435, w_eco109436, w_eco109437, w_eco109438, w_eco109439, w_eco109440, w_eco109441, w_eco109442, w_eco109443, w_eco109444, w_eco109445, w_eco109446, w_eco109447, w_eco109448, w_eco109449, w_eco109450, w_eco109451, w_eco109452, w_eco109453, w_eco109454, w_eco109455, w_eco109456, w_eco109457, w_eco109458, w_eco109459, w_eco109460, w_eco109461, w_eco109462, w_eco109463, w_eco109464, w_eco109465, w_eco109466, w_eco109467, w_eco109468, w_eco109469, w_eco109470, w_eco109471, w_eco109472, w_eco109473, w_eco109474, w_eco109475, w_eco109476, w_eco109477, w_eco109478, w_eco109479, w_eco109480, w_eco109481, w_eco109482, w_eco109483, w_eco109484, w_eco109485, w_eco109486, w_eco109487, w_eco109488, w_eco109489, w_eco109490, w_eco109491, w_eco109492, w_eco109493, w_eco109494, w_eco109495, w_eco109496, w_eco109497, w_eco109498, w_eco109499, w_eco109500, w_eco109501, w_eco109502, w_eco109503, w_eco109504, w_eco109505, w_eco109506, w_eco109507, w_eco109508, w_eco109509, w_eco109510, w_eco109511, w_eco109512, w_eco109513, w_eco109514, w_eco109515, w_eco109516, w_eco109517, w_eco109518, w_eco109519, w_eco109520, w_eco109521, w_eco109522, w_eco109523, w_eco109524, w_eco109525, w_eco109526, w_eco109527, w_eco109528, w_eco109529, w_eco109530, w_eco109531, w_eco109532, w_eco109533, w_eco109534, w_eco109535, w_eco109536, w_eco109537, w_eco109538, w_eco109539, w_eco109540, w_eco109541, w_eco109542, w_eco109543, w_eco109544, w_eco109545, w_eco109546, w_eco109547, w_eco109548, w_eco109549, w_eco109550, w_eco109551, w_eco109552, w_eco109553, w_eco109554, w_eco109555, w_eco109556, w_eco109557, w_eco109558, w_eco109559, w_eco109560, w_eco109561, w_eco109562, w_eco109563, w_eco109564, w_eco109565, w_eco109566, w_eco109567, w_eco109568, w_eco109569, w_eco109570, w_eco109571, w_eco109572, w_eco109573, w_eco109574, w_eco109575, w_eco109576, w_eco109577, w_eco109578, w_eco109579, w_eco109580, w_eco109581, w_eco109582, w_eco109583, w_eco109584, w_eco109585, w_eco109586, w_eco109587, w_eco109588, w_eco109589, w_eco109590, w_eco109591, w_eco109592, w_eco109593, w_eco109594, w_eco109595, w_eco109596, w_eco109597, w_eco109598, w_eco109599, w_eco109600, w_eco109601, w_eco109602, w_eco109603, w_eco109604, w_eco109605, w_eco109606, w_eco109607, w_eco109608, w_eco109609, w_eco109610, w_eco109611, w_eco109612, w_eco109613, w_eco109614, w_eco109615, w_eco109616, w_eco109617, w_eco109618, w_eco109619, w_eco109620, w_eco109621, w_eco109622, w_eco109623, w_eco109624, w_eco109625, w_eco109626, w_eco109627, w_eco109628, w_eco109629, w_eco109630, w_eco109631, w_eco109632, w_eco109633, w_eco109634, w_eco109635, w_eco109636, w_eco109637, w_eco109638, w_eco109639, w_eco109640, w_eco109641, w_eco109642, w_eco109643, w_eco109644, w_eco109645, w_eco109646, w_eco109647, w_eco109648, w_eco109649, w_eco109650, w_eco109651, w_eco109652, w_eco109653, w_eco109654, w_eco109655, w_eco109656, w_eco109657, w_eco109658, w_eco109659, w_eco109660, w_eco109661, w_eco109662, w_eco109663, w_eco109664, w_eco109665, w_eco109666, w_eco109667, w_eco109668, w_eco109669, w_eco109670, w_eco109671, w_eco109672, w_eco109673, w_eco109674, w_eco109675, w_eco109676, w_eco109677, w_eco109678, w_eco109679, w_eco109680, w_eco109681, w_eco109682, w_eco109683, w_eco109684, w_eco109685, w_eco109686, w_eco109687, w_eco109688, w_eco109689, w_eco109690, w_eco109691, w_eco109692, w_eco109693, w_eco109694, w_eco109695, w_eco109696, w_eco109697, w_eco109698, w_eco109699, w_eco109700, w_eco109701, w_eco109702, w_eco109703, w_eco109704, w_eco109705, w_eco109706, w_eco109707, w_eco109708, w_eco109709, w_eco109710, w_eco109711, w_eco109712, w_eco109713, w_eco109714, w_eco109715, w_eco109716, w_eco109717, w_eco109718, w_eco109719, w_eco109720, w_eco109721, w_eco109722, w_eco109723, w_eco109724, w_eco109725, w_eco109726, w_eco109727, w_eco109728, w_eco109729, w_eco109730, w_eco109731, w_eco109732, w_eco109733, w_eco109734, w_eco109735, w_eco109736, w_eco109737, w_eco109738, w_eco109739, w_eco109740, w_eco109741, w_eco109742, w_eco109743, w_eco109744, w_eco109745, w_eco109746, w_eco109747, w_eco109748, w_eco109749, w_eco109750, w_eco109751, w_eco109752, w_eco109753, w_eco109754, w_eco109755, w_eco109756, w_eco109757, w_eco109758, w_eco109759, w_eco109760, w_eco109761, w_eco109762, w_eco109763, w_eco109764, w_eco109765, w_eco109766, w_eco109767, w_eco109768, w_eco109769, w_eco109770, w_eco109771, w_eco109772, w_eco109773, w_eco109774, w_eco109775, w_eco109776, w_eco109777, w_eco109778, w_eco109779, w_eco109780, w_eco109781, w_eco109782, w_eco109783, w_eco109784, w_eco109785, w_eco109786, w_eco109787, w_eco109788, w_eco109789, w_eco109790, w_eco109791, w_eco109792, w_eco109793, w_eco109794, w_eco109795, w_eco109796, w_eco109797, w_eco109798, w_eco109799, w_eco109800, w_eco109801, w_eco109802, w_eco109803, w_eco109804, w_eco109805, w_eco109806, w_eco109807, w_eco109808, w_eco109809, w_eco109810, w_eco109811, w_eco109812, w_eco109813, w_eco109814, w_eco109815, w_eco109816, w_eco109817, w_eco109818, w_eco109819, w_eco109820, w_eco109821, w_eco109822, w_eco109823, w_eco109824, w_eco109825, w_eco109826, w_eco109827, w_eco109828, w_eco109829, w_eco109830, w_eco109831, w_eco109832, w_eco109833, w_eco109834, w_eco109835, w_eco109836, w_eco109837, w_eco109838, w_eco109839, w_eco109840, w_eco109841, w_eco109842, w_eco109843, w_eco109844, w_eco109845, w_eco109846, w_eco109847, w_eco109848, w_eco109849, w_eco109850, w_eco109851, w_eco109852, w_eco109853, w_eco109854, w_eco109855, w_eco109856, w_eco109857, w_eco109858, w_eco109859, w_eco109860, w_eco109861, w_eco109862, w_eco109863, w_eco109864, w_eco109865, w_eco109866, w_eco109867, w_eco109868, w_eco109869, w_eco109870, w_eco109871, w_eco109872, w_eco109873, w_eco109874, w_eco109875, w_eco109876, w_eco109877, w_eco109878, w_eco109879, w_eco109880, w_eco109881, w_eco109882, w_eco109883, w_eco109884, w_eco109885, w_eco109886, w_eco109887, w_eco109888, w_eco109889, w_eco109890, w_eco109891, w_eco109892, w_eco109893, w_eco109894, w_eco109895, w_eco109896, w_eco109897, w_eco109898, w_eco109899, w_eco109900, w_eco109901, w_eco109902, w_eco109903, w_eco109904, w_eco109905, w_eco109906, w_eco109907, w_eco109908, w_eco109909, w_eco109910, w_eco109911, w_eco109912, w_eco109913, w_eco109914, w_eco109915, w_eco109916, w_eco109917, w_eco109918, w_eco109919, w_eco109920, w_eco109921, w_eco109922, w_eco109923, w_eco109924, w_eco109925, w_eco109926, w_eco109927, w_eco109928, w_eco109929, w_eco109930, w_eco109931, w_eco109932, w_eco109933, w_eco109934, w_eco109935, w_eco109936, w_eco109937, w_eco109938, w_eco109939, w_eco109940, w_eco109941, w_eco109942, w_eco109943, w_eco109944, w_eco109945, w_eco109946, w_eco109947, w_eco109948, w_eco109949, w_eco109950, w_eco109951, w_eco109952, w_eco109953, w_eco109954, w_eco109955, w_eco109956, w_eco109957, w_eco109958, w_eco109959, w_eco109960, w_eco109961, w_eco109962, w_eco109963, w_eco109964, w_eco109965, w_eco109966, w_eco109967, w_eco109968, w_eco109969, w_eco109970, w_eco109971, w_eco109972, w_eco109973, w_eco109974, w_eco109975, w_eco109976, w_eco109977, w_eco109978, w_eco109979, w_eco109980, w_eco109981, w_eco109982, w_eco109983, w_eco109984, w_eco109985, w_eco109986, w_eco109987, w_eco109988, w_eco109989, w_eco109990, w_eco109991, w_eco109992, w_eco109993, w_eco109994, w_eco109995, w_eco109996, w_eco109997, w_eco109998, w_eco109999, w_eco110000, w_eco110001, w_eco110002, w_eco110003, w_eco110004, w_eco110005, w_eco110006, w_eco110007, w_eco110008, w_eco110009, w_eco110010, w_eco110011, w_eco110012, w_eco110013, w_eco110014, w_eco110015, w_eco110016, w_eco110017, w_eco110018, w_eco110019, w_eco110020, w_eco110021, w_eco110022, w_eco110023, w_eco110024, w_eco110025, w_eco110026, w_eco110027, w_eco110028, w_eco110029, w_eco110030, w_eco110031, w_eco110032, w_eco110033, w_eco110034, w_eco110035, w_eco110036, w_eco110037, w_eco110038, w_eco110039, w_eco110040, w_eco110041, w_eco110042, w_eco110043, w_eco110044, w_eco110045, w_eco110046, w_eco110047, w_eco110048, w_eco110049, w_eco110050, w_eco110051, w_eco110052, w_eco110053, w_eco110054, w_eco110055, w_eco110056, w_eco110057, w_eco110058, w_eco110059, w_eco110060, w_eco110061, w_eco110062, w_eco110063, w_eco110064, w_eco110065, w_eco110066, w_eco110067, w_eco110068, w_eco110069, w_eco110070, w_eco110071, w_eco110072, w_eco110073, w_eco110074, w_eco110075, w_eco110076, w_eco110077, w_eco110078, w_eco110079, w_eco110080, w_eco110081, w_eco110082, w_eco110083, w_eco110084, w_eco110085, w_eco110086, w_eco110087, w_eco110088, w_eco110089, w_eco110090, w_eco110091, w_eco110092, w_eco110093, w_eco110094, w_eco110095, w_eco110096, w_eco110097, w_eco110098, w_eco110099, w_eco110100, w_eco110101, w_eco110102, w_eco110103, w_eco110104, w_eco110105, w_eco110106, w_eco110107, w_eco110108, w_eco110109, w_eco110110, w_eco110111, w_eco110112, w_eco110113, w_eco110114, w_eco110115, w_eco110116, w_eco110117, w_eco110118, w_eco110119, w_eco110120, w_eco110121, w_eco110122, w_eco110123, w_eco110124, w_eco110125, w_eco110126, w_eco110127, w_eco110128, w_eco110129, w_eco110130, w_eco110131, w_eco110132, w_eco110133, w_eco110134, w_eco110135, w_eco110136, w_eco110137, w_eco110138, w_eco110139, w_eco110140, w_eco110141, w_eco110142, w_eco110143, w_eco110144, w_eco110145, w_eco110146, w_eco110147, w_eco110148, w_eco110149, w_eco110150, w_eco110151, w_eco110152, w_eco110153, w_eco110154, w_eco110155, w_eco110156, w_eco110157, w_eco110158, w_eco110159, w_eco110160, w_eco110161, w_eco110162, w_eco110163, w_eco110164, w_eco110165, w_eco110166, w_eco110167, w_eco110168, w_eco110169, w_eco110170, w_eco110171, w_eco110172, w_eco110173, w_eco110174, w_eco110175, w_eco110176, w_eco110177, w_eco110178, w_eco110179, w_eco110180, w_eco110181, w_eco110182, w_eco110183, w_eco110184, w_eco110185, w_eco110186, w_eco110187, w_eco110188, w_eco110189, w_eco110190, w_eco110191, w_eco110192, w_eco110193, w_eco110194, w_eco110195, w_eco110196, w_eco110197, w_eco110198, w_eco110199, w_eco110200, w_eco110201, w_eco110202, w_eco110203, w_eco110204, w_eco110205, w_eco110206, w_eco110207, w_eco110208, w_eco110209, w_eco110210, w_eco110211, w_eco110212, w_eco110213, w_eco110214, w_eco110215, w_eco110216, w_eco110217, w_eco110218, w_eco110219, w_eco110220, w_eco110221, w_eco110222, w_eco110223, w_eco110224, w_eco110225, w_eco110226, w_eco110227, w_eco110228, w_eco110229, w_eco110230, w_eco110231, w_eco110232, w_eco110233, w_eco110234, w_eco110235, w_eco110236, w_eco110237, w_eco110238, w_eco110239, w_eco110240, w_eco110241, w_eco110242, w_eco110243, w_eco110244, w_eco110245, w_eco110246, w_eco110247, w_eco110248, w_eco110249, w_eco110250, w_eco110251, w_eco110252, w_eco110253, w_eco110254, w_eco110255, w_eco110256, w_eco110257, w_eco110258, w_eco110259, w_eco110260, w_eco110261, w_eco110262, w_eco110263, w_eco110264, w_eco110265, w_eco110266, w_eco110267, w_eco110268, w_eco110269, w_eco110270, w_eco110271, w_eco110272, w_eco110273, w_eco110274, w_eco110275, w_eco110276, w_eco110277, w_eco110278, w_eco110279, w_eco110280, w_eco110281, w_eco110282, w_eco110283, w_eco110284, w_eco110285, w_eco110286, w_eco110287, w_eco110288, w_eco110289, w_eco110290, w_eco110291, w_eco110292, w_eco110293, w_eco110294, w_eco110295, w_eco110296, w_eco110297, w_eco110298, w_eco110299, w_eco110300, w_eco110301, w_eco110302, w_eco110303, w_eco110304, w_eco110305, w_eco110306, w_eco110307, w_eco110308, w_eco110309, w_eco110310, w_eco110311, w_eco110312, w_eco110313, w_eco110314, w_eco110315, w_eco110316, w_eco110317, w_eco110318, w_eco110319, w_eco110320, w_eco110321, w_eco110322, w_eco110323, w_eco110324, w_eco110325, w_eco110326, w_eco110327, w_eco110328, w_eco110329, w_eco110330, w_eco110331, w_eco110332, w_eco110333, w_eco110334, w_eco110335, w_eco110336, w_eco110337, w_eco110338, w_eco110339, w_eco110340, w_eco110341, w_eco110342, w_eco110343, w_eco110344, w_eco110345, w_eco110346, w_eco110347, w_eco110348, w_eco110349, w_eco110350, w_eco110351, w_eco110352, w_eco110353, w_eco110354, w_eco110355, w_eco110356, w_eco110357, w_eco110358, w_eco110359, w_eco110360, w_eco110361, w_eco110362, w_eco110363, w_eco110364, w_eco110365, w_eco110366, w_eco110367, w_eco110368, w_eco110369, w_eco110370, w_eco110371, w_eco110372, w_eco110373, w_eco110374, w_eco110375, w_eco110376, w_eco110377, w_eco110378, w_eco110379, w_eco110380, w_eco110381, w_eco110382, w_eco110383, w_eco110384, w_eco110385, w_eco110386, w_eco110387, w_eco110388, w_eco110389, w_eco110390, w_eco110391, w_eco110392, w_eco110393, w_eco110394, w_eco110395, w_eco110396, w_eco110397, w_eco110398, w_eco110399, w_eco110400, w_eco110401, w_eco110402, w_eco110403, w_eco110404, w_eco110405, w_eco110406, w_eco110407, w_eco110408, w_eco110409, w_eco110410, w_eco110411, w_eco110412, w_eco110413, w_eco110414, w_eco110415, w_eco110416, w_eco110417, w_eco110418, w_eco110419, w_eco110420, w_eco110421, w_eco110422, w_eco110423, w_eco110424, w_eco110425, w_eco110426, w_eco110427, w_eco110428, w_eco110429, w_eco110430, w_eco110431, w_eco110432, w_eco110433, w_eco110434, w_eco110435, w_eco110436, w_eco110437, w_eco110438, w_eco110439, w_eco110440, w_eco110441, w_eco110442, w_eco110443, w_eco110444, w_eco110445, w_eco110446, w_eco110447, w_eco110448, w_eco110449, w_eco110450, w_eco110451, w_eco110452, w_eco110453, w_eco110454, w_eco110455, w_eco110456, w_eco110457, w_eco110458, w_eco110459, w_eco110460, w_eco110461, w_eco110462, w_eco110463, w_eco110464, w_eco110465, w_eco110466, w_eco110467, w_eco110468, w_eco110469, w_eco110470, w_eco110471, w_eco110472, w_eco110473, w_eco110474, w_eco110475, w_eco110476, w_eco110477, w_eco110478, w_eco110479, w_eco110480, w_eco110481, w_eco110482, w_eco110483, w_eco110484, w_eco110485, w_eco110486, w_eco110487, w_eco110488, w_eco110489, w_eco110490, w_eco110491, w_eco110492, w_eco110493, w_eco110494, w_eco110495, w_eco110496, w_eco110497, w_eco110498, w_eco110499, w_eco110500, w_eco110501, w_eco110502, w_eco110503, w_eco110504, w_eco110505, w_eco110506, w_eco110507, w_eco110508, w_eco110509, w_eco110510, w_eco110511, w_eco110512, w_eco110513, w_eco110514, w_eco110515, w_eco110516, w_eco110517, w_eco110518, w_eco110519, w_eco110520, w_eco110521, w_eco110522, w_eco110523, w_eco110524, w_eco110525, w_eco110526, w_eco110527, w_eco110528, w_eco110529, w_eco110530, w_eco110531, w_eco110532, w_eco110533, w_eco110534, w_eco110535, w_eco110536, w_eco110537, w_eco110538, w_eco110539, w_eco110540, w_eco110541, w_eco110542, w_eco110543, w_eco110544, w_eco110545, w_eco110546, w_eco110547, w_eco110548, w_eco110549, w_eco110550, w_eco110551, w_eco110552, w_eco110553, w_eco110554, w_eco110555, w_eco110556, w_eco110557, w_eco110558, w_eco110559, w_eco110560, w_eco110561, w_eco110562, w_eco110563, w_eco110564, w_eco110565, w_eco110566, w_eco110567, w_eco110568, w_eco110569, w_eco110570, w_eco110571, w_eco110572, w_eco110573, w_eco110574, w_eco110575, w_eco110576, w_eco110577, w_eco110578, w_eco110579, w_eco110580, w_eco110581, w_eco110582, w_eco110583, w_eco110584, w_eco110585, w_eco110586, w_eco110587, w_eco110588, w_eco110589, w_eco110590, w_eco110591, w_eco110592, w_eco110593, w_eco110594, w_eco110595, w_eco110596, w_eco110597, w_eco110598, w_eco110599, w_eco110600, w_eco110601, w_eco110602, w_eco110603, w_eco110604, w_eco110605, w_eco110606, w_eco110607, w_eco110608, w_eco110609, w_eco110610, w_eco110611, w_eco110612, w_eco110613, w_eco110614, w_eco110615, w_eco110616, w_eco110617, w_eco110618, w_eco110619, w_eco110620, w_eco110621, w_eco110622, w_eco110623, w_eco110624, w_eco110625, w_eco110626, w_eco110627, w_eco110628, w_eco110629, w_eco110630, w_eco110631, w_eco110632, w_eco110633, w_eco110634, w_eco110635, w_eco110636, w_eco110637, w_eco110638, w_eco110639, w_eco110640, w_eco110641, w_eco110642, w_eco110643, w_eco110644, w_eco110645, w_eco110646, w_eco110647, w_eco110648, w_eco110649, w_eco110650, w_eco110651, w_eco110652, w_eco110653, w_eco110654, w_eco110655, w_eco110656, w_eco110657, w_eco110658, w_eco110659, w_eco110660, w_eco110661, w_eco110662, w_eco110663, w_eco110664, w_eco110665, w_eco110666, w_eco110667, w_eco110668, w_eco110669, w_eco110670, w_eco110671, w_eco110672, w_eco110673, w_eco110674, w_eco110675, w_eco110676, w_eco110677, w_eco110678, w_eco110679, w_eco110680, w_eco110681, w_eco110682, w_eco110683, w_eco110684, w_eco110685, w_eco110686, w_eco110687, w_eco110688, w_eco110689, w_eco110690, w_eco110691, w_eco110692, w_eco110693, w_eco110694, w_eco110695, w_eco110696, w_eco110697, w_eco110698, w_eco110699, w_eco110700, w_eco110701, w_eco110702, w_eco110703, w_eco110704, w_eco110705, w_eco110706, w_eco110707, w_eco110708, w_eco110709, w_eco110710, w_eco110711, w_eco110712, w_eco110713, w_eco110714, w_eco110715, w_eco110716, w_eco110717, w_eco110718, w_eco110719, w_eco110720, w_eco110721, w_eco110722, w_eco110723, w_eco110724, w_eco110725, w_eco110726, w_eco110727, w_eco110728, w_eco110729, w_eco110730, w_eco110731, w_eco110732, w_eco110733, w_eco110734, w_eco110735, w_eco110736, w_eco110737, w_eco110738, w_eco110739, w_eco110740, w_eco110741, w_eco110742, w_eco110743, w_eco110744, w_eco110745, w_eco110746, w_eco110747, w_eco110748, w_eco110749, w_eco110750, w_eco110751, w_eco110752, w_eco110753, w_eco110754, w_eco110755, w_eco110756, w_eco110757, w_eco110758, w_eco110759, w_eco110760, w_eco110761, w_eco110762, w_eco110763, w_eco110764, w_eco110765, w_eco110766, w_eco110767, w_eco110768, w_eco110769, w_eco110770, w_eco110771, w_eco110772, w_eco110773, w_eco110774, w_eco110775, w_eco110776, w_eco110777, w_eco110778, w_eco110779, w_eco110780, w_eco110781, w_eco110782, w_eco110783, w_eco110784, w_eco110785, w_eco110786, w_eco110787, w_eco110788, w_eco110789, w_eco110790, w_eco110791, w_eco110792, w_eco110793, w_eco110794, w_eco110795, w_eco110796, w_eco110797, w_eco110798, w_eco110799, w_eco110800, w_eco110801, w_eco110802, w_eco110803, w_eco110804, w_eco110805, w_eco110806, w_eco110807, w_eco110808, w_eco110809, w_eco110810, w_eco110811, w_eco110812, w_eco110813, w_eco110814, w_eco110815, w_eco110816, w_eco110817, w_eco110818, w_eco110819, w_eco110820, w_eco110821, w_eco110822, w_eco110823, w_eco110824, w_eco110825, w_eco110826, w_eco110827, w_eco110828, w_eco110829, w_eco110830, w_eco110831, w_eco110832, w_eco110833, w_eco110834, w_eco110835, w_eco110836, w_eco110837, w_eco110838, w_eco110839, w_eco110840, w_eco110841, w_eco110842, w_eco110843, w_eco110844, w_eco110845, w_eco110846, w_eco110847, w_eco110848, w_eco110849, w_eco110850, w_eco110851, w_eco110852, w_eco110853, w_eco110854, w_eco110855, w_eco110856, w_eco110857, w_eco110858, w_eco110859, w_eco110860, w_eco110861, w_eco110862, w_eco110863, w_eco110864, w_eco110865, w_eco110866, w_eco110867, w_eco110868, w_eco110869, w_eco110870, w_eco110871, w_eco110872, w_eco110873, w_eco110874, w_eco110875, w_eco110876, w_eco110877, w_eco110878, w_eco110879, w_eco110880, w_eco110881, w_eco110882, w_eco110883, w_eco110884, w_eco110885, w_eco110886, w_eco110887, w_eco110888, w_eco110889, w_eco110890, w_eco110891, w_eco110892, w_eco110893, w_eco110894, w_eco110895, w_eco110896, w_eco110897, w_eco110898, w_eco110899, w_eco110900, w_eco110901, w_eco110902, w_eco110903, w_eco110904, w_eco110905, w_eco110906, w_eco110907, w_eco110908, w_eco110909, w_eco110910, w_eco110911, w_eco110912, w_eco110913, w_eco110914, w_eco110915, w_eco110916, w_eco110917, w_eco110918, w_eco110919, w_eco110920, w_eco110921, w_eco110922, w_eco110923, w_eco110924, w_eco110925, w_eco110926, w_eco110927, w_eco110928, w_eco110929, w_eco110930, w_eco110931, w_eco110932, w_eco110933, w_eco110934, w_eco110935, w_eco110936, w_eco110937, w_eco110938, w_eco110939, w_eco110940, w_eco110941, w_eco110942, w_eco110943, w_eco110944, w_eco110945, w_eco110946, w_eco110947, w_eco110948, w_eco110949, w_eco110950, w_eco110951, w_eco110952, w_eco110953, w_eco110954, w_eco110955, w_eco110956, w_eco110957, w_eco110958, w_eco110959, w_eco110960, w_eco110961, w_eco110962, w_eco110963, w_eco110964, w_eco110965, w_eco110966, w_eco110967, w_eco110968, w_eco110969, w_eco110970, w_eco110971, w_eco110972, w_eco110973, w_eco110974, w_eco110975, w_eco110976, w_eco110977, w_eco110978, w_eco110979, w_eco110980, w_eco110981, w_eco110982, w_eco110983, w_eco110984, w_eco110985, w_eco110986, w_eco110987, w_eco110988, w_eco110989, w_eco110990, w_eco110991, w_eco110992, w_eco110993, w_eco110994, w_eco110995, w_eco110996, w_eco110997, w_eco110998, w_eco110999, w_eco111000, w_eco111001, w_eco111002, w_eco111003, w_eco111004, w_eco111005, w_eco111006, w_eco111007, w_eco111008, w_eco111009, w_eco111010, w_eco111011, w_eco111012, w_eco111013, w_eco111014, w_eco111015, w_eco111016, w_eco111017, w_eco111018, w_eco111019, w_eco111020, w_eco111021, w_eco111022, w_eco111023, w_eco111024, w_eco111025, w_eco111026, w_eco111027, w_eco111028, w_eco111029, w_eco111030, w_eco111031, w_eco111032, w_eco111033, w_eco111034, w_eco111035, w_eco111036, w_eco111037, w_eco111038, w_eco111039, w_eco111040, w_eco111041, w_eco111042, w_eco111043, w_eco111044, w_eco111045, w_eco111046, w_eco111047, w_eco111048, w_eco111049, w_eco111050, w_eco111051, w_eco111052, w_eco111053, w_eco111054, w_eco111055, w_eco111056, w_eco111057, w_eco111058, w_eco111059, w_eco111060, w_eco111061, w_eco111062, w_eco111063, w_eco111064, w_eco111065, w_eco111066, w_eco111067, w_eco111068, w_eco111069, w_eco111070, w_eco111071, w_eco111072, w_eco111073, w_eco111074, w_eco111075, w_eco111076, w_eco111077, w_eco111078, w_eco111079, w_eco111080, w_eco111081, w_eco111082, w_eco111083, w_eco111084, w_eco111085, w_eco111086, w_eco111087, w_eco111088, w_eco111089, w_eco111090, w_eco111091, w_eco111092, w_eco111093, w_eco111094, w_eco111095, w_eco111096, w_eco111097, w_eco111098, w_eco111099, w_eco111100, w_eco111101, w_eco111102, w_eco111103, w_eco111104, w_eco111105, w_eco111106, w_eco111107, w_eco111108, w_eco111109, w_eco111110, w_eco111111, w_eco111112, w_eco111113, w_eco111114, w_eco111115, w_eco111116, w_eco111117, w_eco111118, w_eco111119, w_eco111120, w_eco111121, w_eco111122, w_eco111123, w_eco111124, w_eco111125, w_eco111126, w_eco111127, w_eco111128, w_eco111129, w_eco111130, w_eco111131, w_eco111132, w_eco111133, w_eco111134, w_eco111135, w_eco111136, w_eco111137, w_eco111138, w_eco111139, w_eco111140, w_eco111141, w_eco111142, w_eco111143, w_eco111144, w_eco111145, w_eco111146, w_eco111147, w_eco111148, w_eco111149, w_eco111150, w_eco111151, w_eco111152, w_eco111153, w_eco111154, w_eco111155, w_eco111156, w_eco111157, w_eco111158, w_eco111159, w_eco111160, w_eco111161, w_eco111162, w_eco111163, w_eco111164, w_eco111165, w_eco111166, w_eco111167, w_eco111168, w_eco111169, w_eco111170, w_eco111171, w_eco111172, w_eco111173, w_eco111174, w_eco111175, w_eco111176, w_eco111177, w_eco111178, w_eco111179, w_eco111180, w_eco111181, w_eco111182, w_eco111183, w_eco111184, w_eco111185, w_eco111186, w_eco111187, w_eco111188, w_eco111189, w_eco111190, w_eco111191, w_eco111192, w_eco111193, w_eco111194, w_eco111195, w_eco111196, w_eco111197, w_eco111198, w_eco111199, w_eco111200, w_eco111201, w_eco111202, w_eco111203, w_eco111204, w_eco111205, w_eco111206, w_eco111207, w_eco111208, w_eco111209, w_eco111210, w_eco111211, w_eco111212, w_eco111213, w_eco111214, w_eco111215, w_eco111216, w_eco111217, w_eco111218, w_eco111219, w_eco111220, w_eco111221, w_eco111222, w_eco111223, w_eco111224, w_eco111225, w_eco111226, w_eco111227, w_eco111228, w_eco111229, w_eco111230, w_eco111231, w_eco111232, w_eco111233, w_eco111234, w_eco111235, w_eco111236, w_eco111237, w_eco111238, w_eco111239, w_eco111240, w_eco111241, w_eco111242, w_eco111243, w_eco111244, w_eco111245, w_eco111246, w_eco111247, w_eco111248, w_eco111249, w_eco111250, w_eco111251, w_eco111252, w_eco111253, w_eco111254, w_eco111255, w_eco111256, w_eco111257, w_eco111258, w_eco111259, w_eco111260, w_eco111261, w_eco111262, w_eco111263, w_eco111264, w_eco111265, w_eco111266, w_eco111267, w_eco111268, w_eco111269, w_eco111270, w_eco111271, w_eco111272, w_eco111273, w_eco111274, w_eco111275, w_eco111276, w_eco111277, w_eco111278, w_eco111279, w_eco111280, w_eco111281, w_eco111282, w_eco111283, w_eco111284, w_eco111285, w_eco111286, w_eco111287, w_eco111288, w_eco111289, w_eco111290, w_eco111291, w_eco111292, w_eco111293, w_eco111294, w_eco111295, w_eco111296, w_eco111297, w_eco111298, w_eco111299, w_eco111300, w_eco111301, w_eco111302, w_eco111303, w_eco111304, w_eco111305, w_eco111306, w_eco111307, w_eco111308, w_eco111309, w_eco111310, w_eco111311, w_eco111312, w_eco111313, w_eco111314, w_eco111315, w_eco111316, w_eco111317, w_eco111318, w_eco111319, w_eco111320, w_eco111321, w_eco111322, w_eco111323, w_eco111324, w_eco111325, w_eco111326, w_eco111327, w_eco111328, w_eco111329, w_eco111330, w_eco111331, w_eco111332, w_eco111333, w_eco111334, w_eco111335, w_eco111336, w_eco111337, w_eco111338, w_eco111339, w_eco111340, w_eco111341, w_eco111342, w_eco111343, w_eco111344, w_eco111345, w_eco111346, w_eco111347, w_eco111348, w_eco111349, w_eco111350, w_eco111351, w_eco111352, w_eco111353, w_eco111354, w_eco111355, w_eco111356, w_eco111357, w_eco111358, w_eco111359, w_eco111360, w_eco111361, w_eco111362, w_eco111363, w_eco111364, w_eco111365, w_eco111366, w_eco111367, w_eco111368, w_eco111369, w_eco111370, w_eco111371, w_eco111372, w_eco111373, w_eco111374, w_eco111375, w_eco111376, w_eco111377, w_eco111378, w_eco111379, w_eco111380, w_eco111381, w_eco111382, w_eco111383, w_eco111384, w_eco111385, w_eco111386, w_eco111387, w_eco111388, w_eco111389, w_eco111390, w_eco111391, w_eco111392, w_eco111393, w_eco111394, w_eco111395, w_eco111396, w_eco111397, w_eco111398, w_eco111399, w_eco111400, w_eco111401, w_eco111402, w_eco111403, w_eco111404, w_eco111405, w_eco111406, w_eco111407, w_eco111408, w_eco111409, w_eco111410, w_eco111411, w_eco111412, w_eco111413, w_eco111414, w_eco111415, w_eco111416, w_eco111417, w_eco111418, w_eco111419, w_eco111420, w_eco111421, w_eco111422, w_eco111423, w_eco111424, w_eco111425, w_eco111426, w_eco111427, w_eco111428, w_eco111429, w_eco111430, w_eco111431, w_eco111432, w_eco111433, w_eco111434, w_eco111435, w_eco111436, w_eco111437, w_eco111438, w_eco111439, w_eco111440, w_eco111441, w_eco111442, w_eco111443, w_eco111444, w_eco111445, w_eco111446, w_eco111447, w_eco111448, w_eco111449, w_eco111450, w_eco111451, w_eco111452, w_eco111453, w_eco111454, w_eco111455, w_eco111456, w_eco111457, w_eco111458, w_eco111459, w_eco111460, w_eco111461, w_eco111462, w_eco111463, w_eco111464, w_eco111465, w_eco111466, w_eco111467, w_eco111468, w_eco111469, w_eco111470, w_eco111471, w_eco111472, w_eco111473, w_eco111474, w_eco111475, w_eco111476, w_eco111477, w_eco111478, w_eco111479, w_eco111480, w_eco111481, w_eco111482, w_eco111483, w_eco111484, w_eco111485, w_eco111486, w_eco111487, w_eco111488, w_eco111489, w_eco111490, w_eco111491, w_eco111492, w_eco111493, w_eco111494, w_eco111495, w_eco111496, w_eco111497, w_eco111498, w_eco111499, w_eco111500, w_eco111501, w_eco111502, w_eco111503, w_eco111504, w_eco111505, w_eco111506, w_eco111507, w_eco111508, w_eco111509, w_eco111510, w_eco111511, w_eco111512, w_eco111513, w_eco111514, w_eco111515, w_eco111516, w_eco111517, w_eco111518, w_eco111519, w_eco111520, w_eco111521, w_eco111522, w_eco111523, w_eco111524, w_eco111525, w_eco111526, w_eco111527, w_eco111528, w_eco111529, w_eco111530, w_eco111531, w_eco111532, w_eco111533, w_eco111534, w_eco111535, w_eco111536, w_eco111537, w_eco111538, w_eco111539, w_eco111540, w_eco111541, w_eco111542, w_eco111543, w_eco111544, w_eco111545, w_eco111546, w_eco111547, w_eco111548, w_eco111549, w_eco111550, w_eco111551, w_eco111552, w_eco111553, w_eco111554, w_eco111555, w_eco111556, w_eco111557, w_eco111558, w_eco111559, w_eco111560, w_eco111561, w_eco111562, w_eco111563, w_eco111564, w_eco111565, w_eco111566, w_eco111567, w_eco111568, w_eco111569, w_eco111570, w_eco111571, w_eco111572, w_eco111573, w_eco111574, w_eco111575, w_eco111576, w_eco111577, w_eco111578, w_eco111579, w_eco111580, w_eco111581, w_eco111582, w_eco111583, w_eco111584, w_eco111585, w_eco111586, w_eco111587, w_eco111588, w_eco111589, w_eco111590, w_eco111591, w_eco111592, w_eco111593, w_eco111594, w_eco111595, w_eco111596, w_eco111597, w_eco111598, w_eco111599, w_eco111600, w_eco111601, w_eco111602, w_eco111603, w_eco111604, w_eco111605, w_eco111606, w_eco111607, w_eco111608, w_eco111609, w_eco111610, w_eco111611, w_eco111612, w_eco111613, w_eco111614, w_eco111615, w_eco111616, w_eco111617, w_eco111618, w_eco111619, w_eco111620, w_eco111621, w_eco111622, w_eco111623, w_eco111624, w_eco111625, w_eco111626, w_eco111627, w_eco111628, w_eco111629, w_eco111630, w_eco111631, w_eco111632, w_eco111633, w_eco111634, w_eco111635, w_eco111636, w_eco111637, w_eco111638, w_eco111639, w_eco111640, w_eco111641, w_eco111642, w_eco111643, w_eco111644, w_eco111645, w_eco111646, w_eco111647, w_eco111648, w_eco111649, w_eco111650, w_eco111651, w_eco111652, w_eco111653, w_eco111654, w_eco111655, w_eco111656, w_eco111657, w_eco111658, w_eco111659, w_eco111660, w_eco111661, w_eco111662, w_eco111663, w_eco111664, w_eco111665, w_eco111666, w_eco111667, w_eco111668, w_eco111669, w_eco111670, w_eco111671, w_eco111672, w_eco111673, w_eco111674, w_eco111675, w_eco111676, w_eco111677, w_eco111678, w_eco111679, w_eco111680, w_eco111681, w_eco111682, w_eco111683, w_eco111684, w_eco111685, w_eco111686, w_eco111687, w_eco111688, w_eco111689, w_eco111690, w_eco111691, w_eco111692, w_eco111693, w_eco111694, w_eco111695, w_eco111696, w_eco111697, w_eco111698, w_eco111699, w_eco111700, w_eco111701, w_eco111702, w_eco111703, w_eco111704, w_eco111705, w_eco111706, w_eco111707, w_eco111708, w_eco111709, w_eco111710, w_eco111711, w_eco111712, w_eco111713, w_eco111714, w_eco111715, w_eco111716, w_eco111717, w_eco111718, w_eco111719, w_eco111720, w_eco111721, w_eco111722, w_eco111723, w_eco111724, w_eco111725, w_eco111726, w_eco111727, w_eco111728, w_eco111729, w_eco111730, w_eco111731, w_eco111732, w_eco111733, w_eco111734, w_eco111735, w_eco111736, w_eco111737, w_eco111738, w_eco111739, w_eco111740, w_eco111741, w_eco111742, w_eco111743, w_eco111744, w_eco111745, w_eco111746, w_eco111747, w_eco111748, w_eco111749, w_eco111750, w_eco111751, w_eco111752, w_eco111753, w_eco111754, w_eco111755, w_eco111756, w_eco111757, w_eco111758, w_eco111759, w_eco111760, w_eco111761, w_eco111762, w_eco111763, w_eco111764, w_eco111765, w_eco111766, w_eco111767, w_eco111768, w_eco111769, w_eco111770, w_eco111771, w_eco111772, w_eco111773, w_eco111774, w_eco111775, w_eco111776, w_eco111777, w_eco111778, w_eco111779, w_eco111780, w_eco111781, w_eco111782, w_eco111783, w_eco111784, w_eco111785, w_eco111786, w_eco111787, w_eco111788, w_eco111789, w_eco111790, w_eco111791, w_eco111792, w_eco111793, w_eco111794, w_eco111795, w_eco111796, w_eco111797, w_eco111798, w_eco111799, w_eco111800, w_eco111801, w_eco111802, w_eco111803, w_eco111804, w_eco111805, w_eco111806, w_eco111807, w_eco111808, w_eco111809, w_eco111810, w_eco111811, w_eco111812, w_eco111813, w_eco111814, w_eco111815, w_eco111816, w_eco111817, w_eco111818, w_eco111819, w_eco111820, w_eco111821, w_eco111822, w_eco111823, w_eco111824, w_eco111825, w_eco111826, w_eco111827, w_eco111828, w_eco111829, w_eco111830, w_eco111831, w_eco111832, w_eco111833, w_eco111834, w_eco111835, w_eco111836, w_eco111837, w_eco111838, w_eco111839, w_eco111840, w_eco111841, w_eco111842, w_eco111843, w_eco111844, w_eco111845, w_eco111846, w_eco111847, w_eco111848, w_eco111849, w_eco111850, w_eco111851, w_eco111852, w_eco111853, w_eco111854, w_eco111855, w_eco111856, w_eco111857, w_eco111858, w_eco111859, w_eco111860, w_eco111861, w_eco111862, w_eco111863, w_eco111864, w_eco111865, w_eco111866, w_eco111867, w_eco111868, w_eco111869, w_eco111870, w_eco111871, w_eco111872, w_eco111873, w_eco111874, w_eco111875, w_eco111876, w_eco111877, w_eco111878, w_eco111879, w_eco111880, w_eco111881, w_eco111882, w_eco111883, w_eco111884, w_eco111885, w_eco111886, w_eco111887, w_eco111888, w_eco111889, w_eco111890, w_eco111891, w_eco111892, w_eco111893, w_eco111894, w_eco111895, w_eco111896, w_eco111897, w_eco111898, w_eco111899, w_eco111900, w_eco111901, w_eco111902, w_eco111903, w_eco111904, w_eco111905, w_eco111906, w_eco111907, w_eco111908, w_eco111909, w_eco111910, w_eco111911, w_eco111912, w_eco111913, w_eco111914, w_eco111915, w_eco111916, w_eco111917, w_eco111918, w_eco111919, w_eco111920, w_eco111921, w_eco111922, w_eco111923, w_eco111924, w_eco111925, w_eco111926, w_eco111927, w_eco111928, w_eco111929, w_eco111930, w_eco111931, w_eco111932, w_eco111933, w_eco111934, w_eco111935, w_eco111936, w_eco111937, w_eco111938, w_eco111939, w_eco111940, w_eco111941, w_eco111942, w_eco111943, w_eco111944, w_eco111945, w_eco111946, w_eco111947, w_eco111948, w_eco111949, w_eco111950, w_eco111951, w_eco111952, w_eco111953, w_eco111954, w_eco111955, w_eco111956, w_eco111957, w_eco111958, w_eco111959, w_eco111960, w_eco111961, w_eco111962, w_eco111963, w_eco111964, w_eco111965, w_eco111966, w_eco111967, w_eco111968, w_eco111969, w_eco111970, w_eco111971, w_eco111972, w_eco111973, w_eco111974, w_eco111975, w_eco111976, w_eco111977, w_eco111978, w_eco111979, w_eco111980, w_eco111981, w_eco111982, w_eco111983, w_eco111984, w_eco111985, w_eco111986, w_eco111987, w_eco111988, w_eco111989, w_eco111990, w_eco111991, w_eco111992, w_eco111993, w_eco111994, w_eco111995, w_eco111996, w_eco111997, w_eco111998, w_eco111999, w_eco112000, w_eco112001, w_eco112002, w_eco112003, w_eco112004, w_eco112005, w_eco112006, w_eco112007, w_eco112008, w_eco112009, w_eco112010, w_eco112011, w_eco112012, w_eco112013, w_eco112014, w_eco112015, w_eco112016, w_eco112017, w_eco112018, w_eco112019, w_eco112020, w_eco112021, w_eco112022, w_eco112023, w_eco112024, w_eco112025, w_eco112026, w_eco112027, w_eco112028, w_eco112029, w_eco112030, w_eco112031, w_eco112032, w_eco112033, w_eco112034, w_eco112035, w_eco112036, w_eco112037, w_eco112038, w_eco112039, w_eco112040, w_eco112041, w_eco112042, w_eco112043, w_eco112044, w_eco112045, w_eco112046, w_eco112047, w_eco112048, w_eco112049, w_eco112050, w_eco112051, w_eco112052, w_eco112053, w_eco112054, w_eco112055, w_eco112056, w_eco112057, w_eco112058, w_eco112059, w_eco112060, w_eco112061, w_eco112062, w_eco112063, w_eco112064, w_eco112065, w_eco112066, w_eco112067, w_eco112068, w_eco112069, w_eco112070, w_eco112071, w_eco112072, w_eco112073, w_eco112074, w_eco112075, w_eco112076, w_eco112077, w_eco112078, w_eco112079, w_eco112080, w_eco112081, w_eco112082, w_eco112083, w_eco112084, w_eco112085, w_eco112086, w_eco112087, w_eco112088, w_eco112089, w_eco112090, w_eco112091, w_eco112092, w_eco112093, w_eco112094, w_eco112095, w_eco112096, w_eco112097, w_eco112098, w_eco112099, w_eco112100, w_eco112101, w_eco112102, w_eco112103, w_eco112104, w_eco112105, w_eco112106, w_eco112107, w_eco112108, w_eco112109, w_eco112110, w_eco112111, w_eco112112, w_eco112113, w_eco112114, w_eco112115, w_eco112116, w_eco112117, w_eco112118, w_eco112119, w_eco112120, w_eco112121, w_eco112122, w_eco112123, w_eco112124, w_eco112125, w_eco112126, w_eco112127, w_eco112128, w_eco112129, w_eco112130, w_eco112131, w_eco112132, w_eco112133, w_eco112134, w_eco112135, w_eco112136, w_eco112137, w_eco112138, w_eco112139, w_eco112140, w_eco112141, w_eco112142, w_eco112143, w_eco112144, w_eco112145, w_eco112146, w_eco112147, w_eco112148, w_eco112149, w_eco112150, w_eco112151, w_eco112152, w_eco112153, w_eco112154, w_eco112155, w_eco112156, w_eco112157, w_eco112158, w_eco112159, w_eco112160, w_eco112161, w_eco112162, w_eco112163, w_eco112164, w_eco112165, w_eco112166, w_eco112167, w_eco112168, w_eco112169, w_eco112170, w_eco112171, w_eco112172, w_eco112173, w_eco112174, w_eco112175, w_eco112176, w_eco112177, w_eco112178, w_eco112179, w_eco112180, w_eco112181, w_eco112182, w_eco112183, w_eco112184, w_eco112185, w_eco112186, w_eco112187, w_eco112188, w_eco112189, w_eco112190, w_eco112191, w_eco112192, w_eco112193, w_eco112194, w_eco112195, w_eco112196, w_eco112197, w_eco112198, w_eco112199, w_eco112200, w_eco112201, w_eco112202, w_eco112203, w_eco112204, w_eco112205, w_eco112206, w_eco112207, w_eco112208, w_eco112209, w_eco112210, w_eco112211, w_eco112212, w_eco112213, w_eco112214, w_eco112215, w_eco112216, w_eco112217, w_eco112218, w_eco112219, w_eco112220, w_eco112221, w_eco112222, w_eco112223, w_eco112224, w_eco112225, w_eco112226, w_eco112227, w_eco112228, w_eco112229, w_eco112230, w_eco112231, w_eco112232, w_eco112233, w_eco112234, w_eco112235, w_eco112236, w_eco112237, w_eco112238, w_eco112239, w_eco112240, w_eco112241, w_eco112242, w_eco112243, w_eco112244, w_eco112245, w_eco112246, w_eco112247, w_eco112248, w_eco112249, w_eco112250, w_eco112251, w_eco112252, w_eco112253, w_eco112254, w_eco112255, w_eco112256, w_eco112257, w_eco112258, w_eco112259, w_eco112260, w_eco112261, w_eco112262, w_eco112263, w_eco112264, w_eco112265, w_eco112266, w_eco112267, w_eco112268, w_eco112269, w_eco112270, w_eco112271, w_eco112272, w_eco112273, w_eco112274, w_eco112275, w_eco112276, w_eco112277, w_eco112278, w_eco112279, w_eco112280, w_eco112281, w_eco112282, w_eco112283, w_eco112284, w_eco112285, w_eco112286, w_eco112287, w_eco112288, w_eco112289, w_eco112290, w_eco112291, w_eco112292, w_eco112293, w_eco112294, w_eco112295, w_eco112296, w_eco112297, w_eco112298, w_eco112299, w_eco112300, w_eco112301, w_eco112302, w_eco112303, w_eco112304, w_eco112305, w_eco112306, w_eco112307, w_eco112308, w_eco112309, w_eco112310, w_eco112311, w_eco112312, w_eco112313, w_eco112314, w_eco112315, w_eco112316, w_eco112317, w_eco112318, w_eco112319, w_eco112320, w_eco112321, w_eco112322, w_eco112323, w_eco112324, w_eco112325, w_eco112326, w_eco112327, w_eco112328, w_eco112329, w_eco112330, w_eco112331, w_eco112332, w_eco112333, w_eco112334, w_eco112335, w_eco112336, w_eco112337, w_eco112338, w_eco112339, w_eco112340, w_eco112341, w_eco112342, w_eco112343, w_eco112344, w_eco112345, w_eco112346, w_eco112347, w_eco112348, w_eco112349, w_eco112350, w_eco112351, w_eco112352, w_eco112353, w_eco112354, w_eco112355, w_eco112356, w_eco112357, w_eco112358, w_eco112359, w_eco112360, w_eco112361, w_eco112362, w_eco112363, w_eco112364, w_eco112365, w_eco112366, w_eco112367, w_eco112368, w_eco112369, w_eco112370, w_eco112371, w_eco112372, w_eco112373, w_eco112374, w_eco112375, w_eco112376, w_eco112377, w_eco112378, w_eco112379, w_eco112380, w_eco112381, w_eco112382, w_eco112383, w_eco112384, w_eco112385, w_eco112386, w_eco112387, w_eco112388, w_eco112389, w_eco112390, w_eco112391, w_eco112392, w_eco112393, w_eco112394, w_eco112395, w_eco112396, w_eco112397, w_eco112398, w_eco112399, w_eco112400, w_eco112401, w_eco112402, w_eco112403, w_eco112404, w_eco112405, w_eco112406, w_eco112407, w_eco112408, w_eco112409, w_eco112410, w_eco112411, w_eco112412, w_eco112413, w_eco112414, w_eco112415, w_eco112416, w_eco112417, w_eco112418, w_eco112419, w_eco112420, w_eco112421, w_eco112422, w_eco112423, w_eco112424, w_eco112425, w_eco112426, w_eco112427, w_eco112428, w_eco112429, w_eco112430, w_eco112431, w_eco112432, w_eco112433, w_eco112434, w_eco112435, w_eco112436, w_eco112437, w_eco112438, w_eco112439, w_eco112440, w_eco112441, w_eco112442, w_eco112443, w_eco112444, w_eco112445, w_eco112446, w_eco112447, w_eco112448, w_eco112449, w_eco112450, w_eco112451, w_eco112452, w_eco112453, w_eco112454, w_eco112455, w_eco112456, w_eco112457, w_eco112458, w_eco112459, w_eco112460, w_eco112461, w_eco112462, w_eco112463, w_eco112464, w_eco112465, w_eco112466, w_eco112467, w_eco112468, w_eco112469, w_eco112470, w_eco112471, w_eco112472, w_eco112473, w_eco112474, w_eco112475, w_eco112476, w_eco112477, w_eco112478, w_eco112479, w_eco112480, w_eco112481, w_eco112482, w_eco112483, w_eco112484, w_eco112485, w_eco112486, w_eco112487, w_eco112488, w_eco112489, w_eco112490, w_eco112491, w_eco112492, w_eco112493, w_eco112494, w_eco112495, w_eco112496, w_eco112497, w_eco112498, w_eco112499, w_eco112500, w_eco112501, w_eco112502, w_eco112503, w_eco112504, w_eco112505, w_eco112506, w_eco112507, w_eco112508, w_eco112509, w_eco112510, w_eco112511, w_eco112512, w_eco112513, w_eco112514, w_eco112515, w_eco112516, w_eco112517, w_eco112518, w_eco112519, w_eco112520, w_eco112521, w_eco112522, w_eco112523, w_eco112524, w_eco112525, w_eco112526, w_eco112527, w_eco112528, w_eco112529, w_eco112530, w_eco112531, w_eco112532, w_eco112533, w_eco112534, w_eco112535, w_eco112536, w_eco112537, w_eco112538, w_eco112539, w_eco112540, w_eco112541, w_eco112542, w_eco112543, w_eco112544, w_eco112545, w_eco112546, w_eco112547, w_eco112548, w_eco112549, w_eco112550, w_eco112551, w_eco112552, w_eco112553, w_eco112554, w_eco112555, w_eco112556, w_eco112557, w_eco112558, w_eco112559, w_eco112560, w_eco112561, w_eco112562, w_eco112563, w_eco112564, w_eco112565, w_eco112566, w_eco112567, w_eco112568, w_eco112569, w_eco112570, w_eco112571, w_eco112572, w_eco112573, w_eco112574, w_eco112575, w_eco112576, w_eco112577, w_eco112578, w_eco112579, w_eco112580, w_eco112581, w_eco112582, w_eco112583, w_eco112584, w_eco112585, w_eco112586, w_eco112587, w_eco112588, w_eco112589, w_eco112590, w_eco112591, w_eco112592, w_eco112593, w_eco112594, w_eco112595, w_eco112596, w_eco112597, w_eco112598, w_eco112599, w_eco112600, w_eco112601, w_eco112602, w_eco112603, w_eco112604, w_eco112605, w_eco112606, w_eco112607, w_eco112608, w_eco112609, w_eco112610, w_eco112611, w_eco112612, w_eco112613, w_eco112614, w_eco112615, w_eco112616, w_eco112617, w_eco112618, w_eco112619, w_eco112620, w_eco112621, w_eco112622, w_eco112623, w_eco112624, w_eco112625, w_eco112626, w_eco112627, w_eco112628, w_eco112629, w_eco112630, w_eco112631, w_eco112632, w_eco112633, w_eco112634, w_eco112635, w_eco112636, w_eco112637, w_eco112638, w_eco112639, w_eco112640, w_eco112641, w_eco112642, w_eco112643, w_eco112644, w_eco112645, w_eco112646, w_eco112647, w_eco112648, w_eco112649, w_eco112650, w_eco112651, w_eco112652, w_eco112653, w_eco112654, w_eco112655, w_eco112656, w_eco112657, w_eco112658, w_eco112659, w_eco112660, w_eco112661, w_eco112662, w_eco112663, w_eco112664, w_eco112665, w_eco112666, w_eco112667, w_eco112668, w_eco112669, w_eco112670, w_eco112671, w_eco112672, w_eco112673, w_eco112674, w_eco112675, w_eco112676, w_eco112677, w_eco112678, w_eco112679, w_eco112680, w_eco112681, w_eco112682, w_eco112683, w_eco112684, w_eco112685, w_eco112686, w_eco112687, w_eco112688, w_eco112689, w_eco112690, w_eco112691, w_eco112692, w_eco112693, w_eco112694, w_eco112695, w_eco112696, w_eco112697, w_eco112698, w_eco112699, w_eco112700, w_eco112701, w_eco112702, w_eco112703, w_eco112704, w_eco112705, w_eco112706, w_eco112707, w_eco112708, w_eco112709, w_eco112710, w_eco112711, w_eco112712, w_eco112713, w_eco112714, w_eco112715, w_eco112716, w_eco112717, w_eco112718, w_eco112719, w_eco112720, w_eco112721, w_eco112722, w_eco112723, w_eco112724, w_eco112725, w_eco112726, w_eco112727, w_eco112728, w_eco112729, w_eco112730, w_eco112731, w_eco112732, w_eco112733, w_eco112734, w_eco112735, w_eco112736, w_eco112737, w_eco112738, w_eco112739, w_eco112740, w_eco112741, w_eco112742, w_eco112743, w_eco112744, w_eco112745, w_eco112746, w_eco112747, w_eco112748, w_eco112749, w_eco112750, w_eco112751, w_eco112752, w_eco112753, w_eco112754, w_eco112755, w_eco112756, w_eco112757, w_eco112758, w_eco112759, w_eco112760, w_eco112761, w_eco112762, w_eco112763, w_eco112764, w_eco112765, w_eco112766, w_eco112767, w_eco112768, w_eco112769, w_eco112770, w_eco112771, w_eco112772, w_eco112773, w_eco112774, w_eco112775, w_eco112776, w_eco112777, w_eco112778, w_eco112779, w_eco112780, w_eco112781, w_eco112782, w_eco112783, w_eco112784, w_eco112785, w_eco112786, w_eco112787, w_eco112788, w_eco112789, w_eco112790, w_eco112791, w_eco112792, w_eco112793, w_eco112794, w_eco112795, w_eco112796, w_eco112797, w_eco112798, w_eco112799, w_eco112800, w_eco112801, w_eco112802, w_eco112803, w_eco112804, w_eco112805, w_eco112806, w_eco112807, w_eco112808, w_eco112809, w_eco112810, w_eco112811, w_eco112812, w_eco112813, w_eco112814, w_eco112815, w_eco112816, w_eco112817, w_eco112818, w_eco112819, w_eco112820, w_eco112821, w_eco112822, w_eco112823, w_eco112824, w_eco112825, w_eco112826, w_eco112827, w_eco112828, w_eco112829, w_eco112830, w_eco112831, w_eco112832, w_eco112833, w_eco112834, w_eco112835, w_eco112836, w_eco112837, w_eco112838, w_eco112839, w_eco112840, w_eco112841, w_eco112842, w_eco112843, w_eco112844, w_eco112845, w_eco112846, w_eco112847, w_eco112848, w_eco112849, w_eco112850, w_eco112851, w_eco112852, w_eco112853, w_eco112854, w_eco112855, w_eco112856, w_eco112857, w_eco112858, w_eco112859, w_eco112860, w_eco112861, w_eco112862, w_eco112863, w_eco112864, w_eco112865, w_eco112866, w_eco112867, w_eco112868, w_eco112869, w_eco112870, w_eco112871, w_eco112872, w_eco112873, w_eco112874, w_eco112875, w_eco112876, w_eco112877, w_eco112878, w_eco112879, w_eco112880, w_eco112881, w_eco112882, w_eco112883, w_eco112884, w_eco112885, w_eco112886, w_eco112887, w_eco112888, w_eco112889, w_eco112890, w_eco112891, w_eco112892, w_eco112893, w_eco112894, w_eco112895, w_eco112896, w_eco112897, w_eco112898, w_eco112899, w_eco112900, w_eco112901, w_eco112902, w_eco112903, w_eco112904, w_eco112905, w_eco112906, w_eco112907, w_eco112908, w_eco112909, w_eco112910, w_eco112911, w_eco112912, w_eco112913, w_eco112914, w_eco112915, w_eco112916, w_eco112917, w_eco112918, w_eco112919, w_eco112920, w_eco112921, w_eco112922, w_eco112923, w_eco112924, w_eco112925, w_eco112926, w_eco112927, w_eco112928, w_eco112929, w_eco112930, w_eco112931, w_eco112932, w_eco112933, w_eco112934, w_eco112935, w_eco112936, w_eco112937, w_eco112938, w_eco112939, w_eco112940, w_eco112941, w_eco112942, w_eco112943, w_eco112944, w_eco112945, w_eco112946, w_eco112947, w_eco112948, w_eco112949, w_eco112950, w_eco112951, w_eco112952, w_eco112953, w_eco112954, w_eco112955, w_eco112956, w_eco112957, w_eco112958, w_eco112959, w_eco112960, w_eco112961, w_eco112962, w_eco112963, w_eco112964, w_eco112965, w_eco112966, w_eco112967, w_eco112968, w_eco112969, w_eco112970, w_eco112971, w_eco112972, w_eco112973, w_eco112974, w_eco112975, w_eco112976, w_eco112977, w_eco112978, w_eco112979, w_eco112980, w_eco112981, w_eco112982, w_eco112983, w_eco112984, w_eco112985, w_eco112986, w_eco112987, w_eco112988, w_eco112989, w_eco112990, w_eco112991, w_eco112992, w_eco112993, w_eco112994, w_eco112995, w_eco112996, w_eco112997, w_eco112998, w_eco112999, w_eco113000, w_eco113001, w_eco113002, w_eco113003, w_eco113004, w_eco113005, w_eco113006, w_eco113007, w_eco113008, w_eco113009, w_eco113010, w_eco113011, w_eco113012, w_eco113013, w_eco113014, w_eco113015, w_eco113016, w_eco113017, w_eco113018, w_eco113019, w_eco113020, w_eco113021, w_eco113022, w_eco113023, w_eco113024, w_eco113025, w_eco113026, w_eco113027, w_eco113028, w_eco113029, w_eco113030, w_eco113031, w_eco113032, w_eco113033, w_eco113034, w_eco113035, w_eco113036, w_eco113037, w_eco113038, w_eco113039, w_eco113040, w_eco113041, w_eco113042, w_eco113043, w_eco113044, w_eco113045, w_eco113046, w_eco113047, w_eco113048, w_eco113049, w_eco113050, w_eco113051, w_eco113052, w_eco113053, w_eco113054, w_eco113055, w_eco113056, w_eco113057, w_eco113058, w_eco113059, w_eco113060, w_eco113061, w_eco113062, w_eco113063, w_eco113064, w_eco113065, w_eco113066, w_eco113067, w_eco113068, w_eco113069, w_eco113070, w_eco113071, w_eco113072, w_eco113073, w_eco113074, w_eco113075, w_eco113076, w_eco113077, w_eco113078, w_eco113079, w_eco113080, w_eco113081, w_eco113082, w_eco113083, w_eco113084, w_eco113085, w_eco113086, w_eco113087, w_eco113088, w_eco113089, w_eco113090, w_eco113091, w_eco113092, w_eco113093, w_eco113094, w_eco113095, w_eco113096, w_eco113097, w_eco113098, w_eco113099, w_eco113100, w_eco113101, w_eco113102, w_eco113103, w_eco113104, w_eco113105, w_eco113106, w_eco113107, w_eco113108, w_eco113109, w_eco113110, w_eco113111, w_eco113112, w_eco113113, w_eco113114, w_eco113115, w_eco113116, w_eco113117, w_eco113118, w_eco113119, w_eco113120, w_eco113121, w_eco113122, w_eco113123, w_eco113124, w_eco113125, w_eco113126, w_eco113127, w_eco113128, w_eco113129, w_eco113130, w_eco113131, w_eco113132, w_eco113133, w_eco113134, w_eco113135, w_eco113136, w_eco113137, w_eco113138, w_eco113139, w_eco113140, w_eco113141, w_eco113142, w_eco113143, w_eco113144, w_eco113145, w_eco113146, w_eco113147, w_eco113148, w_eco113149, w_eco113150, w_eco113151, w_eco113152, w_eco113153, w_eco113154, w_eco113155, w_eco113156, w_eco113157, w_eco113158, w_eco113159, w_eco113160, w_eco113161, w_eco113162, w_eco113163, w_eco113164, w_eco113165, w_eco113166, w_eco113167, w_eco113168, w_eco113169, w_eco113170, w_eco113171, w_eco113172, w_eco113173, w_eco113174, w_eco113175, w_eco113176, w_eco113177, w_eco113178, w_eco113179, w_eco113180, w_eco113181, w_eco113182, w_eco113183, w_eco113184, w_eco113185, w_eco113186, w_eco113187, w_eco113188, w_eco113189, w_eco113190, w_eco113191, w_eco113192, w_eco113193, w_eco113194, w_eco113195, w_eco113196, w_eco113197, w_eco113198, w_eco113199, w_eco113200, w_eco113201, w_eco113202, w_eco113203, w_eco113204, w_eco113205, w_eco113206, w_eco113207, w_eco113208, w_eco113209, w_eco113210, w_eco113211, w_eco113212, w_eco113213, w_eco113214, w_eco113215, w_eco113216, w_eco113217, w_eco113218, w_eco113219, w_eco113220, w_eco113221, w_eco113222, w_eco113223, w_eco113224, w_eco113225, w_eco113226, w_eco113227, w_eco113228, w_eco113229, w_eco113230, w_eco113231, w_eco113232, w_eco113233, w_eco113234, w_eco113235, w_eco113236, w_eco113237, w_eco113238, w_eco113239, w_eco113240, w_eco113241, w_eco113242, w_eco113243, w_eco113244, w_eco113245, w_eco113246, w_eco113247, w_eco113248, w_eco113249, w_eco113250, w_eco113251, w_eco113252, w_eco113253, w_eco113254, w_eco113255, w_eco113256, w_eco113257, w_eco113258, w_eco113259, w_eco113260, w_eco113261, w_eco113262, w_eco113263, w_eco113264, w_eco113265, w_eco113266, w_eco113267, w_eco113268, w_eco113269, w_eco113270, w_eco113271, w_eco113272, w_eco113273, w_eco113274, w_eco113275, w_eco113276, w_eco113277, w_eco113278, w_eco113279, w_eco113280, w_eco113281, w_eco113282, w_eco113283, w_eco113284, w_eco113285, w_eco113286, w_eco113287, w_eco113288, w_eco113289, w_eco113290, w_eco113291, w_eco113292, w_eco113293, w_eco113294, w_eco113295, w_eco113296, w_eco113297, w_eco113298, w_eco113299, w_eco113300, w_eco113301, w_eco113302, w_eco113303, w_eco113304, w_eco113305, w_eco113306, w_eco113307, w_eco113308, w_eco113309, w_eco113310, w_eco113311, w_eco113312, w_eco113313, w_eco113314, w_eco113315, w_eco113316, w_eco113317, w_eco113318, w_eco113319, w_eco113320, w_eco113321, w_eco113322, w_eco113323, w_eco113324, w_eco113325, w_eco113326, w_eco113327, w_eco113328, w_eco113329, w_eco113330, w_eco113331, w_eco113332, w_eco113333, w_eco113334, w_eco113335, w_eco113336, w_eco113337, w_eco113338, w_eco113339, w_eco113340, w_eco113341, w_eco113342, w_eco113343, w_eco113344, w_eco113345, w_eco113346, w_eco113347, w_eco113348, w_eco113349, w_eco113350, w_eco113351, w_eco113352, w_eco113353, w_eco113354, w_eco113355, w_eco113356, w_eco113357, w_eco113358, w_eco113359, w_eco113360, w_eco113361, w_eco113362, w_eco113363, w_eco113364, w_eco113365, w_eco113366, w_eco113367, w_eco113368, w_eco113369, w_eco113370, w_eco113371, w_eco113372, w_eco113373, w_eco113374, w_eco113375, w_eco113376, w_eco113377, w_eco113378, w_eco113379, w_eco113380, w_eco113381, w_eco113382, w_eco113383, w_eco113384, w_eco113385, w_eco113386, w_eco113387, w_eco113388, w_eco113389, w_eco113390, w_eco113391, w_eco113392, w_eco113393, w_eco113394, w_eco113395, w_eco113396, w_eco113397, w_eco113398, w_eco113399, w_eco113400, w_eco113401, w_eco113402, w_eco113403, w_eco113404, w_eco113405, w_eco113406, w_eco113407, w_eco113408, w_eco113409, w_eco113410, w_eco113411, w_eco113412, w_eco113413, w_eco113414, w_eco113415, w_eco113416, w_eco113417, w_eco113418, w_eco113419, w_eco113420, w_eco113421, w_eco113422, w_eco113423, w_eco113424, w_eco113425, w_eco113426, w_eco113427, w_eco113428, w_eco113429, w_eco113430, w_eco113431, w_eco113432, w_eco113433, w_eco113434, w_eco113435, w_eco113436, w_eco113437, w_eco113438, w_eco113439, w_eco113440, w_eco113441, w_eco113442, w_eco113443, w_eco113444, w_eco113445, w_eco113446, w_eco113447, w_eco113448, w_eco113449, w_eco113450, w_eco113451, w_eco113452, w_eco113453, w_eco113454, w_eco113455, w_eco113456, w_eco113457, w_eco113458, w_eco113459, w_eco113460, w_eco113461, w_eco113462, w_eco113463, w_eco113464, w_eco113465, w_eco113466, w_eco113467, w_eco113468, w_eco113469, w_eco113470, w_eco113471, w_eco113472, w_eco113473, w_eco113474, w_eco113475, w_eco113476, w_eco113477, w_eco113478, w_eco113479, w_eco113480, w_eco113481, w_eco113482, w_eco113483, w_eco113484, w_eco113485, w_eco113486, w_eco113487, w_eco113488, w_eco113489, w_eco113490, w_eco113491, w_eco113492, w_eco113493, w_eco113494, w_eco113495, w_eco113496, w_eco113497, w_eco113498, w_eco113499, w_eco113500, w_eco113501, w_eco113502, w_eco113503, w_eco113504, w_eco113505, w_eco113506, w_eco113507, w_eco113508, w_eco113509, w_eco113510, w_eco113511, w_eco113512, w_eco113513, w_eco113514, w_eco113515, w_eco113516, w_eco113517, w_eco113518, w_eco113519, w_eco113520, w_eco113521, w_eco113522, w_eco113523, w_eco113524, w_eco113525, w_eco113526, w_eco113527, w_eco113528, w_eco113529, w_eco113530, w_eco113531, w_eco113532, w_eco113533, w_eco113534, w_eco113535, w_eco113536, w_eco113537, w_eco113538, w_eco113539, w_eco113540, w_eco113541, w_eco113542, w_eco113543, w_eco113544, w_eco113545, w_eco113546, w_eco113547, w_eco113548, w_eco113549, w_eco113550, w_eco113551, w_eco113552, w_eco113553, w_eco113554, w_eco113555, w_eco113556, w_eco113557, w_eco113558, w_eco113559, w_eco113560, w_eco113561, w_eco113562, w_eco113563, w_eco113564, w_eco113565, w_eco113566, w_eco113567, w_eco113568, w_eco113569, w_eco113570, w_eco113571, w_eco113572, w_eco113573, w_eco113574, w_eco113575, w_eco113576, w_eco113577, w_eco113578, w_eco113579, w_eco113580, w_eco113581, w_eco113582, w_eco113583, w_eco113584, w_eco113585, w_eco113586, w_eco113587, w_eco113588, w_eco113589, w_eco113590, w_eco113591, w_eco113592, w_eco113593, w_eco113594, w_eco113595, w_eco113596, w_eco113597, w_eco113598, w_eco113599, w_eco113600, w_eco113601, w_eco113602, w_eco113603, w_eco113604, w_eco113605, w_eco113606, w_eco113607, w_eco113608, w_eco113609, w_eco113610, w_eco113611, w_eco113612, w_eco113613, w_eco113614, w_eco113615, w_eco113616, w_eco113617, w_eco113618, w_eco113619, w_eco113620, w_eco113621, w_eco113622, w_eco113623, w_eco113624, w_eco113625, w_eco113626, w_eco113627, w_eco113628, w_eco113629, w_eco113630, w_eco113631, w_eco113632, w_eco113633, w_eco113634, w_eco113635, w_eco113636, w_eco113637, w_eco113638, w_eco113639, w_eco113640, w_eco113641, w_eco113642, w_eco113643, w_eco113644, w_eco113645, w_eco113646, w_eco113647, w_eco113648, w_eco113649, w_eco113650, w_eco113651, w_eco113652, w_eco113653, w_eco113654, w_eco113655, w_eco113656, w_eco113657, w_eco113658, w_eco113659, w_eco113660, w_eco113661, w_eco113662, w_eco113663, w_eco113664, w_eco113665, w_eco113666, w_eco113667, w_eco113668, w_eco113669, w_eco113670, w_eco113671, w_eco113672, w_eco113673, w_eco113674, w_eco113675, w_eco113676, w_eco113677, w_eco113678, w_eco113679, w_eco113680, w_eco113681, w_eco113682, w_eco113683, w_eco113684, w_eco113685, w_eco113686, w_eco113687, w_eco113688, w_eco113689, w_eco113690, w_eco113691, w_eco113692, w_eco113693, w_eco113694, w_eco113695, w_eco113696, w_eco113697, w_eco113698, w_eco113699, w_eco113700, w_eco113701, w_eco113702, w_eco113703, w_eco113704, w_eco113705, w_eco113706, w_eco113707, w_eco113708, w_eco113709, w_eco113710, w_eco113711, w_eco113712, w_eco113713, w_eco113714, w_eco113715, w_eco113716, w_eco113717, w_eco113718, w_eco113719, w_eco113720, w_eco113721, w_eco113722, w_eco113723, w_eco113724, w_eco113725, w_eco113726, w_eco113727, w_eco113728, w_eco113729, w_eco113730, w_eco113731, w_eco113732, w_eco113733, w_eco113734, w_eco113735, w_eco113736, w_eco113737, w_eco113738, w_eco113739, w_eco113740, w_eco113741, w_eco113742, w_eco113743, w_eco113744, w_eco113745, w_eco113746, w_eco113747, w_eco113748, w_eco113749, w_eco113750, w_eco113751, w_eco113752, w_eco113753, w_eco113754, w_eco113755, w_eco113756, w_eco113757, w_eco113758, w_eco113759, w_eco113760, w_eco113761, w_eco113762, w_eco113763, w_eco113764, w_eco113765, w_eco113766, w_eco113767, w_eco113768, w_eco113769, w_eco113770, w_eco113771, w_eco113772, w_eco113773, w_eco113774, w_eco113775, w_eco113776, w_eco113777, w_eco113778, w_eco113779, w_eco113780, w_eco113781, w_eco113782, w_eco113783, w_eco113784, w_eco113785, w_eco113786, w_eco113787, w_eco113788, w_eco113789, w_eco113790, w_eco113791, w_eco113792, w_eco113793, w_eco113794, w_eco113795, w_eco113796, w_eco113797, w_eco113798, w_eco113799, w_eco113800, w_eco113801, w_eco113802, w_eco113803, w_eco113804, w_eco113805, w_eco113806, w_eco113807, w_eco113808, w_eco113809, w_eco113810, w_eco113811, w_eco113812, w_eco113813, w_eco113814, w_eco113815, w_eco113816, w_eco113817, w_eco113818, w_eco113819, w_eco113820, w_eco113821, w_eco113822, w_eco113823, w_eco113824, w_eco113825, w_eco113826, w_eco113827, w_eco113828, w_eco113829, w_eco113830, w_eco113831, w_eco113832, w_eco113833, w_eco113834, w_eco113835, w_eco113836, w_eco113837, w_eco113838, w_eco113839, w_eco113840, w_eco113841, w_eco113842, w_eco113843, w_eco113844, w_eco113845, w_eco113846, w_eco113847, w_eco113848, w_eco113849, w_eco113850, w_eco113851, w_eco113852, w_eco113853, w_eco113854, w_eco113855, w_eco113856, w_eco113857, w_eco113858, w_eco113859, w_eco113860, w_eco113861, w_eco113862, w_eco113863, w_eco113864, w_eco113865, w_eco113866, w_eco113867, w_eco113868, w_eco113869, w_eco113870, w_eco113871, w_eco113872, w_eco113873, w_eco113874, w_eco113875, w_eco113876, w_eco113877, w_eco113878, w_eco113879, w_eco113880, w_eco113881, w_eco113882, w_eco113883, w_eco113884, w_eco113885, w_eco113886, w_eco113887, w_eco113888, w_eco113889, w_eco113890, w_eco113891, w_eco113892, w_eco113893, w_eco113894, w_eco113895, w_eco113896, w_eco113897, w_eco113898, w_eco113899, w_eco113900, w_eco113901, w_eco113902, w_eco113903, w_eco113904, w_eco113905, w_eco113906, w_eco113907, w_eco113908, w_eco113909, w_eco113910, w_eco113911, w_eco113912, w_eco113913, w_eco113914, w_eco113915, w_eco113916, w_eco113917, w_eco113918, w_eco113919, w_eco113920, w_eco113921, w_eco113922, w_eco113923, w_eco113924, w_eco113925, w_eco113926, w_eco113927, w_eco113928, w_eco113929, w_eco113930, w_eco113931, w_eco113932, w_eco113933, w_eco113934, w_eco113935, w_eco113936, w_eco113937, w_eco113938, w_eco113939, w_eco113940, w_eco113941, w_eco113942, w_eco113943, w_eco113944, w_eco113945, w_eco113946, w_eco113947, w_eco113948, w_eco113949, w_eco113950, w_eco113951, w_eco113952, w_eco113953, w_eco113954, w_eco113955, w_eco113956, w_eco113957, w_eco113958, w_eco113959, w_eco113960, w_eco113961, w_eco113962, w_eco113963, w_eco113964, w_eco113965, w_eco113966, w_eco113967, w_eco113968, w_eco113969, w_eco113970, w_eco113971, w_eco113972, w_eco113973, w_eco113974, w_eco113975, w_eco113976, w_eco113977, w_eco113978, w_eco113979, w_eco113980, w_eco113981, w_eco113982, w_eco113983, w_eco113984, w_eco113985, w_eco113986, w_eco113987, w_eco113988, w_eco113989, w_eco113990, w_eco113991, w_eco113992, w_eco113993, w_eco113994, w_eco113995, w_eco113996, w_eco113997, w_eco113998, w_eco113999, w_eco114000, w_eco114001, w_eco114002, w_eco114003, w_eco114004, w_eco114005, w_eco114006, w_eco114007, w_eco114008, w_eco114009, w_eco114010, w_eco114011, w_eco114012, w_eco114013, w_eco114014, w_eco114015, w_eco114016, w_eco114017, w_eco114018, w_eco114019, w_eco114020, w_eco114021, w_eco114022, w_eco114023, w_eco114024, w_eco114025, w_eco114026, w_eco114027, w_eco114028, w_eco114029, w_eco114030, w_eco114031, w_eco114032, w_eco114033, w_eco114034, w_eco114035, w_eco114036, w_eco114037, w_eco114038, w_eco114039, w_eco114040, w_eco114041, w_eco114042, w_eco114043, w_eco114044, w_eco114045, w_eco114046, w_eco114047, w_eco114048, w_eco114049, w_eco114050, w_eco114051, w_eco114052, w_eco114053, w_eco114054, w_eco114055, w_eco114056, w_eco114057, w_eco114058, w_eco114059, w_eco114060, w_eco114061, w_eco114062, w_eco114063, w_eco114064, w_eco114065, w_eco114066, w_eco114067, w_eco114068, w_eco114069, w_eco114070, w_eco114071, w_eco114072, w_eco114073, w_eco114074, w_eco114075, w_eco114076, w_eco114077, w_eco114078, w_eco114079, w_eco114080, w_eco114081, w_eco114082, w_eco114083, w_eco114084, w_eco114085, w_eco114086, w_eco114087, w_eco114088, w_eco114089, w_eco114090, w_eco114091, w_eco114092, w_eco114093, w_eco114094, w_eco114095, w_eco114096, w_eco114097, w_eco114098, w_eco114099, w_eco114100, w_eco114101, w_eco114102, w_eco114103, w_eco114104, w_eco114105, w_eco114106, w_eco114107, w_eco114108, w_eco114109, w_eco114110, w_eco114111, w_eco114112, w_eco114113, w_eco114114, w_eco114115, w_eco114116, w_eco114117, w_eco114118, w_eco114119, w_eco114120, w_eco114121, w_eco114122, w_eco114123, w_eco114124, w_eco114125, w_eco114126, w_eco114127, w_eco114128, w_eco114129, w_eco114130, w_eco114131, w_eco114132, w_eco114133, w_eco114134, w_eco114135, w_eco114136, w_eco114137, w_eco114138, w_eco114139, w_eco114140, w_eco114141, w_eco114142, w_eco114143, w_eco114144, w_eco114145, w_eco114146, w_eco114147, w_eco114148, w_eco114149, w_eco114150, w_eco114151, w_eco114152, w_eco114153, w_eco114154, w_eco114155, w_eco114156, w_eco114157, w_eco114158, w_eco114159, w_eco114160, w_eco114161, w_eco114162, w_eco114163, w_eco114164, w_eco114165, w_eco114166, w_eco114167, w_eco114168, w_eco114169, w_eco114170, w_eco114171, w_eco114172, w_eco114173, w_eco114174, w_eco114175, w_eco114176, w_eco114177, w_eco114178, w_eco114179, w_eco114180, w_eco114181, w_eco114182, w_eco114183, w_eco114184, w_eco114185, w_eco114186, w_eco114187, w_eco114188, w_eco114189, w_eco114190, w_eco114191, w_eco114192, w_eco114193, w_eco114194, w_eco114195, w_eco114196, w_eco114197, w_eco114198, w_eco114199, w_eco114200, w_eco114201, w_eco114202, w_eco114203, w_eco114204, w_eco114205, w_eco114206, w_eco114207, w_eco114208, w_eco114209, w_eco114210, w_eco114211, w_eco114212, w_eco114213, w_eco114214, w_eco114215, w_eco114216, w_eco114217, w_eco114218, w_eco114219, w_eco114220, w_eco114221, w_eco114222, w_eco114223, w_eco114224, w_eco114225, w_eco114226, w_eco114227, w_eco114228, w_eco114229, w_eco114230, w_eco114231, w_eco114232, w_eco114233, w_eco114234, w_eco114235, w_eco114236, w_eco114237, w_eco114238, w_eco114239, w_eco114240, w_eco114241, w_eco114242, w_eco114243, w_eco114244, w_eco114245, w_eco114246, w_eco114247, w_eco114248, w_eco114249, w_eco114250, w_eco114251, w_eco114252, w_eco114253, w_eco114254, w_eco114255, w_eco114256, w_eco114257, w_eco114258, w_eco114259, w_eco114260, w_eco114261, w_eco114262, w_eco114263, w_eco114264, w_eco114265, w_eco114266, w_eco114267, w_eco114268, w_eco114269, w_eco114270, w_eco114271, w_eco114272, w_eco114273, w_eco114274, w_eco114275, w_eco114276, w_eco114277, w_eco114278, w_eco114279, w_eco114280, w_eco114281, w_eco114282, w_eco114283, w_eco114284, w_eco114285, w_eco114286, w_eco114287, w_eco114288, w_eco114289, w_eco114290, w_eco114291, w_eco114292, w_eco114293, w_eco114294, w_eco114295, w_eco114296, w_eco114297, w_eco114298, w_eco114299, w_eco114300, w_eco114301, w_eco114302, w_eco114303, w_eco114304, w_eco114305, w_eco114306, w_eco114307, w_eco114308, w_eco114309, w_eco114310, w_eco114311, w_eco114312, w_eco114313, w_eco114314, w_eco114315, w_eco114316, w_eco114317, w_eco114318, w_eco114319, w_eco114320, w_eco114321, w_eco114322, w_eco114323, w_eco114324, w_eco114325, w_eco114326, w_eco114327, w_eco114328, w_eco114329, w_eco114330, w_eco114331, w_eco114332, w_eco114333, w_eco114334, w_eco114335, w_eco114336, w_eco114337, w_eco114338, w_eco114339, w_eco114340, w_eco114341, w_eco114342, w_eco114343, w_eco114344, w_eco114345, w_eco114346, w_eco114347, w_eco114348, w_eco114349, w_eco114350, w_eco114351, w_eco114352, w_eco114353, w_eco114354, w_eco114355, w_eco114356, w_eco114357, w_eco114358, w_eco114359, w_eco114360, w_eco114361, w_eco114362, w_eco114363, w_eco114364, w_eco114365, w_eco114366, w_eco114367, w_eco114368, w_eco114369, w_eco114370, w_eco114371, w_eco114372, w_eco114373, w_eco114374, w_eco114375, w_eco114376, w_eco114377, w_eco114378, w_eco114379, w_eco114380, w_eco114381, w_eco114382, w_eco114383, w_eco114384, w_eco114385, w_eco114386, w_eco114387, w_eco114388, w_eco114389, w_eco114390, w_eco114391, w_eco114392, w_eco114393, w_eco114394, w_eco114395, w_eco114396, w_eco114397, w_eco114398, w_eco114399, w_eco114400, w_eco114401, w_eco114402, w_eco114403, w_eco114404, w_eco114405, w_eco114406, w_eco114407, w_eco114408, w_eco114409, w_eco114410, w_eco114411, w_eco114412, w_eco114413, w_eco114414, w_eco114415, w_eco114416, w_eco114417, w_eco114418, w_eco114419, w_eco114420, w_eco114421, w_eco114422, w_eco114423, w_eco114424, w_eco114425, w_eco114426, w_eco114427, w_eco114428, w_eco114429, w_eco114430, w_eco114431, w_eco114432, w_eco114433, w_eco114434, w_eco114435, w_eco114436, w_eco114437, w_eco114438, w_eco114439, w_eco114440, w_eco114441, w_eco114442, w_eco114443, w_eco114444, w_eco114445, w_eco114446, w_eco114447, w_eco114448, w_eco114449, w_eco114450, w_eco114451, w_eco114452, w_eco114453, w_eco114454, w_eco114455, w_eco114456, w_eco114457, w_eco114458, w_eco114459, w_eco114460, w_eco114461, w_eco114462, w_eco114463, w_eco114464, w_eco114465, w_eco114466, w_eco114467, w_eco114468, w_eco114469, w_eco114470, w_eco114471, w_eco114472, w_eco114473, w_eco114474, w_eco114475, w_eco114476, w_eco114477, w_eco114478, w_eco114479, w_eco114480, w_eco114481, w_eco114482, w_eco114483, w_eco114484, w_eco114485, w_eco114486, w_eco114487, w_eco114488, w_eco114489, w_eco114490, w_eco114491, w_eco114492, w_eco114493, w_eco114494, w_eco114495, w_eco114496, w_eco114497, w_eco114498, w_eco114499, w_eco114500, w_eco114501, w_eco114502, w_eco114503, w_eco114504, w_eco114505, w_eco114506, w_eco114507, w_eco114508, w_eco114509, w_eco114510, w_eco114511, w_eco114512, w_eco114513, w_eco114514, w_eco114515, w_eco114516, w_eco114517, w_eco114518, w_eco114519, w_eco114520, w_eco114521, w_eco114522, w_eco114523, w_eco114524, w_eco114525, w_eco114526, w_eco114527, w_eco114528, w_eco114529, w_eco114530, w_eco114531, w_eco114532, w_eco114533, w_eco114534, w_eco114535, w_eco114536, w_eco114537, w_eco114538, w_eco114539, w_eco114540, w_eco114541, w_eco114542, w_eco114543, w_eco114544, w_eco114545, w_eco114546, w_eco114547, w_eco114548, w_eco114549, w_eco114550, w_eco114551, w_eco114552, w_eco114553, w_eco114554, w_eco114555, w_eco114556, w_eco114557, w_eco114558, w_eco114559, w_eco114560, w_eco114561, w_eco114562, w_eco114563, w_eco114564, w_eco114565, w_eco114566, w_eco114567, w_eco114568, w_eco114569, w_eco114570, w_eco114571, w_eco114572, w_eco114573, w_eco114574, w_eco114575, w_eco114576, w_eco114577, w_eco114578, w_eco114579, w_eco114580, w_eco114581, w_eco114582, w_eco114583, w_eco114584, w_eco114585, w_eco114586, w_eco114587, w_eco114588, w_eco114589, w_eco114590, w_eco114591, w_eco114592, w_eco114593, w_eco114594, w_eco114595, w_eco114596, w_eco114597, w_eco114598, w_eco114599, w_eco114600, w_eco114601, w_eco114602, w_eco114603, w_eco114604, w_eco114605, w_eco114606, w_eco114607, w_eco114608, w_eco114609, w_eco114610, w_eco114611, w_eco114612, w_eco114613, w_eco114614, w_eco114615, w_eco114616, w_eco114617, w_eco114618, w_eco114619, w_eco114620, w_eco114621, w_eco114622, w_eco114623, w_eco114624, w_eco114625, w_eco114626, w_eco114627, w_eco114628, w_eco114629, w_eco114630, w_eco114631, w_eco114632, w_eco114633, w_eco114634, w_eco114635, w_eco114636, w_eco114637, w_eco114638, w_eco114639, w_eco114640, w_eco114641, w_eco114642, w_eco114643, w_eco114644, w_eco114645, w_eco114646, w_eco114647, w_eco114648, w_eco114649, w_eco114650, w_eco114651, w_eco114652, w_eco114653, w_eco114654, w_eco114655, w_eco114656, w_eco114657, w_eco114658, w_eco114659, w_eco114660, w_eco114661, w_eco114662, w_eco114663, w_eco114664, w_eco114665, w_eco114666, w_eco114667, w_eco114668, w_eco114669, w_eco114670, w_eco114671, w_eco114672, w_eco114673, w_eco114674, w_eco114675, w_eco114676, w_eco114677, w_eco114678, w_eco114679, w_eco114680, w_eco114681, w_eco114682, w_eco114683, w_eco114684, w_eco114685, w_eco114686, w_eco114687, w_eco114688, w_eco114689, w_eco114690, w_eco114691, w_eco114692, w_eco114693, w_eco114694, w_eco114695, w_eco114696, w_eco114697, w_eco114698, w_eco114699, w_eco114700, w_eco114701, w_eco114702, w_eco114703, w_eco114704, w_eco114705, w_eco114706, w_eco114707, w_eco114708, w_eco114709, w_eco114710, w_eco114711, w_eco114712, w_eco114713, w_eco114714, w_eco114715, w_eco114716, w_eco114717, w_eco114718, w_eco114719, w_eco114720, w_eco114721, w_eco114722, w_eco114723, w_eco114724, w_eco114725, w_eco114726, w_eco114727, w_eco114728, w_eco114729, w_eco114730, w_eco114731, w_eco114732, w_eco114733, w_eco114734, w_eco114735, w_eco114736, w_eco114737, w_eco114738, w_eco114739, w_eco114740, w_eco114741, w_eco114742, w_eco114743, w_eco114744, w_eco114745, w_eco114746, w_eco114747, w_eco114748, w_eco114749, w_eco114750, w_eco114751, w_eco114752, w_eco114753, w_eco114754, w_eco114755, w_eco114756, w_eco114757, w_eco114758, w_eco114759, w_eco114760, w_eco114761, w_eco114762, w_eco114763, w_eco114764, w_eco114765, w_eco114766, w_eco114767, w_eco114768, w_eco114769, w_eco114770, w_eco114771, w_eco114772, w_eco114773, w_eco114774, w_eco114775, w_eco114776, w_eco114777, w_eco114778, w_eco114779, w_eco114780, w_eco114781, w_eco114782, w_eco114783, w_eco114784, w_eco114785, w_eco114786, w_eco114787, w_eco114788, w_eco114789, w_eco114790, w_eco114791, w_eco114792, w_eco114793, w_eco114794, w_eco114795, w_eco114796, w_eco114797, w_eco114798, w_eco114799, w_eco114800, w_eco114801, w_eco114802, w_eco114803, w_eco114804, w_eco114805, w_eco114806, w_eco114807, w_eco114808, w_eco114809, w_eco114810, w_eco114811, w_eco114812, w_eco114813, w_eco114814, w_eco114815, w_eco114816, w_eco114817, w_eco114818, w_eco114819, w_eco114820, w_eco114821, w_eco114822, w_eco114823, w_eco114824, w_eco114825, w_eco114826, w_eco114827, w_eco114828, w_eco114829, w_eco114830, w_eco114831, w_eco114832, w_eco114833, w_eco114834, w_eco114835, w_eco114836, w_eco114837, w_eco114838, w_eco114839, w_eco114840, w_eco114841, w_eco114842, w_eco114843, w_eco114844, w_eco114845, w_eco114846, w_eco114847, w_eco114848, w_eco114849, w_eco114850, w_eco114851, w_eco114852, w_eco114853, w_eco114854, w_eco114855, w_eco114856, w_eco114857, w_eco114858, w_eco114859, w_eco114860, w_eco114861, w_eco114862, w_eco114863, w_eco114864, w_eco114865, w_eco114866, w_eco114867, w_eco114868, w_eco114869, w_eco114870, w_eco114871, w_eco114872, w_eco114873, w_eco114874, w_eco114875, w_eco114876, w_eco114877, w_eco114878, w_eco114879, w_eco114880, w_eco114881, w_eco114882, w_eco114883, w_eco114884, w_eco114885, w_eco114886, w_eco114887, w_eco114888, w_eco114889, w_eco114890, w_eco114891, w_eco114892, w_eco114893, w_eco114894, w_eco114895, w_eco114896, w_eco114897, w_eco114898, w_eco114899, w_eco114900, w_eco114901, w_eco114902, w_eco114903, w_eco114904, w_eco114905, w_eco114906, w_eco114907, w_eco114908, w_eco114909, w_eco114910, w_eco114911, w_eco114912, w_eco114913, w_eco114914, w_eco114915, w_eco114916, w_eco114917, w_eco114918, w_eco114919, w_eco114920, w_eco114921, w_eco114922, w_eco114923, w_eco114924, w_eco114925, w_eco114926, w_eco114927, w_eco114928, w_eco114929, w_eco114930, w_eco114931, w_eco114932, w_eco114933, w_eco114934, w_eco114935, w_eco114936, w_eco114937, w_eco114938, w_eco114939, w_eco114940, w_eco114941, w_eco114942, w_eco114943, w_eco114944, w_eco114945, w_eco114946, w_eco114947, w_eco114948, w_eco114949, w_eco114950, w_eco114951, w_eco114952, w_eco114953, w_eco114954, w_eco114955, w_eco114956, w_eco114957, w_eco114958, w_eco114959, w_eco114960, w_eco114961, w_eco114962, w_eco114963, w_eco114964, w_eco114965, w_eco114966, w_eco114967, w_eco114968, w_eco114969, w_eco114970, w_eco114971, w_eco114972, w_eco114973, w_eco114974, w_eco114975, w_eco114976, w_eco114977, w_eco114978, w_eco114979, w_eco114980, w_eco114981, w_eco114982, w_eco114983, w_eco114984, w_eco114985, w_eco114986, w_eco114987, w_eco114988, w_eco114989, w_eco114990, w_eco114991, w_eco114992, w_eco114993, w_eco114994, w_eco114995, w_eco114996, w_eco114997, w_eco114998, w_eco114999, w_eco115000, w_eco115001, w_eco115002, w_eco115003, w_eco115004, w_eco115005, w_eco115006, w_eco115007, w_eco115008, w_eco115009, w_eco115010, w_eco115011, w_eco115012, w_eco115013, w_eco115014, w_eco115015, w_eco115016, w_eco115017, w_eco115018, w_eco115019, w_eco115020, w_eco115021, w_eco115022, w_eco115023, w_eco115024, w_eco115025, w_eco115026, w_eco115027, w_eco115028, w_eco115029, w_eco115030, w_eco115031, w_eco115032, w_eco115033, w_eco115034, w_eco115035, w_eco115036, w_eco115037, w_eco115038, w_eco115039, w_eco115040, w_eco115041, w_eco115042, w_eco115043, w_eco115044, w_eco115045, w_eco115046, w_eco115047, w_eco115048, w_eco115049, w_eco115050, w_eco115051, w_eco115052, w_eco115053, w_eco115054, w_eco115055, w_eco115056, w_eco115057, w_eco115058, w_eco115059, w_eco115060, w_eco115061, w_eco115062, w_eco115063, w_eco115064, w_eco115065, w_eco115066, w_eco115067, w_eco115068, w_eco115069, w_eco115070, w_eco115071, w_eco115072, w_eco115073, w_eco115074, w_eco115075, w_eco115076, w_eco115077, w_eco115078, w_eco115079, w_eco115080, w_eco115081, w_eco115082, w_eco115083, w_eco115084, w_eco115085, w_eco115086, w_eco115087, w_eco115088, w_eco115089, w_eco115090, w_eco115091, w_eco115092, w_eco115093, w_eco115094, w_eco115095, w_eco115096, w_eco115097, w_eco115098, w_eco115099, w_eco115100, w_eco115101, w_eco115102, w_eco115103, w_eco115104, w_eco115105, w_eco115106, w_eco115107, w_eco115108, w_eco115109, w_eco115110, w_eco115111, w_eco115112, w_eco115113, w_eco115114, w_eco115115, w_eco115116, w_eco115117, w_eco115118, w_eco115119, w_eco115120, w_eco115121, w_eco115122, w_eco115123, w_eco115124, w_eco115125, w_eco115126, w_eco115127, w_eco115128, w_eco115129, w_eco115130, w_eco115131, w_eco115132, w_eco115133, w_eco115134, w_eco115135, w_eco115136, w_eco115137, w_eco115138, w_eco115139, w_eco115140, w_eco115141, w_eco115142, w_eco115143, w_eco115144, w_eco115145, w_eco115146, w_eco115147, w_eco115148, w_eco115149, w_eco115150, w_eco115151, w_eco115152, w_eco115153, w_eco115154, w_eco115155, w_eco115156, w_eco115157, w_eco115158, w_eco115159, w_eco115160, w_eco115161, w_eco115162, w_eco115163, w_eco115164, w_eco115165, w_eco115166, w_eco115167, w_eco115168, w_eco115169, w_eco115170, w_eco115171, w_eco115172, w_eco115173, w_eco115174, w_eco115175, w_eco115176, w_eco115177, w_eco115178, w_eco115179, w_eco115180, w_eco115181, w_eco115182, w_eco115183, w_eco115184, w_eco115185, w_eco115186, w_eco115187, w_eco115188, w_eco115189, w_eco115190, w_eco115191, w_eco115192, w_eco115193, w_eco115194, w_eco115195, w_eco115196, w_eco115197, w_eco115198, w_eco115199, w_eco115200, w_eco115201, w_eco115202, w_eco115203, w_eco115204, w_eco115205, w_eco115206, w_eco115207, w_eco115208, w_eco115209, w_eco115210, w_eco115211, w_eco115212, w_eco115213, w_eco115214, w_eco115215, w_eco115216, w_eco115217, w_eco115218, w_eco115219, w_eco115220, w_eco115221, w_eco115222, w_eco115223, w_eco115224, w_eco115225, w_eco115226, w_eco115227, w_eco115228, w_eco115229, w_eco115230, w_eco115231, w_eco115232, w_eco115233, w_eco115234, w_eco115235, w_eco115236, w_eco115237, w_eco115238, w_eco115239, w_eco115240, w_eco115241, w_eco115242, w_eco115243, w_eco115244, w_eco115245, w_eco115246, w_eco115247, w_eco115248, w_eco115249, w_eco115250, w_eco115251, w_eco115252, w_eco115253, w_eco115254, w_eco115255, w_eco115256, w_eco115257, w_eco115258, w_eco115259, w_eco115260, w_eco115261, w_eco115262, w_eco115263, w_eco115264, w_eco115265, w_eco115266, w_eco115267, w_eco115268, w_eco115269, w_eco115270, w_eco115271, w_eco115272, w_eco115273, w_eco115274, w_eco115275, w_eco115276, w_eco115277, w_eco115278, w_eco115279, w_eco115280, w_eco115281, w_eco115282, w_eco115283, w_eco115284, w_eco115285, w_eco115286, w_eco115287, w_eco115288, w_eco115289, w_eco115290, w_eco115291, w_eco115292, w_eco115293, w_eco115294, w_eco115295, w_eco115296, w_eco115297, w_eco115298, w_eco115299, w_eco115300, w_eco115301, w_eco115302, w_eco115303, w_eco115304, w_eco115305, w_eco115306, w_eco115307, w_eco115308, w_eco115309, w_eco115310, w_eco115311, w_eco115312, w_eco115313, w_eco115314, w_eco115315, w_eco115316, w_eco115317, w_eco115318, w_eco115319, w_eco115320, w_eco115321, w_eco115322, w_eco115323, w_eco115324, w_eco115325, w_eco115326, w_eco115327, w_eco115328, w_eco115329, w_eco115330, w_eco115331, w_eco115332, w_eco115333, w_eco115334, w_eco115335, w_eco115336, w_eco115337, w_eco115338, w_eco115339, w_eco115340, w_eco115341, w_eco115342, w_eco115343, w_eco115344, w_eco115345, w_eco115346, w_eco115347, w_eco115348, w_eco115349, w_eco115350, w_eco115351, w_eco115352, w_eco115353, w_eco115354, w_eco115355, w_eco115356, w_eco115357, w_eco115358, w_eco115359, w_eco115360, w_eco115361, w_eco115362, w_eco115363, w_eco115364, w_eco115365, w_eco115366, w_eco115367, w_eco115368, w_eco115369, w_eco115370, w_eco115371, w_eco115372, w_eco115373, w_eco115374, w_eco115375, w_eco115376, w_eco115377, w_eco115378, w_eco115379, w_eco115380, w_eco115381, w_eco115382, w_eco115383, w_eco115384, w_eco115385, w_eco115386, w_eco115387, w_eco115388, w_eco115389, w_eco115390, w_eco115391, w_eco115392, w_eco115393, w_eco115394, w_eco115395, w_eco115396, w_eco115397, w_eco115398, w_eco115399, w_eco115400, w_eco115401, w_eco115402, w_eco115403, w_eco115404, w_eco115405, w_eco115406, w_eco115407, w_eco115408, w_eco115409, w_eco115410, w_eco115411, w_eco115412, w_eco115413, w_eco115414, w_eco115415, w_eco115416, w_eco115417, w_eco115418, w_eco115419, w_eco115420, w_eco115421, w_eco115422, w_eco115423, w_eco115424, w_eco115425, w_eco115426, w_eco115427, w_eco115428, w_eco115429, w_eco115430, w_eco115431, w_eco115432, w_eco115433, w_eco115434, w_eco115435, w_eco115436, w_eco115437, w_eco115438, w_eco115439, w_eco115440, w_eco115441, w_eco115442, w_eco115443, w_eco115444, w_eco115445, w_eco115446, w_eco115447, w_eco115448, w_eco115449, w_eco115450, w_eco115451, w_eco115452, w_eco115453, w_eco115454, w_eco115455, w_eco115456, w_eco115457, w_eco115458, w_eco115459, w_eco115460, w_eco115461, w_eco115462, w_eco115463, w_eco115464, w_eco115465, w_eco115466, w_eco115467, w_eco115468, w_eco115469, w_eco115470, w_eco115471, w_eco115472, w_eco115473, w_eco115474, w_eco115475, w_eco115476, w_eco115477, w_eco115478, w_eco115479, w_eco115480, w_eco115481, w_eco115482, w_eco115483, w_eco115484, w_eco115485, w_eco115486, w_eco115487, w_eco115488, w_eco115489, w_eco115490, w_eco115491, w_eco115492, w_eco115493, w_eco115494, w_eco115495, w_eco115496, w_eco115497, w_eco115498, w_eco115499, w_eco115500, w_eco115501, w_eco115502, w_eco115503, w_eco115504, w_eco115505, w_eco115506, w_eco115507, w_eco115508, w_eco115509, w_eco115510, w_eco115511, w_eco115512, w_eco115513, w_eco115514, w_eco115515, w_eco115516, w_eco115517, w_eco115518, w_eco115519, w_eco115520, w_eco115521, w_eco115522, w_eco115523, w_eco115524, w_eco115525, w_eco115526, w_eco115527, w_eco115528, w_eco115529, w_eco115530, w_eco115531, w_eco115532, w_eco115533, w_eco115534, w_eco115535, w_eco115536, w_eco115537, w_eco115538, w_eco115539, w_eco115540, w_eco115541, w_eco115542, w_eco115543, w_eco115544, w_eco115545, w_eco115546, w_eco115547, w_eco115548, w_eco115549, w_eco115550, w_eco115551, w_eco115552, w_eco115553, w_eco115554, w_eco115555, w_eco115556, w_eco115557, w_eco115558, w_eco115559, w_eco115560, w_eco115561, w_eco115562, w_eco115563, w_eco115564, w_eco115565, w_eco115566, w_eco115567, w_eco115568, w_eco115569, w_eco115570, w_eco115571, w_eco115572, w_eco115573, w_eco115574, w_eco115575, w_eco115576, w_eco115577, w_eco115578, w_eco115579, w_eco115580, w_eco115581, w_eco115582, w_eco115583, w_eco115584, w_eco115585, w_eco115586, w_eco115587, w_eco115588, w_eco115589, w_eco115590, w_eco115591, w_eco115592, w_eco115593, w_eco115594, w_eco115595, w_eco115596, w_eco115597, w_eco115598, w_eco115599, w_eco115600, w_eco115601, w_eco115602, w_eco115603, w_eco115604, w_eco115605, w_eco115606, w_eco115607, w_eco115608, w_eco115609, w_eco115610, w_eco115611, w_eco115612, w_eco115613, w_eco115614, w_eco115615, w_eco115616, w_eco115617, w_eco115618, w_eco115619, w_eco115620, w_eco115621, w_eco115622, w_eco115623, w_eco115624, w_eco115625, w_eco115626, w_eco115627, w_eco115628, w_eco115629, w_eco115630, w_eco115631, w_eco115632, w_eco115633, w_eco115634, w_eco115635, w_eco115636, w_eco115637, w_eco115638, w_eco115639, w_eco115640, w_eco115641, w_eco115642, w_eco115643, w_eco115644, w_eco115645, w_eco115646, w_eco115647, w_eco115648, w_eco115649, w_eco115650, w_eco115651, w_eco115652, w_eco115653, w_eco115654, w_eco115655, w_eco115656, w_eco115657, w_eco115658, w_eco115659, w_eco115660, w_eco115661, w_eco115662, w_eco115663, w_eco115664, w_eco115665, w_eco115666, w_eco115667, w_eco115668, w_eco115669, w_eco115670, w_eco115671, w_eco115672, w_eco115673, w_eco115674, w_eco115675, w_eco115676, w_eco115677, w_eco115678, w_eco115679, w_eco115680, w_eco115681, w_eco115682, w_eco115683, w_eco115684, w_eco115685, w_eco115686, w_eco115687, w_eco115688, w_eco115689, w_eco115690, w_eco115691, w_eco115692, w_eco115693, w_eco115694, w_eco115695, w_eco115696, w_eco115697, w_eco115698, w_eco115699, w_eco115700, w_eco115701, w_eco115702, w_eco115703, w_eco115704, w_eco115705, w_eco115706, w_eco115707, w_eco115708, w_eco115709, w_eco115710, w_eco115711, w_eco115712, w_eco115713, w_eco115714, w_eco115715, w_eco115716, w_eco115717, w_eco115718, w_eco115719, w_eco115720, w_eco115721, w_eco115722, w_eco115723, w_eco115724, w_eco115725, w_eco115726, w_eco115727, w_eco115728, w_eco115729, w_eco115730, w_eco115731, w_eco115732, w_eco115733, w_eco115734, w_eco115735, w_eco115736, w_eco115737, w_eco115738, w_eco115739, w_eco115740, w_eco115741, w_eco115742, w_eco115743, w_eco115744, w_eco115745, w_eco115746, w_eco115747, w_eco115748, w_eco115749, w_eco115750, w_eco115751, w_eco115752, w_eco115753, w_eco115754, w_eco115755, w_eco115756, w_eco115757, w_eco115758, w_eco115759, w_eco115760, w_eco115761, w_eco115762, w_eco115763, w_eco115764, w_eco115765, w_eco115766, w_eco115767, w_eco115768, w_eco115769, w_eco115770, w_eco115771, w_eco115772, w_eco115773, w_eco115774, w_eco115775, w_eco115776, w_eco115777, w_eco115778, w_eco115779, w_eco115780, w_eco115781, w_eco115782, w_eco115783, w_eco115784, w_eco115785, w_eco115786, w_eco115787, w_eco115788, w_eco115789, w_eco115790, w_eco115791, w_eco115792, w_eco115793, w_eco115794, w_eco115795, w_eco115796, w_eco115797, w_eco115798, w_eco115799, w_eco115800, w_eco115801, w_eco115802, w_eco115803, w_eco115804, w_eco115805, w_eco115806, w_eco115807, w_eco115808, w_eco115809, w_eco115810, w_eco115811, w_eco115812, w_eco115813, w_eco115814, w_eco115815, w_eco115816, w_eco115817, w_eco115818, w_eco115819, w_eco115820, w_eco115821, w_eco115822, w_eco115823, w_eco115824, w_eco115825, w_eco115826, w_eco115827, w_eco115828, w_eco115829, w_eco115830, w_eco115831, w_eco115832, w_eco115833, w_eco115834, w_eco115835, w_eco115836, w_eco115837, w_eco115838, w_eco115839, w_eco115840, w_eco115841, w_eco115842, w_eco115843, w_eco115844, w_eco115845, w_eco115846, w_eco115847, w_eco115848, w_eco115849, w_eco115850, w_eco115851, w_eco115852, w_eco115853, w_eco115854, w_eco115855, w_eco115856, w_eco115857, w_eco115858, w_eco115859, w_eco115860, w_eco115861, w_eco115862, w_eco115863, w_eco115864, w_eco115865, w_eco115866, w_eco115867, w_eco115868, w_eco115869, w_eco115870, w_eco115871, w_eco115872, w_eco115873, w_eco115874, w_eco115875, w_eco115876, w_eco115877, w_eco115878, w_eco115879, w_eco115880, w_eco115881, w_eco115882, w_eco115883, w_eco115884, w_eco115885, w_eco115886, w_eco115887, w_eco115888, w_eco115889, w_eco115890, w_eco115891, w_eco115892, w_eco115893, w_eco115894, w_eco115895, w_eco115896, w_eco115897, w_eco115898, w_eco115899, w_eco115900, w_eco115901, w_eco115902, w_eco115903, w_eco115904, w_eco115905, w_eco115906, w_eco115907, w_eco115908, w_eco115909, w_eco115910, w_eco115911, w_eco115912, w_eco115913, w_eco115914, w_eco115915, w_eco115916, w_eco115917, w_eco115918, w_eco115919, w_eco115920, w_eco115921, w_eco115922, w_eco115923, w_eco115924, w_eco115925, w_eco115926, w_eco115927, w_eco115928, w_eco115929, w_eco115930, w_eco115931, w_eco115932, w_eco115933, w_eco115934, w_eco115935, w_eco115936, w_eco115937, w_eco115938, w_eco115939, w_eco115940, w_eco115941, w_eco115942, w_eco115943, w_eco115944, w_eco115945, w_eco115946, w_eco115947, w_eco115948, w_eco115949, w_eco115950, w_eco115951, w_eco115952, w_eco115953, w_eco115954, w_eco115955, w_eco115956, w_eco115957, w_eco115958, w_eco115959, w_eco115960, w_eco115961, w_eco115962, w_eco115963, w_eco115964, w_eco115965, w_eco115966, w_eco115967, w_eco115968, w_eco115969, w_eco115970, w_eco115971, w_eco115972, w_eco115973, w_eco115974, w_eco115975, w_eco115976, w_eco115977, w_eco115978, w_eco115979, w_eco115980, w_eco115981, w_eco115982, w_eco115983, w_eco115984, w_eco115985, w_eco115986, w_eco115987, w_eco115988, w_eco115989, w_eco115990, w_eco115991, w_eco115992, w_eco115993, w_eco115994, w_eco115995, w_eco115996, w_eco115997, w_eco115998, w_eco115999, w_eco116000, w_eco116001, w_eco116002, w_eco116003, w_eco116004, w_eco116005, w_eco116006, w_eco116007, w_eco116008, w_eco116009, w_eco116010, w_eco116011, w_eco116012, w_eco116013, w_eco116014, w_eco116015, w_eco116016, w_eco116017, w_eco116018, w_eco116019, w_eco116020, w_eco116021, w_eco116022, w_eco116023, w_eco116024, w_eco116025, w_eco116026, w_eco116027, w_eco116028, w_eco116029, w_eco116030, w_eco116031, w_eco116032, w_eco116033, w_eco116034, w_eco116035, w_eco116036, w_eco116037, w_eco116038, w_eco116039, w_eco116040, w_eco116041, w_eco116042, w_eco116043, w_eco116044, w_eco116045, w_eco116046, w_eco116047, w_eco116048, w_eco116049, w_eco116050, w_eco116051, w_eco116052, w_eco116053, w_eco116054, w_eco116055, w_eco116056, w_eco116057, w_eco116058, w_eco116059, w_eco116060, w_eco116061, w_eco116062, w_eco116063, w_eco116064, w_eco116065, w_eco116066, w_eco116067, w_eco116068, w_eco116069, w_eco116070, w_eco116071, w_eco116072, w_eco116073, w_eco116074, w_eco116075, w_eco116076, w_eco116077, w_eco116078, w_eco116079, w_eco116080, w_eco116081, w_eco116082, w_eco116083, w_eco116084, w_eco116085, w_eco116086, w_eco116087, w_eco116088, w_eco116089, w_eco116090, w_eco116091, w_eco116092, w_eco116093, w_eco116094, w_eco116095, w_eco116096, w_eco116097, w_eco116098, w_eco116099, w_eco116100, w_eco116101, w_eco116102, w_eco116103, w_eco116104, w_eco116105, w_eco116106, w_eco116107, w_eco116108, w_eco116109, w_eco116110, w_eco116111, w_eco116112, w_eco116113, w_eco116114, w_eco116115, w_eco116116, w_eco116117, w_eco116118, w_eco116119, w_eco116120, w_eco116121, w_eco116122, w_eco116123, w_eco116124, w_eco116125, w_eco116126, w_eco116127, w_eco116128, w_eco116129, w_eco116130, w_eco116131, w_eco116132, w_eco116133, w_eco116134, w_eco116135, w_eco116136, w_eco116137, w_eco116138, w_eco116139, w_eco116140, w_eco116141, w_eco116142, w_eco116143, w_eco116144, w_eco116145, w_eco116146, w_eco116147, w_eco116148, w_eco116149, w_eco116150, w_eco116151, w_eco116152, w_eco116153, w_eco116154, w_eco116155, w_eco116156, w_eco116157, w_eco116158, w_eco116159, w_eco116160, w_eco116161, w_eco116162, w_eco116163, w_eco116164, w_eco116165, w_eco116166, w_eco116167, w_eco116168, w_eco116169, w_eco116170, w_eco116171, w_eco116172, w_eco116173, w_eco116174, w_eco116175, w_eco116176, w_eco116177, w_eco116178, w_eco116179, w_eco116180, w_eco116181, w_eco116182, w_eco116183, w_eco116184, w_eco116185, w_eco116186, w_eco116187, w_eco116188, w_eco116189, w_eco116190, w_eco116191, w_eco116192, w_eco116193, w_eco116194, w_eco116195, w_eco116196, w_eco116197, w_eco116198, w_eco116199, w_eco116200, w_eco116201, w_eco116202, w_eco116203, w_eco116204, w_eco116205, w_eco116206, w_eco116207, w_eco116208, w_eco116209, w_eco116210, w_eco116211, w_eco116212, w_eco116213, w_eco116214, w_eco116215, w_eco116216, w_eco116217, w_eco116218, w_eco116219, w_eco116220, w_eco116221, w_eco116222, w_eco116223, w_eco116224, w_eco116225, w_eco116226, w_eco116227, w_eco116228, w_eco116229, w_eco116230, w_eco116231, w_eco116232, w_eco116233, w_eco116234, w_eco116235, w_eco116236, w_eco116237, w_eco116238, w_eco116239, w_eco116240, w_eco116241, w_eco116242, w_eco116243, w_eco116244, w_eco116245, w_eco116246, w_eco116247, w_eco116248, w_eco116249, w_eco116250, w_eco116251, w_eco116252, w_eco116253, w_eco116254, w_eco116255, w_eco116256, w_eco116257, w_eco116258, w_eco116259, w_eco116260, w_eco116261, w_eco116262, w_eco116263, w_eco116264, w_eco116265, w_eco116266, w_eco116267, w_eco116268, w_eco116269, w_eco116270, w_eco116271, w_eco116272, w_eco116273, w_eco116274, w_eco116275, w_eco116276, w_eco116277, w_eco116278, w_eco116279, w_eco116280, w_eco116281, w_eco116282, w_eco116283, w_eco116284, w_eco116285, w_eco116286, w_eco116287, w_eco116288, w_eco116289, w_eco116290, w_eco116291, w_eco116292, w_eco116293, w_eco116294, w_eco116295, w_eco116296, w_eco116297, w_eco116298, w_eco116299, w_eco116300, w_eco116301, w_eco116302, w_eco116303, w_eco116304, w_eco116305, w_eco116306, w_eco116307, w_eco116308, w_eco116309, w_eco116310, w_eco116311, w_eco116312, w_eco116313, w_eco116314, w_eco116315, w_eco116316, w_eco116317, w_eco116318, w_eco116319, w_eco116320, w_eco116321, w_eco116322, w_eco116323, w_eco116324, w_eco116325, w_eco116326, w_eco116327, w_eco116328, w_eco116329, w_eco116330, w_eco116331, w_eco116332, w_eco116333, w_eco116334, w_eco116335, w_eco116336, w_eco116337, w_eco116338, w_eco116339, w_eco116340, w_eco116341, w_eco116342, w_eco116343, w_eco116344, w_eco116345, w_eco116346, w_eco116347, w_eco116348, w_eco116349, w_eco116350, w_eco116351, w_eco116352, w_eco116353, w_eco116354, w_eco116355, w_eco116356, w_eco116357, w_eco116358, w_eco116359, w_eco116360, w_eco116361, w_eco116362, w_eco116363, w_eco116364, w_eco116365, w_eco116366, w_eco116367, w_eco116368, w_eco116369, w_eco116370, w_eco116371, w_eco116372, w_eco116373, w_eco116374, w_eco116375, w_eco116376, w_eco116377, w_eco116378, w_eco116379, w_eco116380, w_eco116381, w_eco116382, w_eco116383, w_eco116384, w_eco116385, w_eco116386, w_eco116387, w_eco116388, w_eco116389, w_eco116390, w_eco116391, w_eco116392, w_eco116393, w_eco116394, w_eco116395, w_eco116396, w_eco116397, w_eco116398, w_eco116399, w_eco116400, w_eco116401, w_eco116402, w_eco116403, w_eco116404, w_eco116405, w_eco116406, w_eco116407, w_eco116408, w_eco116409, w_eco116410, w_eco116411, w_eco116412, w_eco116413, w_eco116414, w_eco116415, w_eco116416, w_eco116417, w_eco116418, w_eco116419, w_eco116420, w_eco116421, w_eco116422, w_eco116423, w_eco116424, w_eco116425, w_eco116426, w_eco116427, w_eco116428, w_eco116429, w_eco116430, w_eco116431, w_eco116432, w_eco116433, w_eco116434, w_eco116435, w_eco116436, w_eco116437, w_eco116438, w_eco116439, w_eco116440, w_eco116441, w_eco116442, w_eco116443, w_eco116444, w_eco116445, w_eco116446, w_eco116447, w_eco116448, w_eco116449, w_eco116450, w_eco116451, w_eco116452, w_eco116453, w_eco116454, w_eco116455, w_eco116456, w_eco116457, w_eco116458, w_eco116459, w_eco116460, w_eco116461, w_eco116462, w_eco116463, w_eco116464, w_eco116465, w_eco116466, w_eco116467, w_eco116468, w_eco116469, w_eco116470, w_eco116471, w_eco116472, w_eco116473, w_eco116474, w_eco116475, w_eco116476, w_eco116477, w_eco116478, w_eco116479, w_eco116480, w_eco116481, w_eco116482, w_eco116483, w_eco116484, w_eco116485, w_eco116486, w_eco116487, w_eco116488, w_eco116489, w_eco116490, w_eco116491, w_eco116492, w_eco116493, w_eco116494, w_eco116495, w_eco116496, w_eco116497, w_eco116498, w_eco116499, w_eco116500, w_eco116501, w_eco116502, w_eco116503, w_eco116504, w_eco116505, w_eco116506, w_eco116507, w_eco116508, w_eco116509, w_eco116510, w_eco116511, w_eco116512, w_eco116513, w_eco116514, w_eco116515, w_eco116516, w_eco116517, w_eco116518, w_eco116519, w_eco116520, w_eco116521, w_eco116522, w_eco116523, w_eco116524, w_eco116525, w_eco116526, w_eco116527, w_eco116528, w_eco116529, w_eco116530, w_eco116531, w_eco116532, w_eco116533, w_eco116534, w_eco116535, w_eco116536, w_eco116537, w_eco116538, w_eco116539, w_eco116540, w_eco116541, w_eco116542, w_eco116543, w_eco116544, w_eco116545, w_eco116546, w_eco116547, w_eco116548, w_eco116549, w_eco116550, w_eco116551, w_eco116552, w_eco116553, w_eco116554, w_eco116555, w_eco116556, w_eco116557, w_eco116558, w_eco116559, w_eco116560, w_eco116561, w_eco116562, w_eco116563, w_eco116564, w_eco116565, w_eco116566, w_eco116567, w_eco116568, w_eco116569, w_eco116570, w_eco116571, w_eco116572, w_eco116573, w_eco116574, w_eco116575, w_eco116576, w_eco116577, w_eco116578, w_eco116579, w_eco116580, w_eco116581, w_eco116582, w_eco116583, w_eco116584, w_eco116585, w_eco116586, w_eco116587, w_eco116588, w_eco116589, w_eco116590, w_eco116591, w_eco116592, w_eco116593, w_eco116594, w_eco116595, w_eco116596, w_eco116597, w_eco116598, w_eco116599, w_eco116600, w_eco116601, w_eco116602, w_eco116603, w_eco116604, w_eco116605, w_eco116606, w_eco116607, w_eco116608, w_eco116609, w_eco116610, w_eco116611, w_eco116612, w_eco116613, w_eco116614, w_eco116615, w_eco116616, w_eco116617, w_eco116618, w_eco116619, w_eco116620, w_eco116621, w_eco116622, w_eco116623, w_eco116624, w_eco116625, w_eco116626, w_eco116627, w_eco116628, w_eco116629, w_eco116630, w_eco116631, w_eco116632, w_eco116633, w_eco116634, w_eco116635, w_eco116636, w_eco116637, w_eco116638, w_eco116639, w_eco116640, w_eco116641, w_eco116642, w_eco116643, w_eco116644, w_eco116645, w_eco116646, w_eco116647, w_eco116648, w_eco116649, w_eco116650, w_eco116651, w_eco116652, w_eco116653, w_eco116654, w_eco116655, w_eco116656, w_eco116657, w_eco116658, w_eco116659, w_eco116660, w_eco116661, w_eco116662, w_eco116663, w_eco116664, w_eco116665, w_eco116666, w_eco116667, w_eco116668, w_eco116669, w_eco116670, w_eco116671, w_eco116672, w_eco116673, w_eco116674, w_eco116675, w_eco116676, w_eco116677, w_eco116678, w_eco116679, w_eco116680, w_eco116681, w_eco116682, w_eco116683, w_eco116684, w_eco116685, w_eco116686, w_eco116687, w_eco116688, w_eco116689, w_eco116690, w_eco116691, w_eco116692, w_eco116693, w_eco116694, w_eco116695, w_eco116696, w_eco116697, w_eco116698, w_eco116699, w_eco116700, w_eco116701, w_eco116702, w_eco116703, w_eco116704, w_eco116705, w_eco116706, w_eco116707, w_eco116708, w_eco116709, w_eco116710, w_eco116711, w_eco116712, w_eco116713, w_eco116714, w_eco116715, w_eco116716, w_eco116717, w_eco116718, w_eco116719, w_eco116720, w_eco116721, w_eco116722, w_eco116723, w_eco116724, w_eco116725, w_eco116726, w_eco116727, w_eco116728, w_eco116729, w_eco116730, w_eco116731, w_eco116732, w_eco116733, w_eco116734, w_eco116735, w_eco116736, w_eco116737, w_eco116738, w_eco116739, w_eco116740, w_eco116741, w_eco116742, w_eco116743, w_eco116744, w_eco116745, w_eco116746, w_eco116747, w_eco116748, w_eco116749, w_eco116750, w_eco116751, w_eco116752, w_eco116753, w_eco116754, w_eco116755, w_eco116756, w_eco116757, w_eco116758, w_eco116759, w_eco116760, w_eco116761, w_eco116762, w_eco116763, w_eco116764, w_eco116765, w_eco116766, w_eco116767, w_eco116768, w_eco116769, w_eco116770, w_eco116771, w_eco116772, w_eco116773, w_eco116774, w_eco116775, w_eco116776, w_eco116777, w_eco116778, w_eco116779, w_eco116780, w_eco116781, w_eco116782, w_eco116783, w_eco116784, w_eco116785, w_eco116786, w_eco116787, w_eco116788, w_eco116789, w_eco116790, w_eco116791, w_eco116792, w_eco116793, w_eco116794, w_eco116795, w_eco116796, w_eco116797, w_eco116798, w_eco116799, w_eco116800, w_eco116801, w_eco116802, w_eco116803, w_eco116804, w_eco116805, w_eco116806, w_eco116807, w_eco116808, w_eco116809, w_eco116810, w_eco116811, w_eco116812, w_eco116813, w_eco116814, w_eco116815, w_eco116816, w_eco116817, w_eco116818, w_eco116819, w_eco116820, w_eco116821, w_eco116822, w_eco116823, w_eco116824, w_eco116825, w_eco116826, w_eco116827, w_eco116828, w_eco116829, w_eco116830, w_eco116831, w_eco116832, w_eco116833, w_eco116834, w_eco116835, w_eco116836, w_eco116837, w_eco116838, w_eco116839, w_eco116840, w_eco116841, w_eco116842, w_eco116843, w_eco116844, w_eco116845, w_eco116846, w_eco116847, w_eco116848, w_eco116849, w_eco116850, w_eco116851, w_eco116852, w_eco116853, w_eco116854, w_eco116855, w_eco116856, w_eco116857, w_eco116858, w_eco116859, w_eco116860, w_eco116861, w_eco116862, w_eco116863, w_eco116864, w_eco116865, w_eco116866, w_eco116867, w_eco116868, w_eco116869, w_eco116870, w_eco116871, w_eco116872, w_eco116873, w_eco116874, w_eco116875, w_eco116876, w_eco116877, w_eco116878, w_eco116879, w_eco116880, w_eco116881, w_eco116882, w_eco116883, w_eco116884, w_eco116885, w_eco116886, w_eco116887, w_eco116888, w_eco116889, w_eco116890, w_eco116891, w_eco116892, w_eco116893, w_eco116894, w_eco116895, w_eco116896, w_eco116897, w_eco116898, w_eco116899, w_eco116900, w_eco116901, w_eco116902, w_eco116903, w_eco116904, w_eco116905, w_eco116906, w_eco116907, w_eco116908, w_eco116909, w_eco116910, w_eco116911, w_eco116912, w_eco116913, w_eco116914, w_eco116915, w_eco116916, w_eco116917, w_eco116918, w_eco116919, w_eco116920, w_eco116921, w_eco116922, w_eco116923, w_eco116924, w_eco116925, w_eco116926, w_eco116927, w_eco116928, w_eco116929, w_eco116930, w_eco116931, w_eco116932, w_eco116933, w_eco116934, w_eco116935, w_eco116936, w_eco116937, w_eco116938, w_eco116939, w_eco116940, w_eco116941, w_eco116942, w_eco116943, w_eco116944, w_eco116945, w_eco116946, w_eco116947, w_eco116948, w_eco116949, w_eco116950, w_eco116951, w_eco116952, w_eco116953, w_eco116954, w_eco116955, w_eco116956, w_eco116957, w_eco116958, w_eco116959, w_eco116960, w_eco116961, w_eco116962, w_eco116963, w_eco116964, w_eco116965, w_eco116966, w_eco116967, w_eco116968, w_eco116969, w_eco116970, w_eco116971, w_eco116972, w_eco116973, w_eco116974, w_eco116975, w_eco116976, w_eco116977, w_eco116978, w_eco116979, w_eco116980, w_eco116981, w_eco116982, w_eco116983, w_eco116984, w_eco116985, w_eco116986, w_eco116987, w_eco116988, w_eco116989, w_eco116990, w_eco116991, w_eco116992, w_eco116993, w_eco116994, w_eco116995, w_eco116996, w_eco116997, w_eco116998, w_eco116999, w_eco117000, w_eco117001, w_eco117002, w_eco117003, w_eco117004, w_eco117005, w_eco117006, w_eco117007, w_eco117008, w_eco117009, w_eco117010, w_eco117011, w_eco117012, w_eco117013, w_eco117014, w_eco117015, w_eco117016, w_eco117017, w_eco117018, w_eco117019, w_eco117020, w_eco117021, w_eco117022, w_eco117023, w_eco117024, w_eco117025, w_eco117026, w_eco117027, w_eco117028, w_eco117029, w_eco117030, w_eco117031, w_eco117032, w_eco117033, w_eco117034, w_eco117035, w_eco117036, w_eco117037, w_eco117038, w_eco117039, w_eco117040, w_eco117041, w_eco117042, w_eco117043, w_eco117044, w_eco117045, w_eco117046, w_eco117047, w_eco117048, w_eco117049, w_eco117050, w_eco117051, w_eco117052, w_eco117053, w_eco117054, w_eco117055, w_eco117056, w_eco117057, w_eco117058, w_eco117059, w_eco117060, w_eco117061, w_eco117062, w_eco117063, w_eco117064, w_eco117065, w_eco117066, w_eco117067, w_eco117068, w_eco117069, w_eco117070, w_eco117071, w_eco117072, w_eco117073, w_eco117074, w_eco117075, w_eco117076, w_eco117077, w_eco117078, w_eco117079, w_eco117080, w_eco117081, w_eco117082, w_eco117083, w_eco117084, w_eco117085, w_eco117086, w_eco117087, w_eco117088, w_eco117089, w_eco117090, w_eco117091, w_eco117092, w_eco117093, w_eco117094, w_eco117095, w_eco117096, w_eco117097, w_eco117098, w_eco117099, w_eco117100, w_eco117101, w_eco117102, w_eco117103, w_eco117104, w_eco117105, w_eco117106, w_eco117107, w_eco117108, w_eco117109, w_eco117110, w_eco117111, w_eco117112, w_eco117113, w_eco117114, w_eco117115, w_eco117116, w_eco117117, w_eco117118, w_eco117119, w_eco117120, w_eco117121, w_eco117122, w_eco117123, w_eco117124, w_eco117125, w_eco117126, w_eco117127, w_eco117128, w_eco117129, w_eco117130, w_eco117131, w_eco117132, w_eco117133, w_eco117134, w_eco117135, w_eco117136, w_eco117137, w_eco117138, w_eco117139, w_eco117140, w_eco117141, w_eco117142, w_eco117143, w_eco117144, w_eco117145, w_eco117146, w_eco117147, w_eco117148, w_eco117149, w_eco117150, w_eco117151, w_eco117152, w_eco117153, w_eco117154, w_eco117155, w_eco117156, w_eco117157, w_eco117158, w_eco117159, w_eco117160, w_eco117161, w_eco117162, w_eco117163, w_eco117164, w_eco117165, w_eco117166, w_eco117167, w_eco117168, w_eco117169, w_eco117170, w_eco117171, w_eco117172, w_eco117173, w_eco117174, w_eco117175, w_eco117176, w_eco117177, w_eco117178, w_eco117179, w_eco117180, w_eco117181, w_eco117182, w_eco117183, w_eco117184, w_eco117185, w_eco117186, w_eco117187, w_eco117188, w_eco117189, w_eco117190, w_eco117191, w_eco117192, w_eco117193, w_eco117194, w_eco117195, w_eco117196, w_eco117197, w_eco117198, w_eco117199, w_eco117200, w_eco117201, w_eco117202, w_eco117203, w_eco117204, w_eco117205, w_eco117206, w_eco117207, w_eco117208, w_eco117209, w_eco117210, w_eco117211, w_eco117212, w_eco117213, w_eco117214, w_eco117215, w_eco117216, w_eco117217, w_eco117218, w_eco117219, w_eco117220, w_eco117221, w_eco117222, w_eco117223, w_eco117224, w_eco117225, w_eco117226, w_eco117227, w_eco117228, w_eco117229, w_eco117230, w_eco117231, w_eco117232, w_eco117233, w_eco117234, w_eco117235, w_eco117236, w_eco117237, w_eco117238, w_eco117239, w_eco117240, w_eco117241, w_eco117242, w_eco117243, w_eco117244, w_eco117245, w_eco117246, w_eco117247, w_eco117248, w_eco117249, w_eco117250, w_eco117251, w_eco117252, w_eco117253, w_eco117254, w_eco117255, w_eco117256, w_eco117257, w_eco117258, w_eco117259, w_eco117260, w_eco117261, w_eco117262, w_eco117263, w_eco117264, w_eco117265, w_eco117266, w_eco117267, w_eco117268, w_eco117269, w_eco117270, w_eco117271, w_eco117272, w_eco117273, w_eco117274, w_eco117275, w_eco117276, w_eco117277, w_eco117278, w_eco117279, w_eco117280, w_eco117281, w_eco117282, w_eco117283, w_eco117284, w_eco117285, w_eco117286, w_eco117287, w_eco117288, w_eco117289, w_eco117290, w_eco117291, w_eco117292, w_eco117293, w_eco117294, w_eco117295, w_eco117296, w_eco117297, w_eco117298, w_eco117299, w_eco117300, w_eco117301, w_eco117302, w_eco117303, w_eco117304, w_eco117305, w_eco117306, w_eco117307, w_eco117308, w_eco117309, w_eco117310, w_eco117311, w_eco117312, w_eco117313, w_eco117314, w_eco117315, w_eco117316, w_eco117317, w_eco117318, w_eco117319, w_eco117320, w_eco117321, w_eco117322, w_eco117323, w_eco117324, w_eco117325, w_eco117326, w_eco117327, w_eco117328, w_eco117329, w_eco117330, w_eco117331, w_eco117332, w_eco117333, w_eco117334, w_eco117335, w_eco117336, w_eco117337, w_eco117338, w_eco117339, w_eco117340, w_eco117341, w_eco117342, w_eco117343, w_eco117344, w_eco117345, w_eco117346, w_eco117347, w_eco117348, w_eco117349, w_eco117350, w_eco117351, w_eco117352, w_eco117353, w_eco117354, w_eco117355, w_eco117356, w_eco117357, w_eco117358, w_eco117359, w_eco117360, w_eco117361, w_eco117362, w_eco117363, w_eco117364, w_eco117365, w_eco117366, w_eco117367, w_eco117368, w_eco117369, w_eco117370, w_eco117371, w_eco117372, w_eco117373, w_eco117374, w_eco117375, w_eco117376, w_eco117377, w_eco117378, w_eco117379, w_eco117380, w_eco117381, w_eco117382, w_eco117383, w_eco117384, w_eco117385, w_eco117386, w_eco117387, w_eco117388, w_eco117389, w_eco117390, w_eco117391, w_eco117392, w_eco117393, w_eco117394, w_eco117395, w_eco117396, w_eco117397, w_eco117398, w_eco117399, w_eco117400, w_eco117401, w_eco117402, w_eco117403, w_eco117404, w_eco117405, w_eco117406, w_eco117407, w_eco117408, w_eco117409, w_eco117410, w_eco117411, w_eco117412, w_eco117413, w_eco117414, w_eco117415, w_eco117416, w_eco117417, w_eco117418, w_eco117419, w_eco117420, w_eco117421, w_eco117422, w_eco117423, w_eco117424, w_eco117425, w_eco117426, w_eco117427, w_eco117428, w_eco117429, w_eco117430, w_eco117431, w_eco117432, w_eco117433, w_eco117434, w_eco117435, w_eco117436, w_eco117437, w_eco117438, w_eco117439, w_eco117440, w_eco117441, w_eco117442, w_eco117443, w_eco117444, w_eco117445, w_eco117446, w_eco117447, w_eco117448, w_eco117449, w_eco117450, w_eco117451, w_eco117452, w_eco117453, w_eco117454, w_eco117455, w_eco117456, w_eco117457, w_eco117458, w_eco117459, w_eco117460, w_eco117461, w_eco117462, w_eco117463, w_eco117464, w_eco117465, w_eco117466, w_eco117467, w_eco117468, w_eco117469, w_eco117470, w_eco117471, w_eco117472, w_eco117473, w_eco117474, w_eco117475, w_eco117476, w_eco117477, w_eco117478, w_eco117479, w_eco117480, w_eco117481, w_eco117482, w_eco117483, w_eco117484, w_eco117485, w_eco117486, w_eco117487, w_eco117488, w_eco117489, w_eco117490, w_eco117491, w_eco117492, w_eco117493, w_eco117494, w_eco117495, w_eco117496, w_eco117497, w_eco117498, w_eco117499, w_eco117500, w_eco117501, w_eco117502, w_eco117503, w_eco117504, w_eco117505, w_eco117506, w_eco117507, w_eco117508, w_eco117509, w_eco117510, w_eco117511, w_eco117512, w_eco117513, w_eco117514, w_eco117515, w_eco117516, w_eco117517, w_eco117518, w_eco117519, w_eco117520, w_eco117521, w_eco117522, w_eco117523, w_eco117524, w_eco117525, w_eco117526, w_eco117527, w_eco117528, w_eco117529, w_eco117530, w_eco117531, w_eco117532, w_eco117533, w_eco117534, w_eco117535, w_eco117536, w_eco117537, w_eco117538, w_eco117539, w_eco117540, w_eco117541, w_eco117542, w_eco117543, w_eco117544, w_eco117545, w_eco117546, w_eco117547, w_eco117548, w_eco117549, w_eco117550, w_eco117551, w_eco117552, w_eco117553, w_eco117554, w_eco117555, w_eco117556, w_eco117557, w_eco117558, w_eco117559, w_eco117560, w_eco117561, w_eco117562, w_eco117563, w_eco117564, w_eco117565, w_eco117566, w_eco117567, w_eco117568, w_eco117569, w_eco117570, w_eco117571, w_eco117572, w_eco117573, w_eco117574, w_eco117575, w_eco117576, w_eco117577, w_eco117578, w_eco117579, w_eco117580, w_eco117581, w_eco117582, w_eco117583, w_eco117584, w_eco117585, w_eco117586, w_eco117587, w_eco117588, w_eco117589, w_eco117590, w_eco117591, w_eco117592, w_eco117593, w_eco117594, w_eco117595, w_eco117596, w_eco117597, w_eco117598, w_eco117599, w_eco117600, w_eco117601, w_eco117602, w_eco117603, w_eco117604, w_eco117605, w_eco117606, w_eco117607, w_eco117608, w_eco117609, w_eco117610, w_eco117611, w_eco117612, w_eco117613, w_eco117614, w_eco117615, w_eco117616, w_eco117617, w_eco117618, w_eco117619, w_eco117620, w_eco117621, w_eco117622, w_eco117623, w_eco117624, w_eco117625, w_eco117626, w_eco117627, w_eco117628, w_eco117629, w_eco117630, w_eco117631, w_eco117632, w_eco117633, w_eco117634, w_eco117635, w_eco117636, w_eco117637, w_eco117638, w_eco117639, w_eco117640, w_eco117641, w_eco117642, w_eco117643, w_eco117644, w_eco117645, w_eco117646, w_eco117647, w_eco117648, w_eco117649, w_eco117650, w_eco117651, w_eco117652, w_eco117653, w_eco117654, w_eco117655, w_eco117656, w_eco117657, w_eco117658, w_eco117659, w_eco117660, w_eco117661, w_eco117662, w_eco117663, w_eco117664, w_eco117665, w_eco117666, w_eco117667, w_eco117668, w_eco117669, w_eco117670, w_eco117671, w_eco117672, w_eco117673, w_eco117674, w_eco117675, w_eco117676, w_eco117677, w_eco117678, w_eco117679, w_eco117680, w_eco117681, w_eco117682, w_eco117683, w_eco117684, w_eco117685, w_eco117686, w_eco117687, w_eco117688, w_eco117689, w_eco117690, w_eco117691, w_eco117692, w_eco117693, w_eco117694, w_eco117695, w_eco117696, w_eco117697, w_eco117698, w_eco117699, w_eco117700, w_eco117701, w_eco117702, w_eco117703, w_eco117704, w_eco117705, w_eco117706, w_eco117707, w_eco117708, w_eco117709, w_eco117710, w_eco117711, w_eco117712, w_eco117713, w_eco117714, w_eco117715, w_eco117716, w_eco117717, w_eco117718, w_eco117719, w_eco117720, w_eco117721, w_eco117722, w_eco117723, w_eco117724, w_eco117725, w_eco117726, w_eco117727, w_eco117728, w_eco117729, w_eco117730, w_eco117731, w_eco117732, w_eco117733, w_eco117734, w_eco117735, w_eco117736, w_eco117737, w_eco117738, w_eco117739, w_eco117740, w_eco117741, w_eco117742, w_eco117743, w_eco117744, w_eco117745, w_eco117746, w_eco117747, w_eco117748, w_eco117749, w_eco117750, w_eco117751, w_eco117752, w_eco117753, w_eco117754, w_eco117755, w_eco117756, w_eco117757, w_eco117758, w_eco117759, w_eco117760, w_eco117761, w_eco117762, w_eco117763, w_eco117764, w_eco117765, w_eco117766, w_eco117767, w_eco117768, w_eco117769, w_eco117770, w_eco117771, w_eco117772, w_eco117773, w_eco117774, w_eco117775, w_eco117776, w_eco117777, w_eco117778, w_eco117779, w_eco117780, w_eco117781, w_eco117782, w_eco117783, w_eco117784, w_eco117785, w_eco117786, w_eco117787, w_eco117788, w_eco117789, w_eco117790, w_eco117791, w_eco117792, w_eco117793, w_eco117794, w_eco117795, w_eco117796, w_eco117797, w_eco117798, w_eco117799, w_eco117800, w_eco117801, w_eco117802, w_eco117803, w_eco117804, w_eco117805, w_eco117806, w_eco117807, w_eco117808, w_eco117809, w_eco117810, w_eco117811, w_eco117812, w_eco117813, w_eco117814, w_eco117815, w_eco117816, w_eco117817, w_eco117818, w_eco117819, w_eco117820, w_eco117821, w_eco117822, w_eco117823, w_eco117824, w_eco117825, w_eco117826, w_eco117827, w_eco117828, w_eco117829, w_eco117830, w_eco117831, w_eco117832, w_eco117833, w_eco117834, w_eco117835, w_eco117836, w_eco117837, w_eco117838, w_eco117839, w_eco117840, w_eco117841, w_eco117842, w_eco117843, w_eco117844, w_eco117845, w_eco117846, w_eco117847, w_eco117848, w_eco117849, w_eco117850, w_eco117851, w_eco117852, w_eco117853, w_eco117854, w_eco117855, w_eco117856, w_eco117857, w_eco117858, w_eco117859, w_eco117860, w_eco117861, w_eco117862, w_eco117863, w_eco117864, w_eco117865, w_eco117866, w_eco117867, w_eco117868, w_eco117869, w_eco117870, w_eco117871, w_eco117872, w_eco117873, w_eco117874, w_eco117875, w_eco117876, w_eco117877, w_eco117878, w_eco117879, w_eco117880, w_eco117881, w_eco117882, w_eco117883, w_eco117884, w_eco117885, w_eco117886, w_eco117887, w_eco117888, w_eco117889, w_eco117890, w_eco117891, w_eco117892, w_eco117893, w_eco117894, w_eco117895, w_eco117896, w_eco117897, w_eco117898, w_eco117899, w_eco117900, w_eco117901, w_eco117902, w_eco117903, w_eco117904, w_eco117905, w_eco117906, w_eco117907, w_eco117908, w_eco117909, w_eco117910, w_eco117911, w_eco117912, w_eco117913, w_eco117914, w_eco117915, w_eco117916, w_eco117917, w_eco117918, w_eco117919, w_eco117920, w_eco117921, w_eco117922, w_eco117923, w_eco117924, w_eco117925, w_eco117926, w_eco117927, w_eco117928, w_eco117929, w_eco117930, w_eco117931, w_eco117932, w_eco117933, w_eco117934, w_eco117935, w_eco117936, w_eco117937, w_eco117938, w_eco117939, w_eco117940, w_eco117941, w_eco117942, w_eco117943, w_eco117944, w_eco117945, w_eco117946, w_eco117947, w_eco117948, w_eco117949, w_eco117950, w_eco117951, w_eco117952, w_eco117953, w_eco117954, w_eco117955, w_eco117956, w_eco117957, w_eco117958, w_eco117959, w_eco117960, w_eco117961, w_eco117962, w_eco117963, w_eco117964, w_eco117965, w_eco117966, w_eco117967, w_eco117968, w_eco117969, w_eco117970, w_eco117971, w_eco117972, w_eco117973, w_eco117974, w_eco117975, w_eco117976, w_eco117977, w_eco117978, w_eco117979, w_eco117980, w_eco117981, w_eco117982, w_eco117983, w_eco117984, w_eco117985, w_eco117986, w_eco117987, w_eco117988, w_eco117989, w_eco117990, w_eco117991, w_eco117992, w_eco117993, w_eco117994, w_eco117995, w_eco117996, w_eco117997, w_eco117998, w_eco117999, w_eco118000, w_eco118001, w_eco118002, w_eco118003, w_eco118004, w_eco118005, w_eco118006, w_eco118007, w_eco118008, w_eco118009, w_eco118010, w_eco118011, w_eco118012, w_eco118013, w_eco118014, w_eco118015, w_eco118016, w_eco118017, w_eco118018, w_eco118019, w_eco118020, w_eco118021, w_eco118022, w_eco118023, w_eco118024, w_eco118025, w_eco118026, w_eco118027, w_eco118028, w_eco118029, w_eco118030, w_eco118031, w_eco118032, w_eco118033, w_eco118034, w_eco118035, w_eco118036, w_eco118037, w_eco118038, w_eco118039, w_eco118040, w_eco118041, w_eco118042, w_eco118043, w_eco118044, w_eco118045, w_eco118046, w_eco118047, w_eco118048, w_eco118049, w_eco118050, w_eco118051, w_eco118052, w_eco118053, w_eco118054, w_eco118055, w_eco118056, w_eco118057, w_eco118058, w_eco118059, w_eco118060, w_eco118061, w_eco118062, w_eco118063, w_eco118064, w_eco118065, w_eco118066, w_eco118067, w_eco118068, w_eco118069, w_eco118070, w_eco118071, w_eco118072, w_eco118073, w_eco118074, w_eco118075, w_eco118076, w_eco118077, w_eco118078, w_eco118079, w_eco118080, w_eco118081, w_eco118082, w_eco118083, w_eco118084, w_eco118085, w_eco118086, w_eco118087, w_eco118088, w_eco118089, w_eco118090, w_eco118091, w_eco118092, w_eco118093, w_eco118094, w_eco118095, w_eco118096, w_eco118097, w_eco118098, w_eco118099, w_eco118100, w_eco118101, w_eco118102, w_eco118103, w_eco118104, w_eco118105, w_eco118106, w_eco118107, w_eco118108, w_eco118109, w_eco118110, w_eco118111, w_eco118112, w_eco118113, w_eco118114, w_eco118115, w_eco118116, w_eco118117, w_eco118118, w_eco118119, w_eco118120, w_eco118121, w_eco118122, w_eco118123, w_eco118124, w_eco118125, w_eco118126, w_eco118127, w_eco118128, w_eco118129, w_eco118130, w_eco118131, w_eco118132, w_eco118133, w_eco118134, w_eco118135, w_eco118136, w_eco118137, w_eco118138, w_eco118139, w_eco118140, w_eco118141, w_eco118142, w_eco118143, w_eco118144, w_eco118145, w_eco118146, w_eco118147, w_eco118148, w_eco118149, w_eco118150, w_eco118151, w_eco118152, w_eco118153, w_eco118154, w_eco118155, w_eco118156, w_eco118157, w_eco118158, w_eco118159, w_eco118160, w_eco118161, w_eco118162, w_eco118163, w_eco118164, w_eco118165, w_eco118166, w_eco118167, w_eco118168, w_eco118169, w_eco118170, w_eco118171, w_eco118172, w_eco118173, w_eco118174, w_eco118175, w_eco118176, w_eco118177, w_eco118178, w_eco118179, w_eco118180, w_eco118181, w_eco118182, w_eco118183, w_eco118184, w_eco118185, w_eco118186, w_eco118187, w_eco118188, w_eco118189, w_eco118190, w_eco118191, w_eco118192, w_eco118193, w_eco118194, w_eco118195, w_eco118196, w_eco118197, w_eco118198, w_eco118199, w_eco118200, w_eco118201, w_eco118202, w_eco118203, w_eco118204, w_eco118205, w_eco118206, w_eco118207, w_eco118208, w_eco118209, w_eco118210, w_eco118211, w_eco118212, w_eco118213, w_eco118214, w_eco118215, w_eco118216, w_eco118217, w_eco118218, w_eco118219, w_eco118220, w_eco118221, w_eco118222, w_eco118223, w_eco118224, w_eco118225, w_eco118226, w_eco118227, w_eco118228, w_eco118229, w_eco118230, w_eco118231, w_eco118232, w_eco118233, w_eco118234, w_eco118235, w_eco118236, w_eco118237, w_eco118238, w_eco118239, w_eco118240, w_eco118241, w_eco118242, w_eco118243, w_eco118244, w_eco118245, w_eco118246, w_eco118247, w_eco118248, w_eco118249, w_eco118250, w_eco118251, w_eco118252, w_eco118253, w_eco118254, w_eco118255, w_eco118256, w_eco118257, w_eco118258, w_eco118259, w_eco118260, w_eco118261, w_eco118262, w_eco118263, w_eco118264, w_eco118265, w_eco118266, w_eco118267, w_eco118268, w_eco118269, w_eco118270, w_eco118271, w_eco118272, w_eco118273, w_eco118274, w_eco118275, w_eco118276, w_eco118277, w_eco118278, w_eco118279, w_eco118280, w_eco118281, w_eco118282, w_eco118283, w_eco118284, w_eco118285, w_eco118286, w_eco118287, w_eco118288, w_eco118289, w_eco118290, w_eco118291, w_eco118292, w_eco118293, w_eco118294, w_eco118295, w_eco118296, w_eco118297, w_eco118298, w_eco118299, w_eco118300, w_eco118301, w_eco118302, w_eco118303, w_eco118304, w_eco118305, w_eco118306, w_eco118307, w_eco118308, w_eco118309, w_eco118310, w_eco118311, w_eco118312, w_eco118313, w_eco118314, w_eco118315, w_eco118316, w_eco118317, w_eco118318, w_eco118319, w_eco118320, w_eco118321, w_eco118322, w_eco118323, w_eco118324, w_eco118325, w_eco118326, w_eco118327, w_eco118328, w_eco118329, w_eco118330, w_eco118331, w_eco118332, w_eco118333, w_eco118334, w_eco118335, w_eco118336, w_eco118337, w_eco118338, w_eco118339, w_eco118340, w_eco118341, w_eco118342, w_eco118343, w_eco118344, w_eco118345, w_eco118346, w_eco118347, w_eco118348, w_eco118349, w_eco118350, w_eco118351, w_eco118352, w_eco118353, w_eco118354, w_eco118355, w_eco118356, w_eco118357, w_eco118358, w_eco118359, w_eco118360, w_eco118361, w_eco118362, w_eco118363, w_eco118364, w_eco118365, w_eco118366, w_eco118367, w_eco118368, w_eco118369, w_eco118370, w_eco118371, w_eco118372, w_eco118373, w_eco118374, w_eco118375, w_eco118376, w_eco118377, w_eco118378, w_eco118379, w_eco118380, w_eco118381, w_eco118382, w_eco118383, w_eco118384, w_eco118385, w_eco118386, w_eco118387, w_eco118388, w_eco118389, w_eco118390, w_eco118391, w_eco118392, w_eco118393, w_eco118394, w_eco118395, w_eco118396, w_eco118397, w_eco118398, w_eco118399, w_eco118400, w_eco118401, w_eco118402, w_eco118403, w_eco118404, w_eco118405, w_eco118406, w_eco118407, w_eco118408, w_eco118409, w_eco118410, w_eco118411, w_eco118412, w_eco118413, w_eco118414, w_eco118415, w_eco118416, w_eco118417, w_eco118418, w_eco118419, w_eco118420, w_eco118421, w_eco118422, w_eco118423, w_eco118424, w_eco118425, w_eco118426, w_eco118427, w_eco118428, w_eco118429, w_eco118430, w_eco118431, w_eco118432, w_eco118433, w_eco118434, w_eco118435, w_eco118436, w_eco118437, w_eco118438, w_eco118439, w_eco118440, w_eco118441, w_eco118442, w_eco118443, w_eco118444, w_eco118445, w_eco118446, w_eco118447, w_eco118448, w_eco118449, w_eco118450, w_eco118451, w_eco118452, w_eco118453, w_eco118454, w_eco118455, w_eco118456, w_eco118457, w_eco118458, w_eco118459, w_eco118460, w_eco118461, w_eco118462, w_eco118463, w_eco118464, w_eco118465, w_eco118466, w_eco118467, w_eco118468, w_eco118469, w_eco118470, w_eco118471, w_eco118472, w_eco118473, w_eco118474, w_eco118475, w_eco118476, w_eco118477, w_eco118478, w_eco118479, w_eco118480, w_eco118481, w_eco118482, w_eco118483, w_eco118484, w_eco118485, w_eco118486, w_eco118487, w_eco118488, w_eco118489, w_eco118490, w_eco118491, w_eco118492, w_eco118493, w_eco118494, w_eco118495, w_eco118496, w_eco118497, w_eco118498, w_eco118499, w_eco118500, w_eco118501, w_eco118502, w_eco118503, w_eco118504, w_eco118505, w_eco118506, w_eco118507, w_eco118508, w_eco118509, w_eco118510, w_eco118511, w_eco118512, w_eco118513, w_eco118514, w_eco118515, w_eco118516, w_eco118517, w_eco118518, w_eco118519, w_eco118520, w_eco118521, w_eco118522, w_eco118523, w_eco118524, w_eco118525, w_eco118526, w_eco118527, w_eco118528, w_eco118529, w_eco118530, w_eco118531, w_eco118532, w_eco118533, w_eco118534, w_eco118535, w_eco118536, w_eco118537, w_eco118538, w_eco118539, w_eco118540, w_eco118541, w_eco118542, w_eco118543, w_eco118544, w_eco118545, w_eco118546, w_eco118547, w_eco118548, w_eco118549, w_eco118550, w_eco118551, w_eco118552, w_eco118553, w_eco118554, w_eco118555, w_eco118556, w_eco118557, w_eco118558, w_eco118559, w_eco118560, w_eco118561, w_eco118562, w_eco118563, w_eco118564, w_eco118565, w_eco118566, w_eco118567, w_eco118568, w_eco118569, w_eco118570, w_eco118571, w_eco118572, w_eco118573, w_eco118574, w_eco118575, w_eco118576, w_eco118577, w_eco118578, w_eco118579, w_eco118580, w_eco118581, w_eco118582, w_eco118583, w_eco118584, w_eco118585, w_eco118586, w_eco118587, w_eco118588, w_eco118589, w_eco118590, w_eco118591, w_eco118592, w_eco118593, w_eco118594, w_eco118595, w_eco118596, w_eco118597, w_eco118598, w_eco118599, w_eco118600, w_eco118601, w_eco118602, w_eco118603, w_eco118604, w_eco118605, w_eco118606, w_eco118607, w_eco118608, w_eco118609, w_eco118610, w_eco118611, w_eco118612, w_eco118613, w_eco118614, w_eco118615, w_eco118616, w_eco118617, w_eco118618, w_eco118619, w_eco118620, w_eco118621, w_eco118622, w_eco118623, w_eco118624, w_eco118625, w_eco118626, w_eco118627, w_eco118628, w_eco118629, w_eco118630, w_eco118631, w_eco118632, w_eco118633, w_eco118634, w_eco118635, w_eco118636, w_eco118637, w_eco118638, w_eco118639, w_eco118640, w_eco118641, w_eco118642, w_eco118643, w_eco118644, w_eco118645, w_eco118646, w_eco118647, w_eco118648, w_eco118649, w_eco118650, w_eco118651, w_eco118652, w_eco118653, w_eco118654, w_eco118655, w_eco118656, w_eco118657, w_eco118658, w_eco118659, w_eco118660, w_eco118661, w_eco118662, w_eco118663, w_eco118664, w_eco118665, w_eco118666, w_eco118667, w_eco118668, w_eco118669, w_eco118670, w_eco118671, w_eco118672, w_eco118673, w_eco118674, w_eco118675, w_eco118676, w_eco118677, w_eco118678, w_eco118679, w_eco118680, w_eco118681, w_eco118682, w_eco118683, w_eco118684, w_eco118685, w_eco118686, w_eco118687, w_eco118688, w_eco118689, w_eco118690, w_eco118691, w_eco118692, w_eco118693, w_eco118694, w_eco118695, w_eco118696, w_eco118697, w_eco118698, w_eco118699, w_eco118700, w_eco118701, w_eco118702, w_eco118703, w_eco118704, w_eco118705, w_eco118706, w_eco118707, w_eco118708, w_eco118709, w_eco118710, w_eco118711, w_eco118712, w_eco118713, w_eco118714, w_eco118715, w_eco118716, w_eco118717, w_eco118718, w_eco118719, w_eco118720, w_eco118721, w_eco118722, w_eco118723, w_eco118724, w_eco118725, w_eco118726, w_eco118727, w_eco118728, w_eco118729, w_eco118730, w_eco118731, w_eco118732, w_eco118733, w_eco118734, w_eco118735, w_eco118736, w_eco118737, w_eco118738, w_eco118739, w_eco118740, w_eco118741, w_eco118742, w_eco118743, w_eco118744, w_eco118745, w_eco118746, w_eco118747, w_eco118748, w_eco118749, w_eco118750, w_eco118751, w_eco118752, w_eco118753, w_eco118754, w_eco118755, w_eco118756, w_eco118757, w_eco118758, w_eco118759, w_eco118760, w_eco118761, w_eco118762, w_eco118763, w_eco118764, w_eco118765, w_eco118766, w_eco118767, w_eco118768, w_eco118769, w_eco118770, w_eco118771, w_eco118772, w_eco118773, w_eco118774, w_eco118775, w_eco118776, w_eco118777, w_eco118778, w_eco118779, w_eco118780, w_eco118781, w_eco118782, w_eco118783, w_eco118784, w_eco118785, w_eco118786, w_eco118787, w_eco118788, w_eco118789, w_eco118790, w_eco118791, w_eco118792, w_eco118793, w_eco118794, w_eco118795, w_eco118796, w_eco118797, w_eco118798, w_eco118799, w_eco118800, w_eco118801, w_eco118802, w_eco118803, w_eco118804, w_eco118805, w_eco118806, w_eco118807, w_eco118808, w_eco118809, w_eco118810, w_eco118811, w_eco118812, w_eco118813, w_eco118814, w_eco118815, w_eco118816, w_eco118817, w_eco118818, w_eco118819, w_eco118820, w_eco118821, w_eco118822, w_eco118823, w_eco118824, w_eco118825, w_eco118826, w_eco118827, w_eco118828, w_eco118829, w_eco118830, w_eco118831, w_eco118832, w_eco118833, w_eco118834, w_eco118835, w_eco118836, w_eco118837, w_eco118838, w_eco118839, w_eco118840, w_eco118841, w_eco118842, w_eco118843, w_eco118844, w_eco118845, w_eco118846, w_eco118847, w_eco118848, w_eco118849, w_eco118850, w_eco118851, w_eco118852, w_eco118853, w_eco118854, w_eco118855, w_eco118856, w_eco118857, w_eco118858, w_eco118859, w_eco118860, w_eco118861, w_eco118862, w_eco118863, w_eco118864, w_eco118865, w_eco118866, w_eco118867, w_eco118868, w_eco118869, w_eco118870, w_eco118871, w_eco118872, w_eco118873, w_eco118874, w_eco118875, w_eco118876, w_eco118877, w_eco118878, w_eco118879, w_eco118880, w_eco118881, w_eco118882, w_eco118883, w_eco118884, w_eco118885, w_eco118886, w_eco118887, w_eco118888, w_eco118889, w_eco118890, w_eco118891, w_eco118892, w_eco118893, w_eco118894, w_eco118895, w_eco118896, w_eco118897, w_eco118898, w_eco118899, w_eco118900, w_eco118901, w_eco118902, w_eco118903, w_eco118904, w_eco118905, w_eco118906, w_eco118907, w_eco118908, w_eco118909, w_eco118910, w_eco118911, w_eco118912, w_eco118913, w_eco118914, w_eco118915, w_eco118916, w_eco118917, w_eco118918, w_eco118919, w_eco118920, w_eco118921, w_eco118922, w_eco118923, w_eco118924, w_eco118925, w_eco118926, w_eco118927, w_eco118928, w_eco118929, w_eco118930, w_eco118931, w_eco118932, w_eco118933, w_eco118934, w_eco118935, w_eco118936, w_eco118937, w_eco118938, w_eco118939, w_eco118940, w_eco118941, w_eco118942, w_eco118943, w_eco118944, w_eco118945, w_eco118946, w_eco118947, w_eco118948, w_eco118949, w_eco118950, w_eco118951, w_eco118952, w_eco118953, w_eco118954, w_eco118955, w_eco118956, w_eco118957, w_eco118958, w_eco118959, w_eco118960, w_eco118961, w_eco118962, w_eco118963, w_eco118964, w_eco118965, w_eco118966, w_eco118967, w_eco118968, w_eco118969, w_eco118970, w_eco118971, w_eco118972, w_eco118973, w_eco118974, w_eco118975, w_eco118976, w_eco118977, w_eco118978, w_eco118979, w_eco118980, w_eco118981, w_eco118982, w_eco118983, w_eco118984, w_eco118985, w_eco118986, w_eco118987, w_eco118988, w_eco118989, w_eco118990, w_eco118991, w_eco118992, w_eco118993, w_eco118994, w_eco118995, w_eco118996, w_eco118997, w_eco118998, w_eco118999, w_eco119000, w_eco119001, w_eco119002, w_eco119003, w_eco119004, w_eco119005, w_eco119006, w_eco119007, w_eco119008, w_eco119009, w_eco119010, w_eco119011, w_eco119012, w_eco119013, w_eco119014, w_eco119015, w_eco119016, w_eco119017, w_eco119018, w_eco119019, w_eco119020, w_eco119021, w_eco119022, w_eco119023, w_eco119024, w_eco119025, w_eco119026, w_eco119027, w_eco119028, w_eco119029, w_eco119030, w_eco119031, w_eco119032, w_eco119033, w_eco119034, w_eco119035, w_eco119036, w_eco119037, w_eco119038, w_eco119039, w_eco119040, w_eco119041, w_eco119042, w_eco119043, w_eco119044, w_eco119045, w_eco119046, w_eco119047, w_eco119048, w_eco119049, w_eco119050, w_eco119051, w_eco119052, w_eco119053, w_eco119054, w_eco119055, w_eco119056, w_eco119057, w_eco119058, w_eco119059, w_eco119060, w_eco119061, w_eco119062, w_eco119063, w_eco119064, w_eco119065, w_eco119066, w_eco119067, w_eco119068, w_eco119069, w_eco119070, w_eco119071, w_eco119072, w_eco119073, w_eco119074, w_eco119075, w_eco119076, w_eco119077, w_eco119078, w_eco119079, w_eco119080, w_eco119081, w_eco119082, w_eco119083, w_eco119084, w_eco119085, w_eco119086, w_eco119087, w_eco119088, w_eco119089, w_eco119090, w_eco119091, w_eco119092, w_eco119093, w_eco119094, w_eco119095, w_eco119096, w_eco119097, w_eco119098, w_eco119099, w_eco119100, w_eco119101, w_eco119102, w_eco119103, w_eco119104, w_eco119105, w_eco119106, w_eco119107, w_eco119108, w_eco119109, w_eco119110, w_eco119111, w_eco119112, w_eco119113, w_eco119114, w_eco119115, w_eco119116, w_eco119117, w_eco119118, w_eco119119, w_eco119120, w_eco119121, w_eco119122, w_eco119123, w_eco119124, w_eco119125, w_eco119126, w_eco119127, w_eco119128, w_eco119129, w_eco119130, w_eco119131, w_eco119132, w_eco119133, w_eco119134, w_eco119135, w_eco119136, w_eco119137, w_eco119138, w_eco119139, w_eco119140, w_eco119141, w_eco119142, w_eco119143, w_eco119144, w_eco119145, w_eco119146, w_eco119147, w_eco119148, w_eco119149, w_eco119150, w_eco119151, w_eco119152, w_eco119153, w_eco119154, w_eco119155, w_eco119156, w_eco119157, w_eco119158, w_eco119159, w_eco119160, w_eco119161, w_eco119162, w_eco119163, w_eco119164, w_eco119165, w_eco119166, w_eco119167, w_eco119168, w_eco119169, w_eco119170, w_eco119171, w_eco119172, w_eco119173, w_eco119174, w_eco119175, w_eco119176, w_eco119177, w_eco119178, w_eco119179, w_eco119180, w_eco119181, w_eco119182, w_eco119183, w_eco119184, w_eco119185, w_eco119186, w_eco119187, w_eco119188, w_eco119189, w_eco119190, w_eco119191, w_eco119192, w_eco119193, w_eco119194, w_eco119195, w_eco119196, w_eco119197, w_eco119198, w_eco119199, w_eco119200, w_eco119201, w_eco119202, w_eco119203, w_eco119204, w_eco119205, w_eco119206, w_eco119207, w_eco119208, w_eco119209, w_eco119210, w_eco119211, w_eco119212, w_eco119213, w_eco119214, w_eco119215, w_eco119216, w_eco119217, w_eco119218, w_eco119219, w_eco119220, w_eco119221, w_eco119222, w_eco119223, w_eco119224, w_eco119225, w_eco119226, w_eco119227, w_eco119228, w_eco119229, w_eco119230, w_eco119231, w_eco119232, w_eco119233, w_eco119234, w_eco119235, w_eco119236, w_eco119237, w_eco119238, w_eco119239, w_eco119240, w_eco119241, w_eco119242, w_eco119243, w_eco119244, w_eco119245, w_eco119246, w_eco119247, w_eco119248, w_eco119249, w_eco119250, w_eco119251, w_eco119252, w_eco119253, w_eco119254, w_eco119255, w_eco119256, w_eco119257, w_eco119258, w_eco119259, w_eco119260, w_eco119261, w_eco119262, w_eco119263, w_eco119264, w_eco119265, w_eco119266, w_eco119267, w_eco119268, w_eco119269, w_eco119270, w_eco119271, w_eco119272, w_eco119273, w_eco119274, w_eco119275, w_eco119276, w_eco119277, w_eco119278, w_eco119279, w_eco119280, w_eco119281, w_eco119282, w_eco119283, w_eco119284, w_eco119285, w_eco119286, w_eco119287, w_eco119288, w_eco119289, w_eco119290, w_eco119291, w_eco119292, w_eco119293, w_eco119294, w_eco119295, w_eco119296, w_eco119297, w_eco119298, w_eco119299, w_eco119300, w_eco119301, w_eco119302, w_eco119303, w_eco119304, w_eco119305, w_eco119306, w_eco119307, w_eco119308, w_eco119309, w_eco119310, w_eco119311, w_eco119312, w_eco119313, w_eco119314, w_eco119315, w_eco119316, w_eco119317, w_eco119318, w_eco119319, w_eco119320, w_eco119321, w_eco119322, w_eco119323, w_eco119324, w_eco119325, w_eco119326, w_eco119327, w_eco119328, w_eco119329, w_eco119330, w_eco119331, w_eco119332, w_eco119333, w_eco119334, w_eco119335, w_eco119336, w_eco119337, w_eco119338, w_eco119339, w_eco119340, w_eco119341, w_eco119342, w_eco119343, w_eco119344, w_eco119345, w_eco119346, w_eco119347, w_eco119348, w_eco119349, w_eco119350, w_eco119351, w_eco119352, w_eco119353, w_eco119354, w_eco119355, w_eco119356, w_eco119357, w_eco119358, w_eco119359, w_eco119360, w_eco119361, w_eco119362, w_eco119363, w_eco119364, w_eco119365, w_eco119366, w_eco119367, w_eco119368, w_eco119369, w_eco119370, w_eco119371, w_eco119372, w_eco119373, w_eco119374, w_eco119375, w_eco119376, w_eco119377, w_eco119378, w_eco119379, w_eco119380, w_eco119381, w_eco119382, w_eco119383, w_eco119384, w_eco119385, w_eco119386, w_eco119387, w_eco119388, w_eco119389, w_eco119390, w_eco119391, w_eco119392, w_eco119393, w_eco119394, w_eco119395, w_eco119396, w_eco119397, w_eco119398, w_eco119399, w_eco119400, w_eco119401, w_eco119402, w_eco119403, w_eco119404, w_eco119405, w_eco119406, w_eco119407, w_eco119408, w_eco119409, w_eco119410, w_eco119411, w_eco119412, w_eco119413, w_eco119414, w_eco119415, w_eco119416, w_eco119417, w_eco119418, w_eco119419, w_eco119420, w_eco119421, w_eco119422, w_eco119423, w_eco119424, w_eco119425, w_eco119426, w_eco119427, w_eco119428, w_eco119429, w_eco119430, w_eco119431, w_eco119432, w_eco119433, w_eco119434, w_eco119435, w_eco119436, w_eco119437, w_eco119438, w_eco119439, w_eco119440, w_eco119441, w_eco119442, w_eco119443, w_eco119444, w_eco119445, w_eco119446, w_eco119447, w_eco119448, w_eco119449, w_eco119450, w_eco119451, w_eco119452, w_eco119453, w_eco119454, w_eco119455, w_eco119456, w_eco119457, w_eco119458, w_eco119459, w_eco119460, w_eco119461, w_eco119462, w_eco119463, w_eco119464, w_eco119465, w_eco119466, w_eco119467, w_eco119468, w_eco119469, w_eco119470, w_eco119471, w_eco119472, w_eco119473, w_eco119474, w_eco119475, w_eco119476, w_eco119477, w_eco119478, w_eco119479, w_eco119480, w_eco119481, w_eco119482, w_eco119483, w_eco119484, w_eco119485, w_eco119486, w_eco119487, w_eco119488, w_eco119489, w_eco119490, w_eco119491, w_eco119492, w_eco119493, w_eco119494, w_eco119495, w_eco119496, w_eco119497, w_eco119498, w_eco119499, w_eco119500, w_eco119501, w_eco119502, w_eco119503, w_eco119504, w_eco119505, w_eco119506, w_eco119507, w_eco119508, w_eco119509, w_eco119510, w_eco119511, w_eco119512, w_eco119513, w_eco119514, w_eco119515, w_eco119516, w_eco119517, w_eco119518, w_eco119519, w_eco119520, w_eco119521, w_eco119522, w_eco119523, w_eco119524, w_eco119525, w_eco119526, w_eco119527, w_eco119528, w_eco119529, w_eco119530, w_eco119531, w_eco119532, w_eco119533, w_eco119534, w_eco119535, w_eco119536, w_eco119537, w_eco119538, w_eco119539, w_eco119540, w_eco119541, w_eco119542, w_eco119543, w_eco119544, w_eco119545, w_eco119546, w_eco119547, w_eco119548, w_eco119549, w_eco119550, w_eco119551, w_eco119552, w_eco119553, w_eco119554, w_eco119555, w_eco119556, w_eco119557, w_eco119558, w_eco119559, w_eco119560, w_eco119561, w_eco119562, w_eco119563, w_eco119564, w_eco119565, w_eco119566, w_eco119567, w_eco119568, w_eco119569, w_eco119570, w_eco119571, w_eco119572, w_eco119573, w_eco119574, w_eco119575, w_eco119576, w_eco119577, w_eco119578, w_eco119579, w_eco119580, w_eco119581, w_eco119582, w_eco119583, w_eco119584, w_eco119585, w_eco119586, w_eco119587, w_eco119588, w_eco119589, w_eco119590, w_eco119591, w_eco119592, w_eco119593, w_eco119594, w_eco119595, w_eco119596, w_eco119597, w_eco119598, w_eco119599, w_eco119600, w_eco119601, w_eco119602, w_eco119603, w_eco119604, w_eco119605, w_eco119606, w_eco119607, w_eco119608, w_eco119609, w_eco119610, w_eco119611, w_eco119612, w_eco119613, w_eco119614, w_eco119615, w_eco119616, w_eco119617, w_eco119618, w_eco119619, w_eco119620, w_eco119621, w_eco119622, w_eco119623, w_eco119624, w_eco119625, w_eco119626, w_eco119627, w_eco119628, w_eco119629, w_eco119630, w_eco119631, w_eco119632, w_eco119633, w_eco119634, w_eco119635, w_eco119636, w_eco119637, w_eco119638, w_eco119639, w_eco119640, w_eco119641, w_eco119642, w_eco119643, w_eco119644, w_eco119645, w_eco119646, w_eco119647, w_eco119648, w_eco119649, w_eco119650, w_eco119651, w_eco119652, w_eco119653, w_eco119654, w_eco119655, w_eco119656, w_eco119657, w_eco119658, w_eco119659, w_eco119660, w_eco119661, w_eco119662, w_eco119663, w_eco119664, w_eco119665, w_eco119666, w_eco119667, w_eco119668, w_eco119669, w_eco119670, w_eco119671, w_eco119672, w_eco119673, w_eco119674, w_eco119675, w_eco119676, w_eco119677, w_eco119678, w_eco119679, w_eco119680, w_eco119681, w_eco119682, w_eco119683, w_eco119684, w_eco119685, w_eco119686, w_eco119687, w_eco119688, w_eco119689, w_eco119690, w_eco119691, w_eco119692, w_eco119693, w_eco119694, w_eco119695, w_eco119696, w_eco119697, w_eco119698, w_eco119699, w_eco119700, w_eco119701, w_eco119702, w_eco119703, w_eco119704, w_eco119705, w_eco119706, w_eco119707, w_eco119708, w_eco119709, w_eco119710, w_eco119711, w_eco119712, w_eco119713, w_eco119714, w_eco119715, w_eco119716, w_eco119717, w_eco119718, w_eco119719, w_eco119720, w_eco119721, w_eco119722, w_eco119723, w_eco119724, w_eco119725, w_eco119726, w_eco119727, w_eco119728, w_eco119729, w_eco119730, w_eco119731, w_eco119732, w_eco119733, w_eco119734, w_eco119735, w_eco119736, w_eco119737, w_eco119738, w_eco119739, w_eco119740, w_eco119741, w_eco119742, w_eco119743, w_eco119744, w_eco119745, w_eco119746, w_eco119747, w_eco119748, w_eco119749, w_eco119750, w_eco119751, w_eco119752, w_eco119753, w_eco119754, w_eco119755, w_eco119756, w_eco119757, w_eco119758, w_eco119759, w_eco119760, w_eco119761, w_eco119762, w_eco119763, w_eco119764, w_eco119765, w_eco119766, w_eco119767, w_eco119768, w_eco119769, w_eco119770, w_eco119771, w_eco119772, w_eco119773, w_eco119774, w_eco119775, w_eco119776, w_eco119777, w_eco119778, w_eco119779, w_eco119780, w_eco119781, w_eco119782, w_eco119783, w_eco119784, w_eco119785, w_eco119786, w_eco119787, w_eco119788, w_eco119789, w_eco119790, w_eco119791, w_eco119792, w_eco119793, w_eco119794, w_eco119795, w_eco119796, w_eco119797, w_eco119798, w_eco119799, w_eco119800, w_eco119801, w_eco119802, w_eco119803, w_eco119804, w_eco119805, w_eco119806, w_eco119807, w_eco119808, w_eco119809, w_eco119810, w_eco119811, w_eco119812, w_eco119813, w_eco119814, w_eco119815, w_eco119816, w_eco119817, w_eco119818, w_eco119819, w_eco119820, w_eco119821, w_eco119822, w_eco119823, w_eco119824, w_eco119825, w_eco119826, w_eco119827, w_eco119828, w_eco119829, w_eco119830, w_eco119831, w_eco119832, w_eco119833, w_eco119834, w_eco119835, w_eco119836, w_eco119837, w_eco119838, w_eco119839, w_eco119840, w_eco119841, w_eco119842, w_eco119843, w_eco119844, w_eco119845, w_eco119846, w_eco119847, w_eco119848, w_eco119849, w_eco119850, w_eco119851, w_eco119852, w_eco119853, w_eco119854, w_eco119855, w_eco119856, w_eco119857, w_eco119858, w_eco119859, w_eco119860, w_eco119861, w_eco119862, w_eco119863, w_eco119864, w_eco119865, w_eco119866, w_eco119867, w_eco119868, w_eco119869, w_eco119870, w_eco119871, w_eco119872, w_eco119873, w_eco119874, w_eco119875, w_eco119876, w_eco119877, w_eco119878, w_eco119879, w_eco119880, w_eco119881, w_eco119882, w_eco119883, w_eco119884, w_eco119885, w_eco119886, w_eco119887, w_eco119888, w_eco119889, w_eco119890, w_eco119891, w_eco119892, w_eco119893, w_eco119894, w_eco119895, w_eco119896, w_eco119897, w_eco119898, w_eco119899, w_eco119900, w_eco119901, w_eco119902, w_eco119903, w_eco119904, w_eco119905, w_eco119906, w_eco119907, w_eco119908, w_eco119909, w_eco119910, w_eco119911, w_eco119912, w_eco119913, w_eco119914, w_eco119915, w_eco119916, w_eco119917, w_eco119918, w_eco119919, w_eco119920, w_eco119921, w_eco119922, w_eco119923, w_eco119924, w_eco119925, w_eco119926, w_eco119927, w_eco119928, w_eco119929, w_eco119930, w_eco119931, w_eco119932, w_eco119933, w_eco119934, w_eco119935, w_eco119936, w_eco119937, w_eco119938, w_eco119939, w_eco119940, w_eco119941, w_eco119942, w_eco119943, w_eco119944, w_eco119945, w_eco119946, w_eco119947, w_eco119948, w_eco119949, w_eco119950, w_eco119951, w_eco119952, w_eco119953, w_eco119954, w_eco119955, w_eco119956, w_eco119957, w_eco119958, w_eco119959, w_eco119960, w_eco119961, w_eco119962, w_eco119963, w_eco119964, w_eco119965, w_eco119966, w_eco119967, w_eco119968, w_eco119969, w_eco119970, w_eco119971, w_eco119972, w_eco119973, w_eco119974, w_eco119975, w_eco119976, w_eco119977, w_eco119978, w_eco119979, w_eco119980, w_eco119981, w_eco119982, w_eco119983, w_eco119984, w_eco119985, w_eco119986, w_eco119987, w_eco119988, w_eco119989, w_eco119990, w_eco119991, w_eco119992, w_eco119993, w_eco119994, w_eco119995, w_eco119996, w_eco119997, w_eco119998, w_eco119999, w_eco120000, w_eco120001, w_eco120002, w_eco120003, w_eco120004, w_eco120005, w_eco120006, w_eco120007, w_eco120008, w_eco120009, w_eco120010, w_eco120011, w_eco120012, w_eco120013, w_eco120014, w_eco120015, w_eco120016, w_eco120017, w_eco120018, w_eco120019, w_eco120020, w_eco120021, w_eco120022, w_eco120023, w_eco120024, w_eco120025, w_eco120026, w_eco120027, w_eco120028, w_eco120029, w_eco120030, w_eco120031, w_eco120032, w_eco120033, w_eco120034, w_eco120035, w_eco120036, w_eco120037, w_eco120038, w_eco120039, w_eco120040, w_eco120041, w_eco120042, w_eco120043, w_eco120044, w_eco120045, w_eco120046, w_eco120047, w_eco120048, w_eco120049, w_eco120050, w_eco120051, w_eco120052, w_eco120053, w_eco120054, w_eco120055, w_eco120056, w_eco120057, w_eco120058, w_eco120059, w_eco120060, w_eco120061, w_eco120062, w_eco120063, w_eco120064, w_eco120065, w_eco120066, w_eco120067, w_eco120068, w_eco120069, w_eco120070, w_eco120071, w_eco120072, w_eco120073, w_eco120074, w_eco120075, w_eco120076, w_eco120077, w_eco120078, w_eco120079, w_eco120080, w_eco120081, w_eco120082, w_eco120083, w_eco120084, w_eco120085, w_eco120086, w_eco120087, w_eco120088, w_eco120089, w_eco120090, w_eco120091, w_eco120092, w_eco120093, w_eco120094, w_eco120095, w_eco120096, w_eco120097, w_eco120098, w_eco120099, w_eco120100, w_eco120101, w_eco120102, w_eco120103, w_eco120104, w_eco120105, w_eco120106, w_eco120107, w_eco120108, w_eco120109, w_eco120110, w_eco120111, w_eco120112, w_eco120113, w_eco120114, w_eco120115, w_eco120116, w_eco120117, w_eco120118, w_eco120119, w_eco120120, w_eco120121, w_eco120122, w_eco120123, w_eco120124, w_eco120125, w_eco120126, w_eco120127, w_eco120128, w_eco120129, w_eco120130, w_eco120131, w_eco120132, w_eco120133, w_eco120134, w_eco120135, w_eco120136, w_eco120137, w_eco120138, w_eco120139, w_eco120140, w_eco120141, w_eco120142, w_eco120143, w_eco120144, w_eco120145, w_eco120146, w_eco120147, w_eco120148, w_eco120149, w_eco120150, w_eco120151, w_eco120152, w_eco120153, w_eco120154, w_eco120155, w_eco120156, w_eco120157, w_eco120158, w_eco120159, w_eco120160, w_eco120161, w_eco120162, w_eco120163, w_eco120164, w_eco120165, w_eco120166, w_eco120167, w_eco120168, w_eco120169, w_eco120170, w_eco120171, w_eco120172, w_eco120173, w_eco120174, w_eco120175, w_eco120176, w_eco120177, w_eco120178, w_eco120179, w_eco120180, w_eco120181, w_eco120182, w_eco120183, w_eco120184, w_eco120185, w_eco120186, w_eco120187, w_eco120188, w_eco120189, w_eco120190, w_eco120191, w_eco120192, w_eco120193, w_eco120194, w_eco120195, w_eco120196, w_eco120197, w_eco120198, w_eco120199, w_eco120200, w_eco120201, w_eco120202, w_eco120203, w_eco120204, w_eco120205, w_eco120206, w_eco120207, w_eco120208, w_eco120209, w_eco120210, w_eco120211, w_eco120212, w_eco120213, w_eco120214, w_eco120215, w_eco120216, w_eco120217, w_eco120218, w_eco120219, w_eco120220, w_eco120221, w_eco120222, w_eco120223, w_eco120224, w_eco120225, w_eco120226, w_eco120227, w_eco120228, w_eco120229, w_eco120230, w_eco120231, w_eco120232, w_eco120233, w_eco120234, w_eco120235, w_eco120236, w_eco120237, w_eco120238, w_eco120239, w_eco120240, w_eco120241, w_eco120242, w_eco120243, w_eco120244, w_eco120245, w_eco120246, w_eco120247, w_eco120248, w_eco120249, w_eco120250, w_eco120251, w_eco120252, w_eco120253, w_eco120254, w_eco120255, w_eco120256, w_eco120257, w_eco120258, w_eco120259, w_eco120260, w_eco120261, w_eco120262, w_eco120263, w_eco120264, w_eco120265, w_eco120266, w_eco120267, w_eco120268, w_eco120269, w_eco120270, w_eco120271, w_eco120272, w_eco120273, w_eco120274, w_eco120275, w_eco120276, w_eco120277, w_eco120278, w_eco120279, w_eco120280, w_eco120281, w_eco120282, w_eco120283, w_eco120284, w_eco120285, w_eco120286, w_eco120287, w_eco120288, w_eco120289, w_eco120290, w_eco120291, w_eco120292, w_eco120293, w_eco120294, w_eco120295, w_eco120296, w_eco120297, w_eco120298, w_eco120299, w_eco120300, w_eco120301, w_eco120302, w_eco120303, w_eco120304, w_eco120305, w_eco120306, w_eco120307, w_eco120308, w_eco120309, w_eco120310, w_eco120311, w_eco120312, w_eco120313, w_eco120314, w_eco120315, w_eco120316, w_eco120317, w_eco120318, w_eco120319, w_eco120320, w_eco120321, w_eco120322, w_eco120323, w_eco120324, w_eco120325, w_eco120326, w_eco120327, w_eco120328, w_eco120329, w_eco120330, w_eco120331, w_eco120332, w_eco120333, w_eco120334, w_eco120335, w_eco120336, w_eco120337, w_eco120338, w_eco120339, w_eco120340, w_eco120341, w_eco120342, w_eco120343, w_eco120344, w_eco120345, w_eco120346, w_eco120347, w_eco120348, w_eco120349, w_eco120350, w_eco120351, w_eco120352, w_eco120353, w_eco120354, w_eco120355, w_eco120356, w_eco120357, w_eco120358, w_eco120359, w_eco120360, w_eco120361, w_eco120362, w_eco120363, w_eco120364, w_eco120365, w_eco120366, w_eco120367, w_eco120368, w_eco120369, w_eco120370, w_eco120371, w_eco120372, w_eco120373, w_eco120374, w_eco120375, w_eco120376, w_eco120377, w_eco120378, w_eco120379, w_eco120380, w_eco120381, w_eco120382, w_eco120383, w_eco120384, w_eco120385, w_eco120386, w_eco120387, w_eco120388, w_eco120389, w_eco120390, w_eco120391, w_eco120392, w_eco120393, w_eco120394, w_eco120395, w_eco120396, w_eco120397, w_eco120398, w_eco120399, w_eco120400, w_eco120401, w_eco120402, w_eco120403, w_eco120404, w_eco120405, w_eco120406, w_eco120407, w_eco120408, w_eco120409, w_eco120410, w_eco120411, w_eco120412, w_eco120413, w_eco120414, w_eco120415, w_eco120416, w_eco120417, w_eco120418, w_eco120419, w_eco120420, w_eco120421, w_eco120422, w_eco120423, w_eco120424, w_eco120425, w_eco120426, w_eco120427, w_eco120428, w_eco120429, w_eco120430, w_eco120431, w_eco120432, w_eco120433, w_eco120434, w_eco120435, w_eco120436, w_eco120437, w_eco120438, w_eco120439, w_eco120440, w_eco120441, w_eco120442, w_eco120443, w_eco120444, w_eco120445, w_eco120446, w_eco120447, w_eco120448, w_eco120449, w_eco120450, w_eco120451, w_eco120452, w_eco120453, w_eco120454, w_eco120455, w_eco120456, w_eco120457, w_eco120458, w_eco120459, w_eco120460, w_eco120461, w_eco120462, w_eco120463, w_eco120464, w_eco120465, w_eco120466, w_eco120467, w_eco120468, w_eco120469, w_eco120470, w_eco120471, w_eco120472, w_eco120473, w_eco120474, w_eco120475, w_eco120476, w_eco120477, w_eco120478, w_eco120479, w_eco120480, w_eco120481, w_eco120482, w_eco120483, w_eco120484, w_eco120485, w_eco120486, w_eco120487, w_eco120488, w_eco120489, w_eco120490, w_eco120491, w_eco120492, w_eco120493, w_eco120494, w_eco120495, w_eco120496, w_eco120497, w_eco120498, w_eco120499, w_eco120500, w_eco120501, w_eco120502, w_eco120503, w_eco120504, w_eco120505, w_eco120506, w_eco120507, w_eco120508, w_eco120509, w_eco120510, w_eco120511, w_eco120512, w_eco120513, w_eco120514, w_eco120515, w_eco120516, w_eco120517, w_eco120518, w_eco120519, w_eco120520, w_eco120521, w_eco120522, w_eco120523, w_eco120524, w_eco120525, w_eco120526, w_eco120527, w_eco120528, w_eco120529, w_eco120530, w_eco120531, w_eco120532, w_eco120533, w_eco120534, w_eco120535, w_eco120536, w_eco120537, w_eco120538, w_eco120539, w_eco120540, w_eco120541, w_eco120542, w_eco120543, w_eco120544, w_eco120545, w_eco120546, w_eco120547, w_eco120548, w_eco120549, w_eco120550, w_eco120551, w_eco120552, w_eco120553, w_eco120554, w_eco120555, w_eco120556, w_eco120557, w_eco120558, w_eco120559, w_eco120560, w_eco120561, w_eco120562, w_eco120563, w_eco120564, w_eco120565, w_eco120566, w_eco120567, w_eco120568, w_eco120569, w_eco120570, w_eco120571, w_eco120572, w_eco120573, w_eco120574, w_eco120575, w_eco120576, w_eco120577, w_eco120578, w_eco120579, w_eco120580, w_eco120581, w_eco120582, w_eco120583, w_eco120584, w_eco120585, w_eco120586, w_eco120587, w_eco120588, w_eco120589, w_eco120590, w_eco120591, w_eco120592, w_eco120593, w_eco120594, w_eco120595, w_eco120596, w_eco120597, w_eco120598, w_eco120599, w_eco120600, w_eco120601, w_eco120602, w_eco120603, w_eco120604, w_eco120605, w_eco120606, w_eco120607, w_eco120608, w_eco120609, w_eco120610, w_eco120611, w_eco120612, w_eco120613, w_eco120614, w_eco120615, w_eco120616, w_eco120617, w_eco120618, w_eco120619, w_eco120620, w_eco120621, w_eco120622, w_eco120623, w_eco120624, w_eco120625, w_eco120626, w_eco120627, w_eco120628, w_eco120629, w_eco120630, w_eco120631, w_eco120632, w_eco120633, w_eco120634, w_eco120635, w_eco120636, w_eco120637, w_eco120638, w_eco120639, w_eco120640, w_eco120641, w_eco120642, w_eco120643, w_eco120644, w_eco120645, w_eco120646, w_eco120647, w_eco120648, w_eco120649, w_eco120650, w_eco120651, w_eco120652, w_eco120653, w_eco120654, w_eco120655, w_eco120656, w_eco120657, w_eco120658, w_eco120659, w_eco120660, w_eco120661, w_eco120662, w_eco120663, w_eco120664, w_eco120665, w_eco120666, w_eco120667, w_eco120668, w_eco120669, w_eco120670, w_eco120671, w_eco120672, w_eco120673, w_eco120674, w_eco120675, w_eco120676, w_eco120677, w_eco120678, w_eco120679, w_eco120680, w_eco120681, w_eco120682, w_eco120683, w_eco120684, w_eco120685, w_eco120686, w_eco120687, w_eco120688, w_eco120689, w_eco120690, w_eco120691, w_eco120692, w_eco120693, w_eco120694, w_eco120695, w_eco120696, w_eco120697, w_eco120698, w_eco120699, w_eco120700, w_eco120701, w_eco120702, w_eco120703, w_eco120704, w_eco120705, w_eco120706, w_eco120707, w_eco120708, w_eco120709, w_eco120710, w_eco120711, w_eco120712, w_eco120713, w_eco120714, w_eco120715, w_eco120716, w_eco120717, w_eco120718, w_eco120719, w_eco120720, w_eco120721, w_eco120722, w_eco120723, w_eco120724, w_eco120725, w_eco120726, w_eco120727, w_eco120728, w_eco120729, w_eco120730, w_eco120731, w_eco120732, w_eco120733, w_eco120734, w_eco120735, w_eco120736, w_eco120737, w_eco120738, w_eco120739, w_eco120740, w_eco120741, w_eco120742, w_eco120743, w_eco120744, w_eco120745, w_eco120746, w_eco120747, w_eco120748, w_eco120749, w_eco120750, w_eco120751, w_eco120752, w_eco120753, w_eco120754, w_eco120755, w_eco120756, w_eco120757, w_eco120758, w_eco120759, w_eco120760, w_eco120761, w_eco120762, w_eco120763, w_eco120764, w_eco120765, w_eco120766, w_eco120767, w_eco120768, w_eco120769, w_eco120770, w_eco120771, w_eco120772, w_eco120773, w_eco120774, w_eco120775, w_eco120776, w_eco120777, w_eco120778, w_eco120779, w_eco120780, w_eco120781, w_eco120782, w_eco120783, w_eco120784, w_eco120785, w_eco120786, w_eco120787, w_eco120788, w_eco120789, w_eco120790, w_eco120791, w_eco120792, w_eco120793, w_eco120794, w_eco120795, w_eco120796, w_eco120797, w_eco120798, w_eco120799, w_eco120800, w_eco120801, w_eco120802, w_eco120803, w_eco120804, w_eco120805, w_eco120806, w_eco120807, w_eco120808, w_eco120809, w_eco120810, w_eco120811, w_eco120812, w_eco120813, w_eco120814, w_eco120815, w_eco120816, w_eco120817, w_eco120818, w_eco120819, w_eco120820, w_eco120821, w_eco120822, w_eco120823, w_eco120824, w_eco120825, w_eco120826, w_eco120827, w_eco120828, w_eco120829, w_eco120830, w_eco120831, w_eco120832, w_eco120833, w_eco120834, w_eco120835, w_eco120836, w_eco120837, w_eco120838, w_eco120839, w_eco120840, w_eco120841, w_eco120842, w_eco120843, w_eco120844, w_eco120845, w_eco120846, w_eco120847, w_eco120848, w_eco120849, w_eco120850, w_eco120851, w_eco120852, w_eco120853, w_eco120854, w_eco120855, w_eco120856, w_eco120857, w_eco120858, w_eco120859, w_eco120860, w_eco120861, w_eco120862, w_eco120863, w_eco120864, w_eco120865, w_eco120866, w_eco120867, w_eco120868, w_eco120869, w_eco120870, w_eco120871, w_eco120872, w_eco120873, w_eco120874, w_eco120875, w_eco120876, w_eco120877, w_eco120878, w_eco120879, w_eco120880, w_eco120881, w_eco120882, w_eco120883, w_eco120884, w_eco120885, w_eco120886, w_eco120887, w_eco120888, w_eco120889, w_eco120890, w_eco120891, w_eco120892, w_eco120893, w_eco120894, w_eco120895, w_eco120896, w_eco120897, w_eco120898, w_eco120899, w_eco120900, w_eco120901, w_eco120902, w_eco120903, w_eco120904, w_eco120905, w_eco120906, w_eco120907, w_eco120908, w_eco120909, w_eco120910, w_eco120911, w_eco120912, w_eco120913, w_eco120914, w_eco120915, w_eco120916, w_eco120917, w_eco120918, w_eco120919, w_eco120920, w_eco120921, w_eco120922, w_eco120923, w_eco120924, w_eco120925, w_eco120926, w_eco120927, w_eco120928, w_eco120929, w_eco120930, w_eco120931, w_eco120932, w_eco120933, w_eco120934, w_eco120935, w_eco120936, w_eco120937, w_eco120938, w_eco120939, w_eco120940, w_eco120941, w_eco120942, w_eco120943, w_eco120944, w_eco120945, w_eco120946, w_eco120947, w_eco120948, w_eco120949, w_eco120950, w_eco120951, w_eco120952, w_eco120953, w_eco120954, w_eco120955, w_eco120956, w_eco120957, w_eco120958, w_eco120959, w_eco120960, w_eco120961, w_eco120962, w_eco120963, w_eco120964, w_eco120965, w_eco120966, w_eco120967, w_eco120968, w_eco120969, w_eco120970, w_eco120971, w_eco120972, w_eco120973, w_eco120974, w_eco120975, w_eco120976, w_eco120977, w_eco120978, w_eco120979, w_eco120980, w_eco120981, w_eco120982, w_eco120983, w_eco120984, w_eco120985, w_eco120986, w_eco120987, w_eco120988, w_eco120989, w_eco120990, w_eco120991, w_eco120992, w_eco120993, w_eco120994, w_eco120995, w_eco120996, w_eco120997, w_eco120998, w_eco120999, w_eco121000, w_eco121001, w_eco121002, w_eco121003, w_eco121004, w_eco121005, w_eco121006, w_eco121007, w_eco121008, w_eco121009, w_eco121010, w_eco121011, w_eco121012, w_eco121013, w_eco121014, w_eco121015, w_eco121016, w_eco121017, w_eco121018, w_eco121019, w_eco121020, w_eco121021, w_eco121022, w_eco121023, w_eco121024, w_eco121025, w_eco121026, w_eco121027, w_eco121028, w_eco121029, w_eco121030, w_eco121031, w_eco121032, w_eco121033, w_eco121034, w_eco121035, w_eco121036, w_eco121037, w_eco121038, w_eco121039, w_eco121040, w_eco121041, w_eco121042, w_eco121043, w_eco121044, w_eco121045, w_eco121046, w_eco121047, w_eco121048, w_eco121049, w_eco121050, w_eco121051, w_eco121052, w_eco121053, w_eco121054, w_eco121055, w_eco121056, w_eco121057, w_eco121058, w_eco121059, w_eco121060, w_eco121061, w_eco121062, w_eco121063, w_eco121064, w_eco121065, w_eco121066, w_eco121067, w_eco121068, w_eco121069, w_eco121070, w_eco121071, w_eco121072, w_eco121073, w_eco121074, w_eco121075, w_eco121076, w_eco121077, w_eco121078, w_eco121079, w_eco121080, w_eco121081, w_eco121082, w_eco121083, w_eco121084, w_eco121085, w_eco121086, w_eco121087, w_eco121088, w_eco121089, w_eco121090, w_eco121091, w_eco121092, w_eco121093, w_eco121094, w_eco121095, w_eco121096, w_eco121097, w_eco121098, w_eco121099, w_eco121100, w_eco121101, w_eco121102, w_eco121103, w_eco121104, w_eco121105, w_eco121106, w_eco121107, w_eco121108, w_eco121109, w_eco121110, w_eco121111, w_eco121112, w_eco121113, w_eco121114, w_eco121115, w_eco121116, w_eco121117, w_eco121118, w_eco121119, w_eco121120, w_eco121121, w_eco121122, w_eco121123, w_eco121124, w_eco121125, w_eco121126, w_eco121127, w_eco121128, w_eco121129, w_eco121130, w_eco121131, w_eco121132, w_eco121133, w_eco121134, w_eco121135, w_eco121136, w_eco121137, w_eco121138, w_eco121139, w_eco121140, w_eco121141, w_eco121142, w_eco121143, w_eco121144, w_eco121145, w_eco121146, w_eco121147, w_eco121148, w_eco121149, w_eco121150, w_eco121151, w_eco121152, w_eco121153, w_eco121154, w_eco121155, w_eco121156, w_eco121157, w_eco121158, w_eco121159, w_eco121160, w_eco121161, w_eco121162, w_eco121163, w_eco121164, w_eco121165, w_eco121166, w_eco121167, w_eco121168, w_eco121169, w_eco121170, w_eco121171, w_eco121172, w_eco121173, w_eco121174, w_eco121175, w_eco121176, w_eco121177, w_eco121178, w_eco121179, w_eco121180, w_eco121181, w_eco121182, w_eco121183, w_eco121184, w_eco121185, w_eco121186, w_eco121187, w_eco121188, w_eco121189, w_eco121190, w_eco121191, w_eco121192, w_eco121193, w_eco121194, w_eco121195, w_eco121196, w_eco121197, w_eco121198, w_eco121199, w_eco121200, w_eco121201, w_eco121202, w_eco121203, w_eco121204, w_eco121205, w_eco121206, w_eco121207, w_eco121208, w_eco121209, w_eco121210, w_eco121211, w_eco121212, w_eco121213, w_eco121214, w_eco121215, w_eco121216, w_eco121217, w_eco121218, w_eco121219, w_eco121220, w_eco121221, w_eco121222, w_eco121223, w_eco121224, w_eco121225, w_eco121226, w_eco121227, w_eco121228, w_eco121229, w_eco121230, w_eco121231, w_eco121232, w_eco121233, w_eco121234, w_eco121235, w_eco121236, w_eco121237, w_eco121238, w_eco121239, w_eco121240, w_eco121241, w_eco121242, w_eco121243, w_eco121244, w_eco121245, w_eco121246, w_eco121247, w_eco121248, w_eco121249, w_eco121250, w_eco121251, w_eco121252, w_eco121253, w_eco121254, w_eco121255, w_eco121256, w_eco121257, w_eco121258, w_eco121259, w_eco121260, w_eco121261, w_eco121262, w_eco121263, w_eco121264, w_eco121265, w_eco121266, w_eco121267, w_eco121268, w_eco121269, w_eco121270, w_eco121271, w_eco121272, w_eco121273, w_eco121274, w_eco121275, w_eco121276, w_eco121277, w_eco121278, w_eco121279, w_eco121280, w_eco121281, w_eco121282, w_eco121283, w_eco121284, w_eco121285, w_eco121286, w_eco121287, w_eco121288, w_eco121289, w_eco121290, w_eco121291, w_eco121292, w_eco121293, w_eco121294, w_eco121295, w_eco121296, w_eco121297, w_eco121298, w_eco121299, w_eco121300, w_eco121301, w_eco121302, w_eco121303, w_eco121304, w_eco121305, w_eco121306, w_eco121307, w_eco121308, w_eco121309, w_eco121310, w_eco121311, w_eco121312, w_eco121313, w_eco121314, w_eco121315, w_eco121316, w_eco121317, w_eco121318, w_eco121319, w_eco121320, w_eco121321, w_eco121322, w_eco121323, w_eco121324, w_eco121325, w_eco121326, w_eco121327, w_eco121328, w_eco121329, w_eco121330, w_eco121331, w_eco121332, w_eco121333, w_eco121334, w_eco121335, w_eco121336, w_eco121337, w_eco121338, w_eco121339, w_eco121340, w_eco121341, w_eco121342, w_eco121343, w_eco121344, w_eco121345, w_eco121346, w_eco121347, w_eco121348, w_eco121349, w_eco121350, w_eco121351, w_eco121352, w_eco121353, w_eco121354, w_eco121355, w_eco121356, w_eco121357, w_eco121358, w_eco121359, w_eco121360, w_eco121361, w_eco121362, w_eco121363, w_eco121364, w_eco121365, w_eco121366, w_eco121367, w_eco121368, w_eco121369, w_eco121370, w_eco121371, w_eco121372, w_eco121373, w_eco121374, w_eco121375, w_eco121376, w_eco121377, w_eco121378, w_eco121379, w_eco121380, w_eco121381, w_eco121382, w_eco121383, w_eco121384, w_eco121385, w_eco121386, w_eco121387, w_eco121388, w_eco121389, w_eco121390, w_eco121391, w_eco121392, w_eco121393, w_eco121394, w_eco121395, w_eco121396, w_eco121397, w_eco121398, w_eco121399, w_eco121400, w_eco121401, w_eco121402, w_eco121403, w_eco121404, w_eco121405, w_eco121406, w_eco121407, w_eco121408, w_eco121409, w_eco121410, w_eco121411, w_eco121412, w_eco121413, w_eco121414, w_eco121415, w_eco121416, w_eco121417, w_eco121418, w_eco121419, w_eco121420, w_eco121421, w_eco121422, w_eco121423, w_eco121424, w_eco121425, w_eco121426, w_eco121427, w_eco121428, w_eco121429, w_eco121430, w_eco121431, w_eco121432, w_eco121433, w_eco121434, w_eco121435, w_eco121436, w_eco121437, w_eco121438, w_eco121439, w_eco121440, w_eco121441, w_eco121442, w_eco121443, w_eco121444, w_eco121445, w_eco121446, w_eco121447, w_eco121448, w_eco121449, w_eco121450, w_eco121451, w_eco121452, w_eco121453, w_eco121454, w_eco121455, w_eco121456, w_eco121457, w_eco121458, w_eco121459, w_eco121460, w_eco121461, w_eco121462, w_eco121463, w_eco121464, w_eco121465, w_eco121466, w_eco121467, w_eco121468, w_eco121469, w_eco121470, w_eco121471, w_eco121472, w_eco121473, w_eco121474, w_eco121475, w_eco121476, w_eco121477, w_eco121478, w_eco121479, w_eco121480, w_eco121481, w_eco121482, w_eco121483, w_eco121484, w_eco121485, w_eco121486, w_eco121487, w_eco121488, w_eco121489, w_eco121490, w_eco121491, w_eco121492, w_eco121493, w_eco121494, w_eco121495, w_eco121496, w_eco121497, w_eco121498, w_eco121499, w_eco121500, w_eco121501, w_eco121502, w_eco121503, w_eco121504, w_eco121505, w_eco121506, w_eco121507, w_eco121508, w_eco121509, w_eco121510, w_eco121511, w_eco121512, w_eco121513, w_eco121514, w_eco121515, w_eco121516, w_eco121517, w_eco121518, w_eco121519, w_eco121520, w_eco121521, w_eco121522, w_eco121523, w_eco121524, w_eco121525, w_eco121526, w_eco121527, w_eco121528, w_eco121529, w_eco121530, w_eco121531, w_eco121532, w_eco121533, w_eco121534, w_eco121535, w_eco121536, w_eco121537, w_eco121538, w_eco121539, w_eco121540, w_eco121541, w_eco121542, w_eco121543, w_eco121544, w_eco121545, w_eco121546, w_eco121547, w_eco121548, w_eco121549, w_eco121550, w_eco121551, w_eco121552, w_eco121553, w_eco121554, w_eco121555, w_eco121556, w_eco121557, w_eco121558, w_eco121559, w_eco121560, w_eco121561, w_eco121562, w_eco121563, w_eco121564, w_eco121565, w_eco121566, w_eco121567, w_eco121568, w_eco121569, w_eco121570, w_eco121571, w_eco121572, w_eco121573, w_eco121574, w_eco121575, w_eco121576, w_eco121577, w_eco121578, w_eco121579, w_eco121580, w_eco121581, w_eco121582, w_eco121583, w_eco121584, w_eco121585, w_eco121586, w_eco121587, w_eco121588, w_eco121589, w_eco121590, w_eco121591, w_eco121592, w_eco121593, w_eco121594, w_eco121595, w_eco121596, w_eco121597, w_eco121598, w_eco121599, w_eco121600, w_eco121601, w_eco121602, w_eco121603, w_eco121604, w_eco121605, w_eco121606, w_eco121607, w_eco121608, w_eco121609, w_eco121610, w_eco121611, w_eco121612, w_eco121613, w_eco121614, w_eco121615, w_eco121616, w_eco121617, w_eco121618, w_eco121619, w_eco121620, w_eco121621, w_eco121622, w_eco121623, w_eco121624, w_eco121625, w_eco121626, w_eco121627, w_eco121628, w_eco121629, w_eco121630, w_eco121631, w_eco121632, w_eco121633, w_eco121634, w_eco121635, w_eco121636, w_eco121637, w_eco121638, w_eco121639, w_eco121640, w_eco121641, w_eco121642, w_eco121643, w_eco121644, w_eco121645, w_eco121646, w_eco121647, w_eco121648, w_eco121649, w_eco121650, w_eco121651, w_eco121652, w_eco121653, w_eco121654, w_eco121655, w_eco121656, w_eco121657, w_eco121658, w_eco121659, w_eco121660, w_eco121661, w_eco121662, w_eco121663, w_eco121664, w_eco121665, w_eco121666, w_eco121667, w_eco121668, w_eco121669, w_eco121670, w_eco121671, w_eco121672, w_eco121673, w_eco121674, w_eco121675, w_eco121676, w_eco121677, w_eco121678, w_eco121679, w_eco121680, w_eco121681, w_eco121682, w_eco121683, w_eco121684, w_eco121685, w_eco121686, w_eco121687, w_eco121688, w_eco121689, w_eco121690, w_eco121691, w_eco121692, w_eco121693, w_eco121694, w_eco121695, w_eco121696, w_eco121697, w_eco121698, w_eco121699, w_eco121700, w_eco121701, w_eco121702, w_eco121703, w_eco121704, w_eco121705, w_eco121706, w_eco121707, w_eco121708, w_eco121709, w_eco121710, w_eco121711, w_eco121712, w_eco121713, w_eco121714, w_eco121715, w_eco121716, w_eco121717, w_eco121718, w_eco121719, w_eco121720, w_eco121721, w_eco121722, w_eco121723, w_eco121724, w_eco121725, w_eco121726, w_eco121727, w_eco121728, w_eco121729, w_eco121730, w_eco121731, w_eco121732, w_eco121733, w_eco121734, w_eco121735, w_eco121736, w_eco121737, w_eco121738, w_eco121739, w_eco121740, w_eco121741, w_eco121742, w_eco121743, w_eco121744, w_eco121745, w_eco121746, w_eco121747, w_eco121748, w_eco121749, w_eco121750, w_eco121751, w_eco121752, w_eco121753, w_eco121754, w_eco121755, w_eco121756, w_eco121757, w_eco121758, w_eco121759, w_eco121760, w_eco121761, w_eco121762, w_eco121763, w_eco121764, w_eco121765, w_eco121766, w_eco121767, w_eco121768, w_eco121769, w_eco121770, w_eco121771, w_eco121772, w_eco121773, w_eco121774, w_eco121775, w_eco121776, w_eco121777, w_eco121778, w_eco121779, w_eco121780, w_eco121781, w_eco121782, w_eco121783, w_eco121784, w_eco121785, w_eco121786, w_eco121787, w_eco121788, w_eco121789, w_eco121790, w_eco121791, w_eco121792, w_eco121793, w_eco121794, w_eco121795, w_eco121796, w_eco121797, w_eco121798, w_eco121799, w_eco121800, w_eco121801, w_eco121802, w_eco121803, w_eco121804, w_eco121805, w_eco121806, w_eco121807, w_eco121808, w_eco121809, w_eco121810, w_eco121811, w_eco121812, w_eco121813, w_eco121814, w_eco121815, w_eco121816, w_eco121817, w_eco121818, w_eco121819, w_eco121820, w_eco121821, w_eco121822, w_eco121823, w_eco121824, w_eco121825, w_eco121826, w_eco121827, w_eco121828, w_eco121829, w_eco121830, w_eco121831, w_eco121832, w_eco121833, w_eco121834, w_eco121835, w_eco121836, w_eco121837, w_eco121838, w_eco121839, w_eco121840, w_eco121841, w_eco121842, w_eco121843, w_eco121844, w_eco121845, w_eco121846, w_eco121847, w_eco121848, w_eco121849, w_eco121850, w_eco121851, w_eco121852, w_eco121853, w_eco121854, w_eco121855, w_eco121856, w_eco121857, w_eco121858, w_eco121859, w_eco121860, w_eco121861, w_eco121862, w_eco121863, w_eco121864, w_eco121865, w_eco121866, w_eco121867, w_eco121868, w_eco121869, w_eco121870, w_eco121871, w_eco121872, w_eco121873, w_eco121874, w_eco121875, w_eco121876, w_eco121877, w_eco121878, w_eco121879, w_eco121880, w_eco121881, w_eco121882, w_eco121883, w_eco121884, w_eco121885, w_eco121886, w_eco121887, w_eco121888, w_eco121889, w_eco121890, w_eco121891, w_eco121892, w_eco121893, w_eco121894, w_eco121895, w_eco121896, w_eco121897, w_eco121898, w_eco121899, w_eco121900, w_eco121901, w_eco121902, w_eco121903, w_eco121904, w_eco121905, w_eco121906, w_eco121907, w_eco121908, w_eco121909, w_eco121910, w_eco121911, w_eco121912, w_eco121913, w_eco121914, w_eco121915, w_eco121916, w_eco121917, w_eco121918, w_eco121919, w_eco121920, w_eco121921, w_eco121922, w_eco121923, w_eco121924, w_eco121925, w_eco121926, w_eco121927, w_eco121928, w_eco121929, w_eco121930, w_eco121931, w_eco121932, w_eco121933, w_eco121934, w_eco121935, w_eco121936, w_eco121937, w_eco121938, w_eco121939, w_eco121940, w_eco121941, w_eco121942, w_eco121943, w_eco121944, w_eco121945, w_eco121946, w_eco121947, w_eco121948, w_eco121949, w_eco121950, w_eco121951, w_eco121952, w_eco121953, w_eco121954, w_eco121955, w_eco121956, w_eco121957, w_eco121958, w_eco121959, w_eco121960, w_eco121961, w_eco121962, w_eco121963, w_eco121964, w_eco121965, w_eco121966, w_eco121967, w_eco121968, w_eco121969, w_eco121970, w_eco121971, w_eco121972, w_eco121973, w_eco121974, w_eco121975, w_eco121976, w_eco121977, w_eco121978, w_eco121979, w_eco121980, w_eco121981, w_eco121982, w_eco121983, w_eco121984, w_eco121985, w_eco121986, w_eco121987, w_eco121988, w_eco121989, w_eco121990, w_eco121991, w_eco121992, w_eco121993, w_eco121994, w_eco121995, w_eco121996, w_eco121997, w_eco121998, w_eco121999, w_eco122000, w_eco122001, w_eco122002, w_eco122003, w_eco122004, w_eco122005, w_eco122006, w_eco122007, w_eco122008, w_eco122009, w_eco122010, w_eco122011, w_eco122012, w_eco122013, w_eco122014, w_eco122015, w_eco122016, w_eco122017, w_eco122018, w_eco122019, w_eco122020, w_eco122021, w_eco122022, w_eco122023, w_eco122024, w_eco122025, w_eco122026, w_eco122027, w_eco122028, w_eco122029, w_eco122030, w_eco122031, w_eco122032, w_eco122033, w_eco122034, w_eco122035, w_eco122036, w_eco122037, w_eco122038, w_eco122039, w_eco122040, w_eco122041, w_eco122042, w_eco122043, w_eco122044, w_eco122045, w_eco122046, w_eco122047, w_eco122048, w_eco122049, w_eco122050, w_eco122051, w_eco122052, w_eco122053, w_eco122054, w_eco122055, w_eco122056, w_eco122057, w_eco122058, w_eco122059, w_eco122060, w_eco122061, w_eco122062, w_eco122063, w_eco122064, w_eco122065, w_eco122066, w_eco122067, w_eco122068, w_eco122069, w_eco122070, w_eco122071, w_eco122072, w_eco122073, w_eco122074, w_eco122075, w_eco122076, w_eco122077, w_eco122078, w_eco122079, w_eco122080, w_eco122081, w_eco122082, w_eco122083, w_eco122084, w_eco122085, w_eco122086, w_eco122087, w_eco122088, w_eco122089, w_eco122090, w_eco122091, w_eco122092, w_eco122093, w_eco122094, w_eco122095, w_eco122096, w_eco122097, w_eco122098, w_eco122099, w_eco122100, w_eco122101, w_eco122102, w_eco122103, w_eco122104, w_eco122105, w_eco122106, w_eco122107, w_eco122108, w_eco122109, w_eco122110, w_eco122111, w_eco122112, w_eco122113, w_eco122114, w_eco122115, w_eco122116, w_eco122117, w_eco122118, w_eco122119, w_eco122120, w_eco122121, w_eco122122, w_eco122123, w_eco122124, w_eco122125, w_eco122126, w_eco122127, w_eco122128, w_eco122129, w_eco122130, w_eco122131, w_eco122132, w_eco122133, w_eco122134, w_eco122135, w_eco122136, w_eco122137, w_eco122138, w_eco122139, w_eco122140, w_eco122141, w_eco122142, w_eco122143, w_eco122144, w_eco122145, w_eco122146, w_eco122147, w_eco122148, w_eco122149, w_eco122150, w_eco122151, w_eco122152, w_eco122153, w_eco122154, w_eco122155, w_eco122156, w_eco122157, w_eco122158, w_eco122159, w_eco122160, w_eco122161, w_eco122162, w_eco122163, w_eco122164, w_eco122165, w_eco122166, w_eco122167, w_eco122168, w_eco122169, w_eco122170, w_eco122171, w_eco122172, w_eco122173, w_eco122174, w_eco122175, w_eco122176, w_eco122177, w_eco122178, w_eco122179, w_eco122180, w_eco122181, w_eco122182, w_eco122183, w_eco122184, w_eco122185, w_eco122186, w_eco122187, w_eco122188, w_eco122189, w_eco122190, w_eco122191, w_eco122192, w_eco122193, w_eco122194, w_eco122195, w_eco122196, w_eco122197, w_eco122198, w_eco122199, w_eco122200, w_eco122201, w_eco122202, w_eco122203, w_eco122204, w_eco122205, w_eco122206, w_eco122207, w_eco122208, w_eco122209, w_eco122210, w_eco122211, w_eco122212, w_eco122213, w_eco122214, w_eco122215, w_eco122216, w_eco122217, w_eco122218, w_eco122219, w_eco122220, w_eco122221, w_eco122222, w_eco122223, w_eco122224, w_eco122225, w_eco122226, w_eco122227, w_eco122228, w_eco122229, w_eco122230, w_eco122231, w_eco122232, w_eco122233, w_eco122234, w_eco122235, w_eco122236, w_eco122237, w_eco122238, w_eco122239, w_eco122240, w_eco122241, w_eco122242, w_eco122243, w_eco122244, w_eco122245, w_eco122246, w_eco122247, w_eco122248, w_eco122249, w_eco122250, w_eco122251, w_eco122252, w_eco122253, w_eco122254, w_eco122255, w_eco122256, w_eco122257, w_eco122258, w_eco122259, w_eco122260, w_eco122261, w_eco122262, w_eco122263, w_eco122264, w_eco122265, w_eco122266, w_eco122267, w_eco122268, w_eco122269, w_eco122270, w_eco122271, w_eco122272, w_eco122273, w_eco122274, w_eco122275, w_eco122276, w_eco122277, w_eco122278, w_eco122279, w_eco122280, w_eco122281, w_eco122282, w_eco122283, w_eco122284, w_eco122285, w_eco122286, w_eco122287, w_eco122288, w_eco122289, w_eco122290, w_eco122291, w_eco122292, w_eco122293, w_eco122294, w_eco122295, w_eco122296, w_eco122297, w_eco122298, w_eco122299, w_eco122300, w_eco122301, w_eco122302, w_eco122303, w_eco122304, w_eco122305, w_eco122306, w_eco122307, w_eco122308, w_eco122309, w_eco122310, w_eco122311, w_eco122312, w_eco122313, w_eco122314, w_eco122315, w_eco122316, w_eco122317, w_eco122318, w_eco122319, w_eco122320, w_eco122321, w_eco122322, w_eco122323, w_eco122324, w_eco122325, w_eco122326, w_eco122327, w_eco122328, w_eco122329, w_eco122330, w_eco122331, w_eco122332, w_eco122333, w_eco122334, w_eco122335, w_eco122336, w_eco122337, w_eco122338, w_eco122339, w_eco122340, w_eco122341, w_eco122342, w_eco122343, w_eco122344, w_eco122345, w_eco122346, w_eco122347, w_eco122348, w_eco122349, w_eco122350, w_eco122351, w_eco122352, w_eco122353, w_eco122354, w_eco122355, w_eco122356, w_eco122357, w_eco122358, w_eco122359, w_eco122360, w_eco122361, w_eco122362, w_eco122363, w_eco122364, w_eco122365, w_eco122366, w_eco122367, w_eco122368, w_eco122369, w_eco122370, w_eco122371, w_eco122372, w_eco122373, w_eco122374, w_eco122375, w_eco122376, w_eco122377, w_eco122378, w_eco122379, w_eco122380, w_eco122381, w_eco122382, w_eco122383, w_eco122384, w_eco122385, w_eco122386, w_eco122387, w_eco122388, w_eco122389, w_eco122390, w_eco122391, w_eco122392, w_eco122393, w_eco122394, w_eco122395, w_eco122396, w_eco122397, w_eco122398, w_eco122399, w_eco122400, w_eco122401, w_eco122402, w_eco122403, w_eco122404, w_eco122405, w_eco122406, w_eco122407, w_eco122408, w_eco122409, w_eco122410, w_eco122411, w_eco122412, w_eco122413, w_eco122414, w_eco122415, w_eco122416, w_eco122417, w_eco122418, w_eco122419, w_eco122420, w_eco122421, w_eco122422, w_eco122423, w_eco122424, w_eco122425, w_eco122426, w_eco122427, w_eco122428, w_eco122429, w_eco122430, w_eco122431, w_eco122432, w_eco122433, w_eco122434, w_eco122435, w_eco122436, w_eco122437, w_eco122438, w_eco122439, w_eco122440, w_eco122441, w_eco122442, w_eco122443, w_eco122444, w_eco122445, w_eco122446, w_eco122447, w_eco122448, w_eco122449, w_eco122450, w_eco122451, w_eco122452, w_eco122453, w_eco122454, w_eco122455, w_eco122456, w_eco122457, w_eco122458, w_eco122459, w_eco122460, w_eco122461, w_eco122462, w_eco122463, w_eco122464, w_eco122465, w_eco122466, w_eco122467, w_eco122468, w_eco122469, w_eco122470, w_eco122471, w_eco122472, w_eco122473, w_eco122474, w_eco122475, w_eco122476, w_eco122477, w_eco122478, w_eco122479, w_eco122480, w_eco122481, w_eco122482, w_eco122483, w_eco122484, w_eco122485, w_eco122486, w_eco122487, w_eco122488, w_eco122489, w_eco122490, w_eco122491, w_eco122492, w_eco122493, w_eco122494, w_eco122495, w_eco122496, w_eco122497, w_eco122498, w_eco122499, w_eco122500, w_eco122501, w_eco122502, w_eco122503, w_eco122504, w_eco122505, w_eco122506, w_eco122507, w_eco122508, w_eco122509, w_eco122510, w_eco122511, w_eco122512, w_eco122513, w_eco122514, w_eco122515, w_eco122516, w_eco122517, w_eco122518, w_eco122519, w_eco122520, w_eco122521, w_eco122522, w_eco122523, w_eco122524, w_eco122525, w_eco122526, w_eco122527, w_eco122528, w_eco122529, w_eco122530, w_eco122531, w_eco122532, w_eco122533, w_eco122534, w_eco122535, w_eco122536, w_eco122537, w_eco122538, w_eco122539, w_eco122540, w_eco122541, w_eco122542, w_eco122543, w_eco122544, w_eco122545, w_eco122546, w_eco122547, w_eco122548, w_eco122549, w_eco122550, w_eco122551, w_eco122552, w_eco122553, w_eco122554, w_eco122555, w_eco122556, w_eco122557, w_eco122558, w_eco122559, w_eco122560, w_eco122561, w_eco122562, w_eco122563, w_eco122564, w_eco122565, w_eco122566, w_eco122567, w_eco122568, w_eco122569, w_eco122570, w_eco122571, w_eco122572, w_eco122573, w_eco122574, w_eco122575, w_eco122576, w_eco122577, w_eco122578, w_eco122579, w_eco122580, w_eco122581, w_eco122582, w_eco122583, w_eco122584, w_eco122585, w_eco122586, w_eco122587, w_eco122588, w_eco122589, w_eco122590, w_eco122591, w_eco122592, w_eco122593, w_eco122594, w_eco122595, w_eco122596, w_eco122597, w_eco122598, w_eco122599, w_eco122600, w_eco122601, w_eco122602, w_eco122603, w_eco122604, w_eco122605, w_eco122606, w_eco122607, w_eco122608, w_eco122609, w_eco122610, w_eco122611, w_eco122612, w_eco122613, w_eco122614, w_eco122615, w_eco122616, w_eco122617, w_eco122618, w_eco122619, w_eco122620, w_eco122621, w_eco122622, w_eco122623, w_eco122624, w_eco122625, w_eco122626, w_eco122627, w_eco122628, w_eco122629, w_eco122630, w_eco122631, w_eco122632, w_eco122633, w_eco122634, w_eco122635, w_eco122636, w_eco122637, w_eco122638, w_eco122639, w_eco122640, w_eco122641, w_eco122642, w_eco122643, w_eco122644, w_eco122645, w_eco122646, w_eco122647, w_eco122648, w_eco122649, w_eco122650, w_eco122651, w_eco122652, w_eco122653, w_eco122654, w_eco122655, w_eco122656, w_eco122657, w_eco122658, w_eco122659, w_eco122660, w_eco122661, w_eco122662, w_eco122663, w_eco122664, w_eco122665, w_eco122666, w_eco122667, w_eco122668, w_eco122669, w_eco122670, w_eco122671, w_eco122672, w_eco122673, w_eco122674, w_eco122675, w_eco122676, w_eco122677, w_eco122678, w_eco122679, w_eco122680, w_eco122681, w_eco122682, w_eco122683, w_eco122684, w_eco122685, w_eco122686, w_eco122687, w_eco122688, w_eco122689, w_eco122690, w_eco122691, w_eco122692, w_eco122693, w_eco122694, w_eco122695, w_eco122696, w_eco122697, w_eco122698, w_eco122699, w_eco122700, w_eco122701, w_eco122702, w_eco122703, w_eco122704, w_eco122705, w_eco122706, w_eco122707, w_eco122708, w_eco122709, w_eco122710, w_eco122711, w_eco122712, w_eco122713, w_eco122714, w_eco122715, w_eco122716, w_eco122717, w_eco122718, w_eco122719, w_eco122720, w_eco122721, w_eco122722, w_eco122723, w_eco122724, w_eco122725, w_eco122726, w_eco122727, w_eco122728, w_eco122729, w_eco122730, w_eco122731, w_eco122732, w_eco122733, w_eco122734, w_eco122735, w_eco122736, w_eco122737, w_eco122738, w_eco122739, w_eco122740, w_eco122741, w_eco122742, w_eco122743, w_eco122744, w_eco122745, w_eco122746, w_eco122747, w_eco122748, w_eco122749, w_eco122750, w_eco122751, w_eco122752, w_eco122753, w_eco122754, w_eco122755, w_eco122756, w_eco122757, w_eco122758, w_eco122759, w_eco122760, w_eco122761, w_eco122762, w_eco122763, w_eco122764, w_eco122765, w_eco122766, w_eco122767, w_eco122768, w_eco122769, w_eco122770, w_eco122771, w_eco122772, w_eco122773, w_eco122774, w_eco122775, w_eco122776, w_eco122777, w_eco122778, w_eco122779, w_eco122780, w_eco122781, w_eco122782, w_eco122783, w_eco122784, w_eco122785, w_eco122786, w_eco122787, w_eco122788, w_eco122789, w_eco122790, w_eco122791, w_eco122792, w_eco122793, w_eco122794, w_eco122795, w_eco122796, w_eco122797, w_eco122798, w_eco122799, w_eco122800, w_eco122801, w_eco122802, w_eco122803, w_eco122804, w_eco122805, w_eco122806, w_eco122807, w_eco122808, w_eco122809, w_eco122810, w_eco122811, w_eco122812, w_eco122813, w_eco122814, w_eco122815, w_eco122816, w_eco122817, w_eco122818, w_eco122819, w_eco122820, w_eco122821, w_eco122822, w_eco122823, w_eco122824, w_eco122825, w_eco122826, w_eco122827, w_eco122828, w_eco122829, w_eco122830, w_eco122831, w_eco122832, w_eco122833, w_eco122834, w_eco122835, w_eco122836, w_eco122837, w_eco122838, w_eco122839, w_eco122840, w_eco122841, w_eco122842, w_eco122843, w_eco122844, w_eco122845, w_eco122846, w_eco122847, w_eco122848, w_eco122849, w_eco122850, w_eco122851, w_eco122852, w_eco122853, w_eco122854, w_eco122855, w_eco122856, w_eco122857, w_eco122858, w_eco122859, w_eco122860, w_eco122861, w_eco122862, w_eco122863, w_eco122864, w_eco122865, w_eco122866, w_eco122867, w_eco122868, w_eco122869, w_eco122870, w_eco122871, w_eco122872, w_eco122873, w_eco122874, w_eco122875, w_eco122876, w_eco122877, w_eco122878, w_eco122879, w_eco122880, w_eco122881, w_eco122882, w_eco122883, w_eco122884, w_eco122885, w_eco122886, w_eco122887, w_eco122888, w_eco122889, w_eco122890, w_eco122891, w_eco122892, w_eco122893, w_eco122894, w_eco122895, w_eco122896, w_eco122897, w_eco122898, w_eco122899, w_eco122900, w_eco122901, w_eco122902, w_eco122903, w_eco122904, w_eco122905, w_eco122906, w_eco122907, w_eco122908, w_eco122909, w_eco122910, w_eco122911, w_eco122912, w_eco122913, w_eco122914, w_eco122915, w_eco122916, w_eco122917, w_eco122918, w_eco122919, w_eco122920, w_eco122921, w_eco122922, w_eco122923, w_eco122924, w_eco122925, w_eco122926, w_eco122927, w_eco122928, w_eco122929, w_eco122930, w_eco122931, w_eco122932, w_eco122933, w_eco122934, w_eco122935, w_eco122936, w_eco122937, w_eco122938, w_eco122939, w_eco122940, w_eco122941, w_eco122942, w_eco122943, w_eco122944, w_eco122945, w_eco122946, w_eco122947, w_eco122948, w_eco122949, w_eco122950, w_eco122951, w_eco122952, w_eco122953, w_eco122954, w_eco122955, w_eco122956, w_eco122957, w_eco122958, w_eco122959, w_eco122960, w_eco122961, w_eco122962, w_eco122963, w_eco122964, w_eco122965, w_eco122966, w_eco122967, w_eco122968, w_eco122969, w_eco122970, w_eco122971, w_eco122972, w_eco122973, w_eco122974, w_eco122975, w_eco122976, w_eco122977, w_eco122978, w_eco122979, w_eco122980, w_eco122981, w_eco122982, w_eco122983, w_eco122984, w_eco122985, w_eco122986, w_eco122987, w_eco122988, w_eco122989, w_eco122990, w_eco122991, w_eco122992, w_eco122993, w_eco122994, w_eco122995, w_eco122996, w_eco122997, w_eco122998, w_eco122999, w_eco123000, w_eco123001, w_eco123002, w_eco123003, w_eco123004, w_eco123005, w_eco123006, w_eco123007, w_eco123008, w_eco123009, w_eco123010, w_eco123011, w_eco123012, w_eco123013, w_eco123014, w_eco123015, w_eco123016, w_eco123017, w_eco123018, w_eco123019, w_eco123020, w_eco123021, w_eco123022, w_eco123023, w_eco123024, w_eco123025, w_eco123026, w_eco123027, w_eco123028, w_eco123029, w_eco123030, w_eco123031, w_eco123032, w_eco123033, w_eco123034, w_eco123035, w_eco123036, w_eco123037, w_eco123038, w_eco123039, w_eco123040, w_eco123041, w_eco123042, w_eco123043, w_eco123044, w_eco123045, w_eco123046, w_eco123047, w_eco123048, w_eco123049, w_eco123050, w_eco123051, w_eco123052, w_eco123053, w_eco123054, w_eco123055, w_eco123056, w_eco123057, w_eco123058, w_eco123059, w_eco123060, w_eco123061, w_eco123062, w_eco123063, w_eco123064, w_eco123065, w_eco123066, w_eco123067, w_eco123068, w_eco123069, w_eco123070, w_eco123071, w_eco123072, w_eco123073, w_eco123074, w_eco123075, w_eco123076, w_eco123077, w_eco123078, w_eco123079, w_eco123080, w_eco123081, w_eco123082, w_eco123083, w_eco123084, w_eco123085, w_eco123086, w_eco123087, w_eco123088, w_eco123089, w_eco123090, w_eco123091, w_eco123092, w_eco123093, w_eco123094, w_eco123095, w_eco123096, w_eco123097, w_eco123098, w_eco123099, w_eco123100, w_eco123101, w_eco123102, w_eco123103, w_eco123104, w_eco123105, w_eco123106, w_eco123107, w_eco123108, w_eco123109, w_eco123110, w_eco123111, w_eco123112, w_eco123113, w_eco123114, w_eco123115, w_eco123116, w_eco123117, w_eco123118, w_eco123119, w_eco123120, w_eco123121, w_eco123122, w_eco123123, w_eco123124, w_eco123125, w_eco123126, w_eco123127, w_eco123128, w_eco123129, w_eco123130, w_eco123131, w_eco123132, w_eco123133, w_eco123134, w_eco123135, w_eco123136, w_eco123137, w_eco123138, w_eco123139, w_eco123140, w_eco123141, w_eco123142, w_eco123143, w_eco123144, w_eco123145, w_eco123146, w_eco123147, w_eco123148, w_eco123149, w_eco123150, w_eco123151, w_eco123152, w_eco123153, w_eco123154, w_eco123155, w_eco123156, w_eco123157, w_eco123158, w_eco123159, w_eco123160, w_eco123161, w_eco123162, w_eco123163, w_eco123164, w_eco123165, w_eco123166, w_eco123167, w_eco123168, w_eco123169, w_eco123170, w_eco123171, w_eco123172, w_eco123173, w_eco123174, w_eco123175, w_eco123176, w_eco123177, w_eco123178, w_eco123179, w_eco123180, w_eco123181, w_eco123182, w_eco123183, w_eco123184, w_eco123185, w_eco123186, w_eco123187, w_eco123188, w_eco123189, w_eco123190, w_eco123191, w_eco123192, w_eco123193, w_eco123194, w_eco123195, w_eco123196, w_eco123197, w_eco123198, w_eco123199, w_eco123200, w_eco123201, w_eco123202, w_eco123203, w_eco123204, w_eco123205, w_eco123206, w_eco123207, w_eco123208, w_eco123209, w_eco123210, w_eco123211, w_eco123212, w_eco123213, w_eco123214, w_eco123215, w_eco123216, w_eco123217, w_eco123218, w_eco123219, w_eco123220, w_eco123221, w_eco123222, w_eco123223, w_eco123224, w_eco123225, w_eco123226, w_eco123227, w_eco123228, w_eco123229, w_eco123230, w_eco123231, w_eco123232, w_eco123233, w_eco123234, w_eco123235, w_eco123236, w_eco123237, w_eco123238, w_eco123239, w_eco123240, w_eco123241, w_eco123242, w_eco123243, w_eco123244, w_eco123245, w_eco123246, w_eco123247, w_eco123248, w_eco123249, w_eco123250, w_eco123251, w_eco123252, w_eco123253, w_eco123254, w_eco123255, w_eco123256, w_eco123257, w_eco123258, w_eco123259, w_eco123260, w_eco123261, w_eco123262, w_eco123263, w_eco123264, w_eco123265, w_eco123266, w_eco123267, w_eco123268, w_eco123269, w_eco123270, w_eco123271, w_eco123272, w_eco123273, w_eco123274, w_eco123275, w_eco123276, w_eco123277, w_eco123278, w_eco123279, w_eco123280, w_eco123281, w_eco123282, w_eco123283, w_eco123284, w_eco123285, w_eco123286, w_eco123287, w_eco123288, w_eco123289, w_eco123290, w_eco123291, w_eco123292, w_eco123293, w_eco123294, w_eco123295, w_eco123296, w_eco123297, w_eco123298, w_eco123299, w_eco123300, w_eco123301, w_eco123302, w_eco123303, w_eco123304, w_eco123305, w_eco123306, w_eco123307, w_eco123308, w_eco123309, w_eco123310, w_eco123311, w_eco123312, w_eco123313, w_eco123314, w_eco123315, w_eco123316, w_eco123317, w_eco123318, w_eco123319, w_eco123320, w_eco123321, w_eco123322, w_eco123323, w_eco123324, w_eco123325, w_eco123326, w_eco123327, w_eco123328, w_eco123329, w_eco123330, w_eco123331, w_eco123332, w_eco123333, w_eco123334, w_eco123335, w_eco123336, w_eco123337, w_eco123338, w_eco123339, w_eco123340, w_eco123341, w_eco123342, w_eco123343, w_eco123344, w_eco123345, w_eco123346, w_eco123347, w_eco123348, w_eco123349, w_eco123350, w_eco123351, w_eco123352, w_eco123353, w_eco123354, w_eco123355, w_eco123356, w_eco123357, w_eco123358, w_eco123359, w_eco123360, w_eco123361, w_eco123362, w_eco123363, w_eco123364, w_eco123365, w_eco123366, w_eco123367, w_eco123368, w_eco123369, w_eco123370, w_eco123371, w_eco123372, w_eco123373, w_eco123374, w_eco123375, w_eco123376, w_eco123377, w_eco123378, w_eco123379, w_eco123380, w_eco123381, w_eco123382, w_eco123383, w_eco123384, w_eco123385, w_eco123386, w_eco123387, w_eco123388, w_eco123389, w_eco123390, w_eco123391, w_eco123392, w_eco123393, w_eco123394, w_eco123395, w_eco123396, w_eco123397, w_eco123398, w_eco123399, w_eco123400, w_eco123401, w_eco123402, w_eco123403, w_eco123404, w_eco123405, w_eco123406, w_eco123407, w_eco123408, w_eco123409, w_eco123410, w_eco123411, w_eco123412, w_eco123413, w_eco123414, w_eco123415, w_eco123416, w_eco123417, w_eco123418, w_eco123419, w_eco123420, w_eco123421, w_eco123422, w_eco123423, w_eco123424, w_eco123425, w_eco123426, w_eco123427, w_eco123428, w_eco123429, w_eco123430, w_eco123431, w_eco123432, w_eco123433, w_eco123434, w_eco123435, w_eco123436, w_eco123437, w_eco123438, w_eco123439, w_eco123440, w_eco123441, w_eco123442, w_eco123443, w_eco123444, w_eco123445, w_eco123446, w_eco123447, w_eco123448, w_eco123449, w_eco123450, w_eco123451, w_eco123452, w_eco123453, w_eco123454, w_eco123455, w_eco123456, w_eco123457, w_eco123458, w_eco123459, w_eco123460, w_eco123461, w_eco123462, w_eco123463, w_eco123464, w_eco123465, w_eco123466, w_eco123467, w_eco123468, w_eco123469, w_eco123470, w_eco123471, w_eco123472, w_eco123473, w_eco123474, w_eco123475, w_eco123476, w_eco123477, w_eco123478, w_eco123479, w_eco123480, w_eco123481, w_eco123482, w_eco123483, w_eco123484, w_eco123485, w_eco123486, w_eco123487, w_eco123488, w_eco123489, w_eco123490, w_eco123491, w_eco123492, w_eco123493, w_eco123494, w_eco123495, w_eco123496, w_eco123497, w_eco123498, w_eco123499, w_eco123500, w_eco123501, w_eco123502, w_eco123503, w_eco123504, w_eco123505, w_eco123506, w_eco123507, w_eco123508, w_eco123509, w_eco123510, w_eco123511, w_eco123512, w_eco123513, w_eco123514, w_eco123515, w_eco123516, w_eco123517, w_eco123518, w_eco123519, w_eco123520, w_eco123521, w_eco123522, w_eco123523, w_eco123524, w_eco123525, w_eco123526, w_eco123527, w_eco123528, w_eco123529, w_eco123530, w_eco123531, w_eco123532, w_eco123533, w_eco123534, w_eco123535, w_eco123536, w_eco123537, w_eco123538, w_eco123539, w_eco123540, w_eco123541, w_eco123542, w_eco123543, w_eco123544, w_eco123545, w_eco123546, w_eco123547, w_eco123548, w_eco123549, w_eco123550, w_eco123551, w_eco123552, w_eco123553, w_eco123554, w_eco123555, w_eco123556, w_eco123557, w_eco123558, w_eco123559, w_eco123560, w_eco123561, w_eco123562, w_eco123563, w_eco123564, w_eco123565, w_eco123566, w_eco123567, w_eco123568, w_eco123569, w_eco123570, w_eco123571, w_eco123572, w_eco123573, w_eco123574, w_eco123575, w_eco123576, w_eco123577, w_eco123578, w_eco123579, w_eco123580, w_eco123581, w_eco123582, w_eco123583, w_eco123584, w_eco123585, w_eco123586, w_eco123587, w_eco123588, w_eco123589, w_eco123590, w_eco123591, w_eco123592, w_eco123593, w_eco123594, w_eco123595, w_eco123596, w_eco123597, w_eco123598, w_eco123599, w_eco123600, w_eco123601, w_eco123602, w_eco123603, w_eco123604, w_eco123605, w_eco123606, w_eco123607, w_eco123608, w_eco123609, w_eco123610, w_eco123611, w_eco123612, w_eco123613, w_eco123614, w_eco123615, w_eco123616, w_eco123617, w_eco123618, w_eco123619, w_eco123620, w_eco123621, w_eco123622, w_eco123623, w_eco123624, w_eco123625, w_eco123626, w_eco123627, w_eco123628, w_eco123629, w_eco123630, w_eco123631, w_eco123632, w_eco123633, w_eco123634, w_eco123635, w_eco123636, w_eco123637, w_eco123638, w_eco123639, w_eco123640, w_eco123641, w_eco123642, w_eco123643, w_eco123644, w_eco123645, w_eco123646, w_eco123647, w_eco123648, w_eco123649, w_eco123650, w_eco123651, w_eco123652, w_eco123653, w_eco123654, w_eco123655, w_eco123656, w_eco123657, w_eco123658, w_eco123659, w_eco123660, w_eco123661, w_eco123662, w_eco123663, w_eco123664, w_eco123665, w_eco123666, w_eco123667, w_eco123668, w_eco123669, w_eco123670, w_eco123671, w_eco123672, w_eco123673, w_eco123674, w_eco123675, w_eco123676, w_eco123677, w_eco123678, w_eco123679, w_eco123680, w_eco123681, w_eco123682, w_eco123683, w_eco123684, w_eco123685, w_eco123686, w_eco123687, w_eco123688, w_eco123689, w_eco123690, w_eco123691, w_eco123692, w_eco123693, w_eco123694, w_eco123695, w_eco123696, w_eco123697, w_eco123698, w_eco123699, w_eco123700, w_eco123701, w_eco123702, w_eco123703, w_eco123704, w_eco123705, w_eco123706, w_eco123707, w_eco123708, w_eco123709, w_eco123710, w_eco123711, w_eco123712, w_eco123713, w_eco123714, w_eco123715, w_eco123716, w_eco123717, w_eco123718, w_eco123719, w_eco123720, w_eco123721, w_eco123722, w_eco123723, w_eco123724, w_eco123725, w_eco123726, w_eco123727, w_eco123728, w_eco123729, w_eco123730, w_eco123731, w_eco123732, w_eco123733, w_eco123734, w_eco123735, w_eco123736, w_eco123737, w_eco123738, w_eco123739, w_eco123740, w_eco123741, w_eco123742, w_eco123743, w_eco123744, w_eco123745, w_eco123746, w_eco123747, w_eco123748, w_eco123749, w_eco123750, w_eco123751, w_eco123752, w_eco123753, w_eco123754, w_eco123755, w_eco123756, w_eco123757, w_eco123758, w_eco123759, w_eco123760, w_eco123761, w_eco123762, w_eco123763, w_eco123764, w_eco123765, w_eco123766, w_eco123767, w_eco123768, w_eco123769, w_eco123770, w_eco123771, w_eco123772, w_eco123773, w_eco123774, w_eco123775, w_eco123776, w_eco123777, w_eco123778, w_eco123779, w_eco123780, w_eco123781, w_eco123782, w_eco123783, w_eco123784, w_eco123785, w_eco123786, w_eco123787, w_eco123788, w_eco123789, w_eco123790, w_eco123791, w_eco123792, w_eco123793, w_eco123794, w_eco123795, w_eco123796, w_eco123797, w_eco123798, w_eco123799, w_eco123800, w_eco123801, w_eco123802, w_eco123803, w_eco123804, w_eco123805, w_eco123806, w_eco123807, w_eco123808, w_eco123809, w_eco123810, w_eco123811, w_eco123812, w_eco123813, w_eco123814, w_eco123815, w_eco123816, w_eco123817, w_eco123818, w_eco123819, w_eco123820, w_eco123821, w_eco123822, w_eco123823, w_eco123824, w_eco123825, w_eco123826, w_eco123827, w_eco123828, w_eco123829, w_eco123830, w_eco123831, w_eco123832, w_eco123833, w_eco123834, w_eco123835, w_eco123836, w_eco123837, w_eco123838, w_eco123839, w_eco123840, w_eco123841, w_eco123842, w_eco123843, w_eco123844, w_eco123845, w_eco123846, w_eco123847, w_eco123848, w_eco123849, w_eco123850, w_eco123851, w_eco123852, w_eco123853, w_eco123854, w_eco123855, w_eco123856, w_eco123857, w_eco123858, w_eco123859, w_eco123860, w_eco123861, w_eco123862, w_eco123863, w_eco123864, w_eco123865, w_eco123866, w_eco123867, w_eco123868, w_eco123869, w_eco123870, w_eco123871, w_eco123872, w_eco123873, w_eco123874, w_eco123875, w_eco123876, w_eco123877, w_eco123878, w_eco123879, w_eco123880, w_eco123881, w_eco123882, w_eco123883, w_eco123884, w_eco123885, w_eco123886, w_eco123887, w_eco123888, w_eco123889, w_eco123890, w_eco123891, w_eco123892, w_eco123893, w_eco123894, w_eco123895, w_eco123896, w_eco123897, w_eco123898, w_eco123899, w_eco123900, w_eco123901, w_eco123902, w_eco123903, w_eco123904, w_eco123905, w_eco123906, w_eco123907, w_eco123908, w_eco123909, w_eco123910, w_eco123911, w_eco123912, w_eco123913, w_eco123914, w_eco123915, w_eco123916, w_eco123917, w_eco123918, w_eco123919, w_eco123920, w_eco123921, w_eco123922, w_eco123923, w_eco123924, w_eco123925, w_eco123926, w_eco123927, w_eco123928, w_eco123929, w_eco123930, w_eco123931, w_eco123932, w_eco123933, w_eco123934, w_eco123935, w_eco123936, w_eco123937, w_eco123938, w_eco123939, w_eco123940, w_eco123941, w_eco123942, w_eco123943, w_eco123944, w_eco123945, w_eco123946, w_eco123947, w_eco123948, w_eco123949, w_eco123950, w_eco123951, w_eco123952, w_eco123953, w_eco123954, w_eco123955, w_eco123956, w_eco123957, w_eco123958, w_eco123959, w_eco123960, w_eco123961, w_eco123962, w_eco123963, w_eco123964, w_eco123965, w_eco123966, w_eco123967, w_eco123968, w_eco123969, w_eco123970, w_eco123971, w_eco123972, w_eco123973, w_eco123974, w_eco123975, w_eco123976, w_eco123977, w_eco123978, w_eco123979, w_eco123980, w_eco123981, w_eco123982, w_eco123983, w_eco123984, w_eco123985, w_eco123986, w_eco123987, w_eco123988, w_eco123989, w_eco123990, w_eco123991, w_eco123992, w_eco123993, w_eco123994, w_eco123995, w_eco123996, w_eco123997, w_eco123998, w_eco123999, w_eco124000, w_eco124001, w_eco124002, w_eco124003, w_eco124004, w_eco124005, w_eco124006, w_eco124007, w_eco124008, w_eco124009, w_eco124010, w_eco124011, w_eco124012, w_eco124013, w_eco124014, w_eco124015, w_eco124016, w_eco124017, w_eco124018, w_eco124019, w_eco124020, w_eco124021, w_eco124022, w_eco124023, w_eco124024, w_eco124025, w_eco124026, w_eco124027, w_eco124028, w_eco124029, w_eco124030, w_eco124031, w_eco124032, w_eco124033, w_eco124034, w_eco124035, w_eco124036, w_eco124037, w_eco124038, w_eco124039, w_eco124040, w_eco124041, w_eco124042, w_eco124043, w_eco124044, w_eco124045, w_eco124046, w_eco124047, w_eco124048, w_eco124049, w_eco124050, w_eco124051, w_eco124052, w_eco124053, w_eco124054, w_eco124055, w_eco124056, w_eco124057, w_eco124058, w_eco124059, w_eco124060, w_eco124061, w_eco124062, w_eco124063, w_eco124064, w_eco124065, w_eco124066, w_eco124067, w_eco124068, w_eco124069, w_eco124070, w_eco124071, w_eco124072, w_eco124073, w_eco124074, w_eco124075, w_eco124076, w_eco124077, w_eco124078, w_eco124079, w_eco124080, w_eco124081, w_eco124082, w_eco124083, w_eco124084, w_eco124085, w_eco124086, w_eco124087, w_eco124088, w_eco124089, w_eco124090, w_eco124091, w_eco124092, w_eco124093, w_eco124094, w_eco124095, w_eco124096, w_eco124097, w_eco124098, w_eco124099, w_eco124100, w_eco124101, w_eco124102, w_eco124103, w_eco124104, w_eco124105, w_eco124106, w_eco124107, w_eco124108, w_eco124109, w_eco124110, w_eco124111, w_eco124112, w_eco124113, w_eco124114, w_eco124115, w_eco124116, w_eco124117, w_eco124118, w_eco124119, w_eco124120, w_eco124121, w_eco124122, w_eco124123, w_eco124124, w_eco124125, w_eco124126, w_eco124127, w_eco124128, w_eco124129, w_eco124130, w_eco124131, w_eco124132, w_eco124133, w_eco124134, w_eco124135, w_eco124136, w_eco124137, w_eco124138, w_eco124139, w_eco124140, w_eco124141, w_eco124142, w_eco124143, w_eco124144, w_eco124145, w_eco124146, w_eco124147, w_eco124148, w_eco124149, w_eco124150, w_eco124151, w_eco124152, w_eco124153, w_eco124154, w_eco124155, w_eco124156, w_eco124157, w_eco124158, w_eco124159, w_eco124160, w_eco124161, w_eco124162, w_eco124163, w_eco124164, w_eco124165, w_eco124166, w_eco124167, w_eco124168, w_eco124169, w_eco124170, w_eco124171, w_eco124172, w_eco124173, w_eco124174, w_eco124175, w_eco124176, w_eco124177, w_eco124178, w_eco124179, w_eco124180, w_eco124181, w_eco124182, w_eco124183, w_eco124184, w_eco124185, w_eco124186, w_eco124187, w_eco124188, w_eco124189, w_eco124190, w_eco124191, w_eco124192, w_eco124193, w_eco124194, w_eco124195, w_eco124196, w_eco124197, w_eco124198, w_eco124199, w_eco124200, w_eco124201, w_eco124202, w_eco124203, w_eco124204, w_eco124205, w_eco124206, w_eco124207, w_eco124208, w_eco124209, w_eco124210, w_eco124211, w_eco124212, w_eco124213, w_eco124214, w_eco124215, w_eco124216, w_eco124217, w_eco124218, w_eco124219, w_eco124220, w_eco124221, w_eco124222, w_eco124223, w_eco124224, w_eco124225, w_eco124226, w_eco124227, w_eco124228, w_eco124229, w_eco124230, w_eco124231, w_eco124232, w_eco124233, w_eco124234, w_eco124235, w_eco124236, w_eco124237, w_eco124238, w_eco124239, w_eco124240, w_eco124241, w_eco124242, w_eco124243, w_eco124244, w_eco124245, w_eco124246, w_eco124247, w_eco124248, w_eco124249, w_eco124250, w_eco124251, w_eco124252, w_eco124253, w_eco124254, w_eco124255, w_eco124256, w_eco124257, w_eco124258, w_eco124259, w_eco124260, w_eco124261, w_eco124262, w_eco124263, w_eco124264, w_eco124265, w_eco124266, w_eco124267, w_eco124268, w_eco124269, w_eco124270, w_eco124271, w_eco124272, w_eco124273, w_eco124274, w_eco124275, w_eco124276, w_eco124277, w_eco124278, w_eco124279, w_eco124280, w_eco124281, w_eco124282, w_eco124283, w_eco124284, w_eco124285, w_eco124286, w_eco124287, w_eco124288, w_eco124289, w_eco124290, w_eco124291, w_eco124292, w_eco124293, w_eco124294, w_eco124295, w_eco124296, w_eco124297, w_eco124298, w_eco124299, w_eco124300, w_eco124301, w_eco124302, w_eco124303, w_eco124304, w_eco124305, w_eco124306, w_eco124307, w_eco124308, w_eco124309, w_eco124310, w_eco124311, w_eco124312, w_eco124313, w_eco124314, w_eco124315, w_eco124316, w_eco124317, w_eco124318, w_eco124319, w_eco124320, w_eco124321, w_eco124322, w_eco124323, w_eco124324, w_eco124325, w_eco124326, w_eco124327, w_eco124328, w_eco124329, w_eco124330, w_eco124331, w_eco124332, w_eco124333, w_eco124334, w_eco124335, w_eco124336, w_eco124337, w_eco124338, w_eco124339, w_eco124340, w_eco124341, w_eco124342, w_eco124343, w_eco124344, w_eco124345, w_eco124346, w_eco124347, w_eco124348, w_eco124349, w_eco124350, w_eco124351, w_eco124352, w_eco124353, w_eco124354, w_eco124355, w_eco124356, w_eco124357, w_eco124358, w_eco124359, w_eco124360, w_eco124361, w_eco124362, w_eco124363, w_eco124364, w_eco124365, w_eco124366, w_eco124367, w_eco124368, w_eco124369, w_eco124370, w_eco124371, w_eco124372, w_eco124373, w_eco124374, w_eco124375, w_eco124376, w_eco124377, w_eco124378, w_eco124379, w_eco124380, w_eco124381, w_eco124382, w_eco124383, w_eco124384, w_eco124385, w_eco124386, w_eco124387, w_eco124388, w_eco124389, w_eco124390, w_eco124391, w_eco124392, w_eco124393, w_eco124394, w_eco124395, w_eco124396, w_eco124397, w_eco124398, w_eco124399, w_eco124400, w_eco124401, w_eco124402, w_eco124403, w_eco124404, w_eco124405, w_eco124406, w_eco124407, w_eco124408, w_eco124409, w_eco124410, w_eco124411, w_eco124412, w_eco124413, w_eco124414, w_eco124415, w_eco124416, w_eco124417, w_eco124418, w_eco124419, w_eco124420, w_eco124421, w_eco124422, w_eco124423, w_eco124424, w_eco124425, w_eco124426, w_eco124427, w_eco124428, w_eco124429, w_eco124430, w_eco124431, w_eco124432, w_eco124433, w_eco124434, w_eco124435, w_eco124436, w_eco124437, w_eco124438, w_eco124439, w_eco124440, w_eco124441, w_eco124442, w_eco124443, w_eco124444, w_eco124445, w_eco124446, w_eco124447, w_eco124448, w_eco124449, w_eco124450, w_eco124451, w_eco124452, w_eco124453, w_eco124454, w_eco124455, w_eco124456, w_eco124457, w_eco124458, w_eco124459, w_eco124460, w_eco124461, w_eco124462, w_eco124463, w_eco124464, w_eco124465, w_eco124466, w_eco124467, w_eco124468, w_eco124469, w_eco124470, w_eco124471, w_eco124472, w_eco124473, w_eco124474, w_eco124475, w_eco124476, w_eco124477, w_eco124478, w_eco124479, w_eco124480, w_eco124481, w_eco124482, w_eco124483, w_eco124484, w_eco124485, w_eco124486, w_eco124487, w_eco124488, w_eco124489, w_eco124490, w_eco124491, w_eco124492, w_eco124493, w_eco124494, w_eco124495, w_eco124496, w_eco124497, w_eco124498, w_eco124499, w_eco124500, w_eco124501, w_eco124502, w_eco124503, w_eco124504, w_eco124505, w_eco124506, w_eco124507, w_eco124508, w_eco124509, w_eco124510, w_eco124511, w_eco124512, w_eco124513, w_eco124514, w_eco124515, w_eco124516, w_eco124517, w_eco124518, w_eco124519, w_eco124520, w_eco124521, w_eco124522, w_eco124523, w_eco124524, w_eco124525, w_eco124526, w_eco124527, w_eco124528, w_eco124529, w_eco124530, w_eco124531, w_eco124532, w_eco124533, w_eco124534, w_eco124535, w_eco124536, w_eco124537, w_eco124538, w_eco124539, w_eco124540, w_eco124541, w_eco124542, w_eco124543, w_eco124544, w_eco124545, w_eco124546, w_eco124547, w_eco124548, w_eco124549, w_eco124550, w_eco124551, w_eco124552, w_eco124553, w_eco124554, w_eco124555, w_eco124556, w_eco124557, w_eco124558, w_eco124559, w_eco124560, w_eco124561, w_eco124562, w_eco124563, w_eco124564, w_eco124565, w_eco124566, w_eco124567, w_eco124568, w_eco124569, w_eco124570, w_eco124571, w_eco124572, w_eco124573, w_eco124574, w_eco124575, w_eco124576, w_eco124577, w_eco124578, w_eco124579, w_eco124580, w_eco124581, w_eco124582, w_eco124583, w_eco124584, w_eco124585, w_eco124586, w_eco124587, w_eco124588, w_eco124589, w_eco124590, w_eco124591, w_eco124592, w_eco124593, w_eco124594, w_eco124595, w_eco124596, w_eco124597, w_eco124598, w_eco124599, w_eco124600, w_eco124601, w_eco124602, w_eco124603, w_eco124604, w_eco124605, w_eco124606, w_eco124607, w_eco124608, w_eco124609, w_eco124610, w_eco124611, w_eco124612, w_eco124613, w_eco124614, w_eco124615, w_eco124616, w_eco124617, w_eco124618, w_eco124619, w_eco124620, w_eco124621, w_eco124622, w_eco124623, w_eco124624, w_eco124625, w_eco124626, w_eco124627, w_eco124628, w_eco124629, w_eco124630, w_eco124631, w_eco124632, w_eco124633, w_eco124634, w_eco124635, w_eco124636, w_eco124637, w_eco124638, w_eco124639, w_eco124640, w_eco124641, w_eco124642, w_eco124643, w_eco124644, w_eco124645, w_eco124646, w_eco124647, w_eco124648, w_eco124649, w_eco124650, w_eco124651, w_eco124652, w_eco124653, w_eco124654, w_eco124655, w_eco124656, w_eco124657, w_eco124658, w_eco124659, w_eco124660, w_eco124661, w_eco124662, w_eco124663, w_eco124664, w_eco124665, w_eco124666, w_eco124667, w_eco124668, w_eco124669, w_eco124670, w_eco124671, w_eco124672, w_eco124673, w_eco124674, w_eco124675, w_eco124676, w_eco124677, w_eco124678, w_eco124679, w_eco124680, w_eco124681, w_eco124682, w_eco124683, w_eco124684, w_eco124685, w_eco124686, w_eco124687, w_eco124688, w_eco124689, w_eco124690, w_eco124691, w_eco124692, w_eco124693, w_eco124694, w_eco124695, w_eco124696, w_eco124697, w_eco124698, w_eco124699, w_eco124700, w_eco124701, w_eco124702, w_eco124703, w_eco124704, w_eco124705, w_eco124706, w_eco124707, w_eco124708, w_eco124709, w_eco124710, w_eco124711, w_eco124712, w_eco124713, w_eco124714, w_eco124715, w_eco124716, w_eco124717, w_eco124718, w_eco124719, w_eco124720, w_eco124721, w_eco124722, w_eco124723, w_eco124724, w_eco124725, w_eco124726, w_eco124727, w_eco124728, w_eco124729, w_eco124730, w_eco124731, w_eco124732, w_eco124733, w_eco124734, w_eco124735, w_eco124736, w_eco124737, w_eco124738, w_eco124739, w_eco124740, w_eco124741, w_eco124742, w_eco124743, w_eco124744, w_eco124745, w_eco124746, w_eco124747, w_eco124748, w_eco124749, w_eco124750, w_eco124751, w_eco124752, w_eco124753, w_eco124754, w_eco124755, w_eco124756, w_eco124757, w_eco124758, w_eco124759, w_eco124760, w_eco124761, w_eco124762, w_eco124763, w_eco124764, w_eco124765, w_eco124766, w_eco124767, w_eco124768, w_eco124769, w_eco124770, w_eco124771, w_eco124772, w_eco124773, w_eco124774, w_eco124775, w_eco124776, w_eco124777, w_eco124778, w_eco124779, w_eco124780, w_eco124781, w_eco124782, w_eco124783, w_eco124784, w_eco124785, w_eco124786, w_eco124787, w_eco124788, w_eco124789, w_eco124790, w_eco124791, w_eco124792, w_eco124793, w_eco124794, w_eco124795, w_eco124796, w_eco124797, w_eco124798, w_eco124799, w_eco124800, w_eco124801, w_eco124802, w_eco124803, w_eco124804, w_eco124805, w_eco124806, w_eco124807, w_eco124808, w_eco124809, w_eco124810, w_eco124811, w_eco124812, w_eco124813, w_eco124814, w_eco124815, w_eco124816, w_eco124817, w_eco124818, w_eco124819, w_eco124820, w_eco124821, w_eco124822, w_eco124823, w_eco124824, w_eco124825, w_eco124826, w_eco124827, w_eco124828, w_eco124829, w_eco124830, w_eco124831, w_eco124832, w_eco124833, w_eco124834, w_eco124835, w_eco124836, w_eco124837, w_eco124838, w_eco124839, w_eco124840, w_eco124841, w_eco124842, w_eco124843, w_eco124844, w_eco124845, w_eco124846, w_eco124847, w_eco124848, w_eco124849, w_eco124850, w_eco124851, w_eco124852, w_eco124853, w_eco124854, w_eco124855, w_eco124856, w_eco124857, w_eco124858, w_eco124859, w_eco124860, w_eco124861, w_eco124862, w_eco124863, w_eco124864, w_eco124865, w_eco124866, w_eco124867, w_eco124868, w_eco124869, w_eco124870, w_eco124871, w_eco124872, w_eco124873, w_eco124874, w_eco124875, w_eco124876, w_eco124877, w_eco124878, w_eco124879, w_eco124880, w_eco124881, w_eco124882, w_eco124883, w_eco124884, w_eco124885, w_eco124886, w_eco124887, w_eco124888, w_eco124889, w_eco124890, w_eco124891, w_eco124892, w_eco124893, w_eco124894, w_eco124895, w_eco124896, w_eco124897, w_eco124898, w_eco124899, w_eco124900, w_eco124901, w_eco124902, w_eco124903, w_eco124904, w_eco124905, w_eco124906, w_eco124907, w_eco124908, w_eco124909, w_eco124910, w_eco124911, w_eco124912, w_eco124913, w_eco124914, w_eco124915, w_eco124916, w_eco124917, w_eco124918, w_eco124919, w_eco124920, w_eco124921, w_eco124922, w_eco124923, w_eco124924, w_eco124925, w_eco124926, w_eco124927, w_eco124928, w_eco124929, w_eco124930, w_eco124931, w_eco124932, w_eco124933, w_eco124934, w_eco124935, w_eco124936, w_eco124937, w_eco124938, w_eco124939, w_eco124940, w_eco124941, w_eco124942, w_eco124943, w_eco124944, w_eco124945, w_eco124946, w_eco124947, w_eco124948, w_eco124949, w_eco124950, w_eco124951, w_eco124952, w_eco124953, w_eco124954, w_eco124955, w_eco124956, w_eco124957, w_eco124958, w_eco124959, w_eco124960, w_eco124961, w_eco124962, w_eco124963, w_eco124964, w_eco124965, w_eco124966, w_eco124967, w_eco124968, w_eco124969, w_eco124970, w_eco124971, w_eco124972, w_eco124973, w_eco124974, w_eco124975, w_eco124976, w_eco124977, w_eco124978, w_eco124979, w_eco124980, w_eco124981, w_eco124982, w_eco124983, w_eco124984, w_eco124985, w_eco124986, w_eco124987, w_eco124988, w_eco124989, w_eco124990, w_eco124991, w_eco124992, w_eco124993, w_eco124994, w_eco124995, w_eco124996, w_eco124997, w_eco124998, w_eco124999, w_eco125000, w_eco125001, w_eco125002, w_eco125003, w_eco125004, w_eco125005, w_eco125006, w_eco125007, w_eco125008, w_eco125009, w_eco125010, w_eco125011, w_eco125012, w_eco125013, w_eco125014, w_eco125015, w_eco125016, w_eco125017, w_eco125018, w_eco125019, w_eco125020, w_eco125021, w_eco125022, w_eco125023, w_eco125024, w_eco125025, w_eco125026, w_eco125027, w_eco125028, w_eco125029, w_eco125030, w_eco125031, w_eco125032, w_eco125033, w_eco125034, w_eco125035, w_eco125036, w_eco125037, w_eco125038, w_eco125039, w_eco125040, w_eco125041, w_eco125042, w_eco125043, w_eco125044, w_eco125045, w_eco125046, w_eco125047, w_eco125048, w_eco125049, w_eco125050, w_eco125051, w_eco125052, w_eco125053, w_eco125054, w_eco125055, w_eco125056, w_eco125057, w_eco125058, w_eco125059, w_eco125060, w_eco125061, w_eco125062, w_eco125063, w_eco125064, w_eco125065, w_eco125066, w_eco125067, w_eco125068, w_eco125069, w_eco125070, w_eco125071, w_eco125072, w_eco125073, w_eco125074, w_eco125075, w_eco125076, w_eco125077, w_eco125078, w_eco125079, w_eco125080, w_eco125081, w_eco125082, w_eco125083, w_eco125084, w_eco125085, w_eco125086, w_eco125087, w_eco125088, w_eco125089, w_eco125090, w_eco125091, w_eco125092, w_eco125093, w_eco125094, w_eco125095, w_eco125096, w_eco125097, w_eco125098, w_eco125099, w_eco125100, w_eco125101, w_eco125102, w_eco125103, w_eco125104, w_eco125105, w_eco125106, w_eco125107, w_eco125108, w_eco125109, w_eco125110, w_eco125111, w_eco125112, w_eco125113, w_eco125114, w_eco125115, w_eco125116, w_eco125117, w_eco125118, w_eco125119, w_eco125120, w_eco125121, w_eco125122, w_eco125123, w_eco125124, w_eco125125, w_eco125126, w_eco125127, w_eco125128, w_eco125129, w_eco125130, w_eco125131, w_eco125132, w_eco125133, w_eco125134, w_eco125135, w_eco125136, w_eco125137, w_eco125138, w_eco125139, w_eco125140, w_eco125141, w_eco125142, w_eco125143, w_eco125144, w_eco125145, w_eco125146, w_eco125147, w_eco125148, w_eco125149, w_eco125150, w_eco125151, w_eco125152, w_eco125153, w_eco125154, w_eco125155, w_eco125156, w_eco125157, w_eco125158, w_eco125159, w_eco125160, w_eco125161, w_eco125162, w_eco125163, w_eco125164, w_eco125165, w_eco125166, w_eco125167, w_eco125168, w_eco125169, w_eco125170, w_eco125171, w_eco125172, w_eco125173, w_eco125174, w_eco125175, w_eco125176, w_eco125177, w_eco125178, w_eco125179, w_eco125180, w_eco125181, w_eco125182, w_eco125183, w_eco125184, w_eco125185, w_eco125186, w_eco125187, w_eco125188, w_eco125189, w_eco125190, w_eco125191, w_eco125192, w_eco125193, w_eco125194, w_eco125195, w_eco125196, w_eco125197, w_eco125198, w_eco125199, w_eco125200, w_eco125201, w_eco125202, w_eco125203, w_eco125204, w_eco125205, w_eco125206, w_eco125207, w_eco125208, w_eco125209, w_eco125210, w_eco125211, w_eco125212, w_eco125213, w_eco125214, w_eco125215, w_eco125216, w_eco125217, w_eco125218, w_eco125219, w_eco125220, w_eco125221, w_eco125222, w_eco125223, w_eco125224, w_eco125225, w_eco125226, w_eco125227, w_eco125228, w_eco125229, w_eco125230, w_eco125231, w_eco125232, w_eco125233, w_eco125234, w_eco125235, w_eco125236, w_eco125237, w_eco125238, w_eco125239, w_eco125240, w_eco125241, w_eco125242, w_eco125243, w_eco125244, w_eco125245, w_eco125246, w_eco125247, w_eco125248, w_eco125249, w_eco125250, w_eco125251, w_eco125252, w_eco125253, w_eco125254, w_eco125255, w_eco125256, w_eco125257, w_eco125258, w_eco125259, w_eco125260, w_eco125261, w_eco125262, w_eco125263, w_eco125264, w_eco125265, w_eco125266, w_eco125267, w_eco125268, w_eco125269, w_eco125270, w_eco125271, w_eco125272, w_eco125273, w_eco125274, w_eco125275, w_eco125276, w_eco125277, w_eco125278, w_eco125279, w_eco125280, w_eco125281, w_eco125282, w_eco125283, w_eco125284, w_eco125285, w_eco125286, w_eco125287, w_eco125288, w_eco125289, w_eco125290, w_eco125291, w_eco125292, w_eco125293, w_eco125294, w_eco125295, w_eco125296, w_eco125297, w_eco125298, w_eco125299, w_eco125300, w_eco125301, w_eco125302, w_eco125303, w_eco125304, w_eco125305, w_eco125306, w_eco125307, w_eco125308, w_eco125309, w_eco125310, w_eco125311, w_eco125312, w_eco125313, w_eco125314, w_eco125315, w_eco125316, w_eco125317, w_eco125318, w_eco125319, w_eco125320, w_eco125321, w_eco125322, w_eco125323, w_eco125324, w_eco125325, w_eco125326, w_eco125327, w_eco125328, w_eco125329, w_eco125330, w_eco125331, w_eco125332, w_eco125333, w_eco125334, w_eco125335, w_eco125336, w_eco125337, w_eco125338, w_eco125339, w_eco125340, w_eco125341, w_eco125342, w_eco125343, w_eco125344, w_eco125345, w_eco125346, w_eco125347, w_eco125348, w_eco125349, w_eco125350, w_eco125351, w_eco125352, w_eco125353, w_eco125354, w_eco125355, w_eco125356, w_eco125357, w_eco125358, w_eco125359, w_eco125360, w_eco125361, w_eco125362, w_eco125363, w_eco125364, w_eco125365, w_eco125366, w_eco125367, w_eco125368, w_eco125369, w_eco125370, w_eco125371, w_eco125372, w_eco125373, w_eco125374, w_eco125375, w_eco125376, w_eco125377, w_eco125378, w_eco125379, w_eco125380, w_eco125381, w_eco125382, w_eco125383, w_eco125384, w_eco125385, w_eco125386, w_eco125387, w_eco125388, w_eco125389, w_eco125390, w_eco125391, w_eco125392, w_eco125393, w_eco125394, w_eco125395, w_eco125396, w_eco125397, w_eco125398, w_eco125399, w_eco125400, w_eco125401, w_eco125402, w_eco125403, w_eco125404, w_eco125405, w_eco125406, w_eco125407, w_eco125408, w_eco125409, w_eco125410, w_eco125411, w_eco125412, w_eco125413, w_eco125414, w_eco125415, w_eco125416, w_eco125417, w_eco125418, w_eco125419, w_eco125420, w_eco125421, w_eco125422, w_eco125423, w_eco125424, w_eco125425, w_eco125426, w_eco125427, w_eco125428, w_eco125429, w_eco125430, w_eco125431, w_eco125432, w_eco125433, w_eco125434, w_eco125435, w_eco125436, w_eco125437, w_eco125438, w_eco125439, w_eco125440, w_eco125441, w_eco125442, w_eco125443, w_eco125444, w_eco125445, w_eco125446, w_eco125447, w_eco125448, w_eco125449, w_eco125450, w_eco125451, w_eco125452, w_eco125453, w_eco125454, w_eco125455, w_eco125456, w_eco125457, w_eco125458, w_eco125459, w_eco125460, w_eco125461, w_eco125462, w_eco125463, w_eco125464, w_eco125465, w_eco125466, w_eco125467, w_eco125468, w_eco125469, w_eco125470, w_eco125471, w_eco125472, w_eco125473, w_eco125474, w_eco125475, w_eco125476, w_eco125477, w_eco125478, w_eco125479, w_eco125480, w_eco125481, w_eco125482, w_eco125483, w_eco125484, w_eco125485, w_eco125486, w_eco125487, w_eco125488, w_eco125489, w_eco125490, w_eco125491, w_eco125492, w_eco125493, w_eco125494, w_eco125495, w_eco125496, w_eco125497, w_eco125498, w_eco125499, w_eco125500, w_eco125501, w_eco125502, w_eco125503, w_eco125504, w_eco125505, w_eco125506, w_eco125507, w_eco125508, w_eco125509, w_eco125510, w_eco125511, w_eco125512, w_eco125513, w_eco125514, w_eco125515, w_eco125516, w_eco125517, w_eco125518, w_eco125519, w_eco125520, w_eco125521, w_eco125522, w_eco125523, w_eco125524, w_eco125525, w_eco125526, w_eco125527, w_eco125528, w_eco125529, w_eco125530, w_eco125531, w_eco125532, w_eco125533, w_eco125534, w_eco125535, w_eco125536, w_eco125537, w_eco125538, w_eco125539, w_eco125540, w_eco125541, w_eco125542, w_eco125543, w_eco125544, w_eco125545, w_eco125546, w_eco125547, w_eco125548, w_eco125549, w_eco125550, w_eco125551, w_eco125552, w_eco125553, w_eco125554, w_eco125555, w_eco125556, w_eco125557, w_eco125558, w_eco125559, w_eco125560, w_eco125561, w_eco125562, w_eco125563, w_eco125564, w_eco125565, w_eco125566, w_eco125567, w_eco125568, w_eco125569, w_eco125570, w_eco125571, w_eco125572, w_eco125573, w_eco125574, w_eco125575, w_eco125576, w_eco125577, w_eco125578, w_eco125579, w_eco125580, w_eco125581, w_eco125582, w_eco125583, w_eco125584, w_eco125585, w_eco125586, w_eco125587, w_eco125588, w_eco125589, w_eco125590, w_eco125591, w_eco125592, w_eco125593, w_eco125594, w_eco125595, w_eco125596, w_eco125597, w_eco125598, w_eco125599, w_eco125600, w_eco125601, w_eco125602, w_eco125603, w_eco125604, w_eco125605, w_eco125606, w_eco125607, w_eco125608, w_eco125609, w_eco125610, w_eco125611, w_eco125612, w_eco125613, w_eco125614, w_eco125615, w_eco125616, w_eco125617, w_eco125618, w_eco125619, w_eco125620, w_eco125621, w_eco125622, w_eco125623, w_eco125624, w_eco125625, w_eco125626, w_eco125627, w_eco125628, w_eco125629, w_eco125630, w_eco125631, w_eco125632, w_eco125633, w_eco125634, w_eco125635, w_eco125636, w_eco125637, w_eco125638, w_eco125639, w_eco125640, w_eco125641, w_eco125642, w_eco125643, w_eco125644, w_eco125645, w_eco125646, w_eco125647, w_eco125648, w_eco125649, w_eco125650, w_eco125651, w_eco125652, w_eco125653, w_eco125654, w_eco125655, w_eco125656, w_eco125657, w_eco125658, w_eco125659, w_eco125660, w_eco125661, w_eco125662, w_eco125663, w_eco125664, w_eco125665, w_eco125666, w_eco125667, w_eco125668, w_eco125669, w_eco125670, w_eco125671, w_eco125672, w_eco125673, w_eco125674, w_eco125675, w_eco125676, w_eco125677, w_eco125678, w_eco125679, w_eco125680, w_eco125681, w_eco125682, w_eco125683, w_eco125684, w_eco125685, w_eco125686, w_eco125687, w_eco125688, w_eco125689, w_eco125690, w_eco125691, w_eco125692, w_eco125693, w_eco125694, w_eco125695, w_eco125696, w_eco125697, w_eco125698, w_eco125699, w_eco125700, w_eco125701, w_eco125702, w_eco125703, w_eco125704, w_eco125705, w_eco125706, w_eco125707, w_eco125708, w_eco125709, w_eco125710, w_eco125711, w_eco125712, w_eco125713, w_eco125714, w_eco125715, w_eco125716, w_eco125717, w_eco125718, w_eco125719, w_eco125720, w_eco125721, w_eco125722, w_eco125723, w_eco125724, w_eco125725, w_eco125726, w_eco125727, w_eco125728, w_eco125729, w_eco125730, w_eco125731, w_eco125732, w_eco125733, w_eco125734, w_eco125735, w_eco125736, w_eco125737, w_eco125738, w_eco125739, w_eco125740, w_eco125741, w_eco125742, w_eco125743, w_eco125744, w_eco125745, w_eco125746, w_eco125747, w_eco125748, w_eco125749, w_eco125750, w_eco125751, w_eco125752, w_eco125753, w_eco125754, w_eco125755, w_eco125756, w_eco125757, w_eco125758, w_eco125759, w_eco125760, w_eco125761, w_eco125762, w_eco125763, w_eco125764, w_eco125765, w_eco125766, w_eco125767, w_eco125768, w_eco125769, w_eco125770, w_eco125771, w_eco125772, w_eco125773, w_eco125774, w_eco125775, w_eco125776, w_eco125777, w_eco125778, w_eco125779, w_eco125780, w_eco125781, w_eco125782, w_eco125783, w_eco125784, w_eco125785, w_eco125786, w_eco125787, w_eco125788, w_eco125789, w_eco125790, w_eco125791, w_eco125792, w_eco125793, w_eco125794, w_eco125795, w_eco125796, w_eco125797, w_eco125798, w_eco125799, w_eco125800, w_eco125801, w_eco125802, w_eco125803, w_eco125804, w_eco125805, w_eco125806, w_eco125807, w_eco125808, w_eco125809, w_eco125810, w_eco125811, w_eco125812, w_eco125813, w_eco125814, w_eco125815, w_eco125816, w_eco125817, w_eco125818, w_eco125819, w_eco125820, w_eco125821, w_eco125822, w_eco125823, w_eco125824, w_eco125825, w_eco125826, w_eco125827, w_eco125828, w_eco125829, w_eco125830, w_eco125831, w_eco125832, w_eco125833, w_eco125834, w_eco125835, w_eco125836, w_eco125837, w_eco125838, w_eco125839, w_eco125840, w_eco125841, w_eco125842, w_eco125843, w_eco125844, w_eco125845, w_eco125846, w_eco125847, w_eco125848, w_eco125849, w_eco125850, w_eco125851, w_eco125852, w_eco125853, w_eco125854, w_eco125855, w_eco125856, w_eco125857, w_eco125858, w_eco125859, w_eco125860, w_eco125861, w_eco125862, w_eco125863, w_eco125864, w_eco125865, w_eco125866, w_eco125867, w_eco125868, w_eco125869, w_eco125870, w_eco125871, w_eco125872, w_eco125873, w_eco125874, w_eco125875, w_eco125876, w_eco125877, w_eco125878, w_eco125879, w_eco125880, w_eco125881, w_eco125882, w_eco125883, w_eco125884, w_eco125885, w_eco125886, w_eco125887, w_eco125888, w_eco125889, w_eco125890, w_eco125891, w_eco125892, w_eco125893, w_eco125894, w_eco125895, w_eco125896, w_eco125897, w_eco125898, w_eco125899, w_eco125900, w_eco125901, w_eco125902, w_eco125903, w_eco125904, w_eco125905, w_eco125906, w_eco125907, w_eco125908, w_eco125909, w_eco125910, w_eco125911, w_eco125912, w_eco125913, w_eco125914, w_eco125915, w_eco125916, w_eco125917, w_eco125918, w_eco125919, w_eco125920, w_eco125921, w_eco125922, w_eco125923, w_eco125924, w_eco125925, w_eco125926, w_eco125927, w_eco125928, w_eco125929, w_eco125930, w_eco125931, w_eco125932, w_eco125933, w_eco125934, w_eco125935, w_eco125936, w_eco125937, w_eco125938, w_eco125939, w_eco125940, w_eco125941, w_eco125942, w_eco125943, w_eco125944, w_eco125945, w_eco125946, w_eco125947, w_eco125948, w_eco125949, w_eco125950, w_eco125951, w_eco125952, w_eco125953, w_eco125954, w_eco125955, w_eco125956, w_eco125957, w_eco125958, w_eco125959, w_eco125960, w_eco125961, w_eco125962, w_eco125963, w_eco125964, w_eco125965, w_eco125966, w_eco125967, w_eco125968, w_eco125969, w_eco125970, w_eco125971, w_eco125972, w_eco125973, w_eco125974, w_eco125975, w_eco125976, w_eco125977, w_eco125978, w_eco125979, w_eco125980, w_eco125981, w_eco125982, w_eco125983, w_eco125984, w_eco125985, w_eco125986, w_eco125987, w_eco125988, w_eco125989, w_eco125990, w_eco125991, w_eco125992, w_eco125993, w_eco125994, w_eco125995, w_eco125996, w_eco125997, w_eco125998, w_eco125999, w_eco126000, w_eco126001, w_eco126002, w_eco126003, w_eco126004, w_eco126005, w_eco126006, w_eco126007, w_eco126008, w_eco126009, w_eco126010, w_eco126011, w_eco126012, w_eco126013, w_eco126014, w_eco126015, w_eco126016, w_eco126017, w_eco126018, w_eco126019, w_eco126020, w_eco126021, w_eco126022, w_eco126023, w_eco126024, w_eco126025, w_eco126026, w_eco126027, w_eco126028, w_eco126029, w_eco126030, w_eco126031, w_eco126032, w_eco126033, w_eco126034, w_eco126035, w_eco126036, w_eco126037, w_eco126038, w_eco126039, w_eco126040, w_eco126041, w_eco126042, w_eco126043, w_eco126044, w_eco126045, w_eco126046, w_eco126047, w_eco126048, w_eco126049, w_eco126050, w_eco126051, w_eco126052, w_eco126053, w_eco126054, w_eco126055, w_eco126056, w_eco126057, w_eco126058, w_eco126059, w_eco126060, w_eco126061, w_eco126062, w_eco126063, w_eco126064, w_eco126065, w_eco126066, w_eco126067, w_eco126068, w_eco126069, w_eco126070, w_eco126071, w_eco126072, w_eco126073, w_eco126074, w_eco126075, w_eco126076, w_eco126077, w_eco126078, w_eco126079, w_eco126080, w_eco126081, w_eco126082, w_eco126083, w_eco126084, w_eco126085, w_eco126086, w_eco126087, w_eco126088, w_eco126089, w_eco126090, w_eco126091, w_eco126092, w_eco126093, w_eco126094, w_eco126095, w_eco126096, w_eco126097, w_eco126098, w_eco126099, w_eco126100, w_eco126101, w_eco126102, w_eco126103, w_eco126104, w_eco126105, w_eco126106, w_eco126107, w_eco126108, w_eco126109, w_eco126110, w_eco126111, w_eco126112, w_eco126113, w_eco126114, w_eco126115, w_eco126116, w_eco126117, w_eco126118, w_eco126119, w_eco126120, w_eco126121, w_eco126122, w_eco126123, w_eco126124, w_eco126125, w_eco126126, w_eco126127, w_eco126128, w_eco126129, w_eco126130, w_eco126131, w_eco126132, w_eco126133, w_eco126134, w_eco126135, w_eco126136, w_eco126137, w_eco126138, w_eco126139, w_eco126140, w_eco126141, w_eco126142, w_eco126143, w_eco126144, w_eco126145, w_eco126146, w_eco126147, w_eco126148, w_eco126149, w_eco126150, w_eco126151, w_eco126152, w_eco126153, w_eco126154, w_eco126155, w_eco126156, w_eco126157, w_eco126158, w_eco126159, w_eco126160, w_eco126161, w_eco126162, w_eco126163, w_eco126164, w_eco126165, w_eco126166, w_eco126167, w_eco126168, w_eco126169, w_eco126170, w_eco126171, w_eco126172, w_eco126173, w_eco126174, w_eco126175, w_eco126176, w_eco126177, w_eco126178, w_eco126179, w_eco126180, w_eco126181, w_eco126182, w_eco126183, w_eco126184, w_eco126185, w_eco126186, w_eco126187, w_eco126188, w_eco126189, w_eco126190, w_eco126191, w_eco126192, w_eco126193, w_eco126194, w_eco126195, w_eco126196, w_eco126197, w_eco126198, w_eco126199, w_eco126200, w_eco126201, w_eco126202, w_eco126203, w_eco126204, w_eco126205, w_eco126206, w_eco126207, w_eco126208, w_eco126209, w_eco126210, w_eco126211, w_eco126212, w_eco126213, w_eco126214, w_eco126215, w_eco126216, w_eco126217, w_eco126218, w_eco126219, w_eco126220, w_eco126221, w_eco126222, w_eco126223, w_eco126224, w_eco126225, w_eco126226, w_eco126227, w_eco126228, w_eco126229, w_eco126230, w_eco126231, w_eco126232, w_eco126233, w_eco126234, w_eco126235, w_eco126236, w_eco126237, w_eco126238, w_eco126239, w_eco126240, w_eco126241, w_eco126242, w_eco126243, w_eco126244, w_eco126245, w_eco126246, w_eco126247, w_eco126248, w_eco126249, w_eco126250, w_eco126251, w_eco126252, w_eco126253, w_eco126254, w_eco126255, w_eco126256, w_eco126257, w_eco126258, w_eco126259, w_eco126260, w_eco126261, w_eco126262, w_eco126263, w_eco126264, w_eco126265, w_eco126266, w_eco126267, w_eco126268, w_eco126269, w_eco126270, w_eco126271, w_eco126272, w_eco126273, w_eco126274, w_eco126275, w_eco126276, w_eco126277, w_eco126278, w_eco126279, w_eco126280, w_eco126281, w_eco126282, w_eco126283, w_eco126284, w_eco126285, w_eco126286, w_eco126287, w_eco126288, w_eco126289, w_eco126290, w_eco126291, w_eco126292, w_eco126293, w_eco126294, w_eco126295, w_eco126296, w_eco126297, w_eco126298, w_eco126299, w_eco126300, w_eco126301, w_eco126302, w_eco126303, w_eco126304, w_eco126305, w_eco126306, w_eco126307, w_eco126308, w_eco126309, w_eco126310, w_eco126311, w_eco126312, w_eco126313, w_eco126314, w_eco126315, w_eco126316, w_eco126317, w_eco126318, w_eco126319, w_eco126320, w_eco126321, w_eco126322, w_eco126323, w_eco126324, w_eco126325, w_eco126326, w_eco126327, w_eco126328, w_eco126329, w_eco126330, w_eco126331, w_eco126332, w_eco126333, w_eco126334, w_eco126335, w_eco126336, w_eco126337, w_eco126338, w_eco126339, w_eco126340, w_eco126341, w_eco126342, w_eco126343, w_eco126344, w_eco126345, w_eco126346, w_eco126347, w_eco126348, w_eco126349, w_eco126350, w_eco126351, w_eco126352, w_eco126353, w_eco126354, w_eco126355, w_eco126356, w_eco126357, w_eco126358, w_eco126359, w_eco126360, w_eco126361, w_eco126362, w_eco126363, w_eco126364, w_eco126365, w_eco126366, w_eco126367, w_eco126368, w_eco126369, w_eco126370, w_eco126371, w_eco126372, w_eco126373, w_eco126374, w_eco126375, w_eco126376, w_eco126377, w_eco126378, w_eco126379, w_eco126380, w_eco126381, w_eco126382, w_eco126383, w_eco126384, w_eco126385, w_eco126386, w_eco126387, w_eco126388, w_eco126389, w_eco126390, w_eco126391, w_eco126392, w_eco126393, w_eco126394, w_eco126395, w_eco126396, w_eco126397, w_eco126398, w_eco126399, w_eco126400, w_eco126401, w_eco126402, w_eco126403, w_eco126404, w_eco126405, w_eco126406, w_eco126407, w_eco126408, w_eco126409, w_eco126410, w_eco126411, w_eco126412, w_eco126413, w_eco126414, w_eco126415, w_eco126416, w_eco126417, w_eco126418, w_eco126419, w_eco126420, w_eco126421, w_eco126422, w_eco126423, w_eco126424, w_eco126425, w_eco126426, w_eco126427, w_eco126428, w_eco126429, w_eco126430, w_eco126431, w_eco126432, w_eco126433, w_eco126434, w_eco126435, w_eco126436, w_eco126437, w_eco126438, w_eco126439, w_eco126440, w_eco126441, w_eco126442, w_eco126443, w_eco126444, w_eco126445, w_eco126446, w_eco126447, w_eco126448, w_eco126449, w_eco126450, w_eco126451, w_eco126452, w_eco126453, w_eco126454, w_eco126455, w_eco126456, w_eco126457, w_eco126458, w_eco126459, w_eco126460, w_eco126461, w_eco126462, w_eco126463, w_eco126464, w_eco126465, w_eco126466, w_eco126467, w_eco126468, w_eco126469, w_eco126470, w_eco126471, w_eco126472, w_eco126473, w_eco126474, w_eco126475, w_eco126476, w_eco126477, w_eco126478, w_eco126479, w_eco126480, w_eco126481, w_eco126482, w_eco126483, w_eco126484, w_eco126485, w_eco126486, w_eco126487, w_eco126488, w_eco126489, w_eco126490, w_eco126491, w_eco126492, w_eco126493, w_eco126494, w_eco126495, w_eco126496, w_eco126497, w_eco126498, w_eco126499, w_eco126500, w_eco126501, w_eco126502, w_eco126503, w_eco126504, w_eco126505, w_eco126506, w_eco126507, w_eco126508, w_eco126509, w_eco126510, w_eco126511, w_eco126512, w_eco126513, w_eco126514, w_eco126515, w_eco126516, w_eco126517, w_eco126518, w_eco126519, w_eco126520, w_eco126521, w_eco126522, w_eco126523, w_eco126524, w_eco126525, w_eco126526, w_eco126527, w_eco126528, w_eco126529, w_eco126530, w_eco126531, w_eco126532, w_eco126533, w_eco126534, w_eco126535, w_eco126536, w_eco126537, w_eco126538, w_eco126539, w_eco126540, w_eco126541, w_eco126542, w_eco126543, w_eco126544, w_eco126545, w_eco126546, w_eco126547, w_eco126548, w_eco126549, w_eco126550, w_eco126551, w_eco126552, w_eco126553, w_eco126554, w_eco126555, w_eco126556, w_eco126557, w_eco126558, w_eco126559, w_eco126560, w_eco126561, w_eco126562, w_eco126563, w_eco126564, w_eco126565, w_eco126566, w_eco126567, w_eco126568, w_eco126569, w_eco126570, w_eco126571, w_eco126572, w_eco126573, w_eco126574, w_eco126575, w_eco126576, w_eco126577, w_eco126578, w_eco126579, w_eco126580, w_eco126581, w_eco126582, w_eco126583, w_eco126584, w_eco126585, w_eco126586, w_eco126587, w_eco126588, w_eco126589, w_eco126590, w_eco126591, w_eco126592, w_eco126593, w_eco126594, w_eco126595, w_eco126596, w_eco126597, w_eco126598, w_eco126599, w_eco126600, w_eco126601, w_eco126602, w_eco126603, w_eco126604, w_eco126605, w_eco126606, w_eco126607, w_eco126608, w_eco126609, w_eco126610, w_eco126611, w_eco126612, w_eco126613, w_eco126614, w_eco126615, w_eco126616, w_eco126617, w_eco126618, w_eco126619, w_eco126620, w_eco126621, w_eco126622, w_eco126623, w_eco126624, w_eco126625, w_eco126626, w_eco126627, w_eco126628, w_eco126629, w_eco126630, w_eco126631, w_eco126632, w_eco126633, w_eco126634, w_eco126635, w_eco126636, w_eco126637, w_eco126638, w_eco126639, w_eco126640, w_eco126641, w_eco126642, w_eco126643, w_eco126644, w_eco126645, w_eco126646, w_eco126647, w_eco126648, w_eco126649, w_eco126650, w_eco126651, w_eco126652, w_eco126653, w_eco126654, w_eco126655, w_eco126656, w_eco126657, w_eco126658, w_eco126659, w_eco126660, w_eco126661, w_eco126662, w_eco126663, w_eco126664, w_eco126665, w_eco126666, w_eco126667, w_eco126668, w_eco126669, w_eco126670, w_eco126671, w_eco126672, w_eco126673, w_eco126674, w_eco126675, w_eco126676, w_eco126677, w_eco126678, w_eco126679, w_eco126680, w_eco126681, w_eco126682, w_eco126683, w_eco126684, w_eco126685, w_eco126686, w_eco126687, w_eco126688, w_eco126689, w_eco126690, w_eco126691, w_eco126692, w_eco126693, w_eco126694, w_eco126695, w_eco126696, w_eco126697, w_eco126698, w_eco126699, w_eco126700, w_eco126701, w_eco126702, w_eco126703, w_eco126704, w_eco126705, w_eco126706, w_eco126707, w_eco126708, w_eco126709, w_eco126710, w_eco126711, w_eco126712, w_eco126713, w_eco126714, w_eco126715, w_eco126716, w_eco126717, w_eco126718, w_eco126719, w_eco126720, w_eco126721, w_eco126722, w_eco126723, w_eco126724, w_eco126725, w_eco126726, w_eco126727, w_eco126728, w_eco126729, w_eco126730, w_eco126731, w_eco126732, w_eco126733, w_eco126734, w_eco126735, w_eco126736, w_eco126737, w_eco126738, w_eco126739, w_eco126740, w_eco126741, w_eco126742, w_eco126743, w_eco126744, w_eco126745, w_eco126746, w_eco126747, w_eco126748, w_eco126749, w_eco126750, w_eco126751, w_eco126752, w_eco126753, w_eco126754, w_eco126755, w_eco126756, w_eco126757, w_eco126758, w_eco126759, w_eco126760, w_eco126761, w_eco126762, w_eco126763, w_eco126764, w_eco126765, w_eco126766, w_eco126767, w_eco126768, w_eco126769, w_eco126770, w_eco126771, w_eco126772, w_eco126773, w_eco126774, w_eco126775, w_eco126776, w_eco126777, w_eco126778, w_eco126779, w_eco126780, w_eco126781, w_eco126782, w_eco126783, w_eco126784, w_eco126785, w_eco126786, w_eco126787, w_eco126788, w_eco126789, w_eco126790, w_eco126791, w_eco126792, w_eco126793, w_eco126794, w_eco126795, w_eco126796, w_eco126797, w_eco126798, w_eco126799, w_eco126800, w_eco126801, w_eco126802, w_eco126803, w_eco126804, w_eco126805, w_eco126806, w_eco126807, w_eco126808, w_eco126809, w_eco126810, w_eco126811, w_eco126812, w_eco126813, w_eco126814, w_eco126815, w_eco126816, w_eco126817, w_eco126818, w_eco126819, w_eco126820, w_eco126821, w_eco126822, w_eco126823, w_eco126824, w_eco126825, w_eco126826, w_eco126827, w_eco126828, w_eco126829, w_eco126830, w_eco126831, w_eco126832, w_eco126833, w_eco126834, w_eco126835, w_eco126836, w_eco126837, w_eco126838, w_eco126839, w_eco126840, w_eco126841, w_eco126842, w_eco126843, w_eco126844, w_eco126845, w_eco126846, w_eco126847, w_eco126848, w_eco126849, w_eco126850, w_eco126851, w_eco126852, w_eco126853, w_eco126854, w_eco126855, w_eco126856, w_eco126857, w_eco126858, w_eco126859, w_eco126860, w_eco126861, w_eco126862, w_eco126863, w_eco126864, w_eco126865, w_eco126866, w_eco126867, w_eco126868, w_eco126869, w_eco126870, w_eco126871, w_eco126872, w_eco126873, w_eco126874, w_eco126875, w_eco126876, w_eco126877, w_eco126878, w_eco126879, w_eco126880, w_eco126881, w_eco126882, w_eco126883, w_eco126884, w_eco126885, w_eco126886, w_eco126887, w_eco126888, w_eco126889, w_eco126890, w_eco126891, w_eco126892, w_eco126893, w_eco126894, w_eco126895, w_eco126896, w_eco126897, w_eco126898, w_eco126899, w_eco126900, w_eco126901, w_eco126902, w_eco126903, w_eco126904, w_eco126905, w_eco126906, w_eco126907, w_eco126908, w_eco126909, w_eco126910, w_eco126911, w_eco126912, w_eco126913, w_eco126914, w_eco126915, w_eco126916, w_eco126917, w_eco126918, w_eco126919, w_eco126920, w_eco126921, w_eco126922, w_eco126923, w_eco126924, w_eco126925, w_eco126926, w_eco126927, w_eco126928, w_eco126929, w_eco126930, w_eco126931, w_eco126932, w_eco126933, w_eco126934, w_eco126935, w_eco126936, w_eco126937, w_eco126938, w_eco126939, w_eco126940, w_eco126941, w_eco126942, w_eco126943, w_eco126944, w_eco126945, w_eco126946, w_eco126947, w_eco126948, w_eco126949, w_eco126950, w_eco126951, w_eco126952, w_eco126953, w_eco126954, w_eco126955, w_eco126956, w_eco126957, w_eco126958, w_eco126959, w_eco126960, w_eco126961, w_eco126962, w_eco126963, w_eco126964, w_eco126965, w_eco126966, w_eco126967, w_eco126968, w_eco126969, w_eco126970, w_eco126971, w_eco126972, w_eco126973, w_eco126974, w_eco126975, w_eco126976, w_eco126977, w_eco126978, w_eco126979, w_eco126980, w_eco126981, w_eco126982, w_eco126983, w_eco126984, w_eco126985, w_eco126986, w_eco126987, w_eco126988, w_eco126989, w_eco126990, w_eco126991, w_eco126992, w_eco126993, w_eco126994, w_eco126995, w_eco126996, w_eco126997, w_eco126998, w_eco126999, w_eco127000, w_eco127001, w_eco127002, w_eco127003, w_eco127004, w_eco127005, w_eco127006, w_eco127007, w_eco127008, w_eco127009, w_eco127010, w_eco127011, w_eco127012, w_eco127013, w_eco127014, w_eco127015, w_eco127016, w_eco127017, w_eco127018, w_eco127019, w_eco127020, w_eco127021, w_eco127022, w_eco127023, w_eco127024, w_eco127025, w_eco127026, w_eco127027, w_eco127028, w_eco127029, w_eco127030, w_eco127031, w_eco127032, w_eco127033, w_eco127034, w_eco127035, w_eco127036, w_eco127037, w_eco127038, w_eco127039, w_eco127040, w_eco127041, w_eco127042, w_eco127043, w_eco127044, w_eco127045, w_eco127046, w_eco127047, w_eco127048, w_eco127049, w_eco127050, w_eco127051, w_eco127052, w_eco127053, w_eco127054, w_eco127055, w_eco127056, w_eco127057, w_eco127058, w_eco127059, w_eco127060, w_eco127061, w_eco127062, w_eco127063, w_eco127064, w_eco127065, w_eco127066, w_eco127067, w_eco127068, w_eco127069, w_eco127070, w_eco127071, w_eco127072, w_eco127073, w_eco127074, w_eco127075, w_eco127076, w_eco127077, w_eco127078, w_eco127079, w_eco127080, w_eco127081, w_eco127082, w_eco127083, w_eco127084, w_eco127085, w_eco127086, w_eco127087, w_eco127088, w_eco127089, w_eco127090, w_eco127091, w_eco127092, w_eco127093, w_eco127094, w_eco127095, w_eco127096, w_eco127097, w_eco127098, w_eco127099, w_eco127100, w_eco127101, w_eco127102, w_eco127103, w_eco127104, w_eco127105, w_eco127106, w_eco127107, w_eco127108, w_eco127109, w_eco127110, w_eco127111, w_eco127112, w_eco127113, w_eco127114, w_eco127115, w_eco127116, w_eco127117, w_eco127118, w_eco127119, w_eco127120, w_eco127121, w_eco127122, w_eco127123, w_eco127124, w_eco127125, w_eco127126, w_eco127127, w_eco127128, w_eco127129, w_eco127130, w_eco127131, w_eco127132, w_eco127133, w_eco127134, w_eco127135, w_eco127136, w_eco127137, w_eco127138, w_eco127139, w_eco127140, w_eco127141, w_eco127142, w_eco127143, w_eco127144, w_eco127145, w_eco127146, w_eco127147, w_eco127148, w_eco127149, w_eco127150, w_eco127151, w_eco127152, w_eco127153, w_eco127154, w_eco127155, w_eco127156, w_eco127157, w_eco127158, w_eco127159, w_eco127160, w_eco127161, w_eco127162, w_eco127163, w_eco127164, w_eco127165, w_eco127166, w_eco127167, w_eco127168, w_eco127169, w_eco127170, w_eco127171, w_eco127172, w_eco127173, w_eco127174, w_eco127175, w_eco127176, w_eco127177, w_eco127178, w_eco127179, w_eco127180, w_eco127181, w_eco127182, w_eco127183, w_eco127184, w_eco127185, w_eco127186, w_eco127187, w_eco127188, w_eco127189, w_eco127190, w_eco127191, w_eco127192, w_eco127193, w_eco127194, w_eco127195, w_eco127196, w_eco127197, w_eco127198, w_eco127199, w_eco127200, w_eco127201, w_eco127202, w_eco127203, w_eco127204, w_eco127205, w_eco127206, w_eco127207, w_eco127208, w_eco127209, w_eco127210, w_eco127211, w_eco127212, w_eco127213, w_eco127214, w_eco127215, w_eco127216, w_eco127217, w_eco127218, w_eco127219, w_eco127220, w_eco127221, w_eco127222, w_eco127223, w_eco127224, w_eco127225, w_eco127226, w_eco127227, w_eco127228, w_eco127229, w_eco127230, w_eco127231, w_eco127232, w_eco127233, w_eco127234, w_eco127235, w_eco127236, w_eco127237, w_eco127238, w_eco127239, w_eco127240, w_eco127241, w_eco127242, w_eco127243, w_eco127244, w_eco127245, w_eco127246, w_eco127247, w_eco127248, w_eco127249, w_eco127250, w_eco127251, w_eco127252, w_eco127253, w_eco127254, w_eco127255, w_eco127256, w_eco127257, w_eco127258, w_eco127259, w_eco127260, w_eco127261, w_eco127262, w_eco127263, w_eco127264, w_eco127265, w_eco127266, w_eco127267, w_eco127268, w_eco127269, w_eco127270, w_eco127271, w_eco127272, w_eco127273, w_eco127274, w_eco127275, w_eco127276, w_eco127277, w_eco127278, w_eco127279, w_eco127280, w_eco127281, w_eco127282, w_eco127283, w_eco127284, w_eco127285, w_eco127286, w_eco127287, w_eco127288, w_eco127289, w_eco127290, w_eco127291, w_eco127292, w_eco127293, w_eco127294, w_eco127295, w_eco127296, w_eco127297, w_eco127298, w_eco127299, w_eco127300, w_eco127301, w_eco127302, w_eco127303, w_eco127304, w_eco127305, w_eco127306, w_eco127307, w_eco127308, w_eco127309, w_eco127310, w_eco127311, w_eco127312, w_eco127313, w_eco127314, w_eco127315, w_eco127316, w_eco127317, w_eco127318, w_eco127319, w_eco127320, w_eco127321, w_eco127322, w_eco127323, w_eco127324, w_eco127325, w_eco127326, w_eco127327, w_eco127328, w_eco127329, w_eco127330, w_eco127331, w_eco127332, w_eco127333, w_eco127334, w_eco127335, w_eco127336, w_eco127337, w_eco127338, w_eco127339, w_eco127340, w_eco127341, w_eco127342, w_eco127343, w_eco127344, w_eco127345, w_eco127346, w_eco127347, w_eco127348, w_eco127349, w_eco127350, w_eco127351, w_eco127352, w_eco127353, w_eco127354, w_eco127355, w_eco127356, w_eco127357, w_eco127358, w_eco127359, w_eco127360, w_eco127361, w_eco127362, w_eco127363, w_eco127364, w_eco127365, w_eco127366, w_eco127367, w_eco127368, w_eco127369, w_eco127370, w_eco127371, w_eco127372, w_eco127373, w_eco127374, w_eco127375, w_eco127376, w_eco127377, w_eco127378, w_eco127379, w_eco127380, w_eco127381, w_eco127382, w_eco127383, w_eco127384, w_eco127385, w_eco127386, w_eco127387, w_eco127388, w_eco127389, w_eco127390, w_eco127391, w_eco127392, w_eco127393, w_eco127394, w_eco127395, w_eco127396, w_eco127397, w_eco127398, w_eco127399, w_eco127400, w_eco127401, w_eco127402, w_eco127403, w_eco127404, w_eco127405, w_eco127406, w_eco127407, w_eco127408, w_eco127409, w_eco127410, w_eco127411, w_eco127412, w_eco127413, w_eco127414, w_eco127415, w_eco127416, w_eco127417, w_eco127418, w_eco127419, w_eco127420, w_eco127421, w_eco127422, w_eco127423, w_eco127424, w_eco127425, w_eco127426, w_eco127427, w_eco127428, w_eco127429, w_eco127430, w_eco127431, w_eco127432, w_eco127433, w_eco127434, w_eco127435, w_eco127436, w_eco127437, w_eco127438, w_eco127439, w_eco127440, w_eco127441, w_eco127442, w_eco127443, w_eco127444, w_eco127445, w_eco127446, w_eco127447, w_eco127448, w_eco127449, w_eco127450, w_eco127451, w_eco127452, w_eco127453, w_eco127454, w_eco127455, w_eco127456, w_eco127457, w_eco127458, w_eco127459, w_eco127460, w_eco127461, w_eco127462, w_eco127463, w_eco127464, w_eco127465, w_eco127466, w_eco127467, w_eco127468, w_eco127469, w_eco127470, w_eco127471, w_eco127472, w_eco127473, w_eco127474, w_eco127475, w_eco127476, w_eco127477, w_eco127478, w_eco127479, w_eco127480, w_eco127481, w_eco127482, w_eco127483, w_eco127484, w_eco127485, w_eco127486, w_eco127487, w_eco127488, w_eco127489, w_eco127490, w_eco127491, w_eco127492, w_eco127493, w_eco127494, w_eco127495, w_eco127496, w_eco127497, w_eco127498, w_eco127499, w_eco127500, w_eco127501, w_eco127502, w_eco127503, w_eco127504, w_eco127505, w_eco127506, w_eco127507, w_eco127508, w_eco127509, w_eco127510, w_eco127511, w_eco127512, w_eco127513, w_eco127514, w_eco127515, w_eco127516, w_eco127517, w_eco127518, w_eco127519, w_eco127520, w_eco127521, w_eco127522, w_eco127523, w_eco127524, w_eco127525, w_eco127526, w_eco127527, w_eco127528, w_eco127529, w_eco127530, w_eco127531, w_eco127532, w_eco127533, w_eco127534, w_eco127535, w_eco127536, w_eco127537, w_eco127538, w_eco127539, w_eco127540, w_eco127541, w_eco127542, w_eco127543, w_eco127544, w_eco127545, w_eco127546, w_eco127547, w_eco127548, w_eco127549, w_eco127550, w_eco127551, w_eco127552, w_eco127553, w_eco127554, w_eco127555, w_eco127556, w_eco127557, w_eco127558, w_eco127559, w_eco127560, w_eco127561, w_eco127562, w_eco127563, w_eco127564, w_eco127565, w_eco127566, w_eco127567, w_eco127568, w_eco127569, w_eco127570, w_eco127571, w_eco127572, w_eco127573, w_eco127574, w_eco127575, w_eco127576, w_eco127577, w_eco127578, w_eco127579, w_eco127580, w_eco127581, w_eco127582, w_eco127583, w_eco127584, w_eco127585, w_eco127586, w_eco127587, w_eco127588, w_eco127589, w_eco127590, w_eco127591, w_eco127592, w_eco127593, w_eco127594, w_eco127595, w_eco127596, w_eco127597, w_eco127598, w_eco127599, w_eco127600, w_eco127601, w_eco127602, w_eco127603, w_eco127604, w_eco127605, w_eco127606, w_eco127607, w_eco127608, w_eco127609, w_eco127610, w_eco127611, w_eco127612, w_eco127613, w_eco127614, w_eco127615, w_eco127616, w_eco127617, w_eco127618, w_eco127619, w_eco127620, w_eco127621, w_eco127622, w_eco127623, w_eco127624, w_eco127625, w_eco127626, w_eco127627, w_eco127628, w_eco127629, w_eco127630, w_eco127631, w_eco127632, w_eco127633, w_eco127634, w_eco127635, w_eco127636, w_eco127637, w_eco127638, w_eco127639, w_eco127640, w_eco127641, w_eco127642, w_eco127643, w_eco127644, w_eco127645, w_eco127646, w_eco127647, w_eco127648, w_eco127649, w_eco127650, w_eco127651, w_eco127652, w_eco127653, w_eco127654, w_eco127655, w_eco127656, w_eco127657, w_eco127658, w_eco127659, w_eco127660, w_eco127661, w_eco127662, w_eco127663, w_eco127664, w_eco127665, w_eco127666, w_eco127667, w_eco127668, w_eco127669, w_eco127670, w_eco127671, w_eco127672, w_eco127673, w_eco127674, w_eco127675, w_eco127676, w_eco127677, w_eco127678, w_eco127679, w_eco127680, w_eco127681, w_eco127682, w_eco127683, w_eco127684, w_eco127685, w_eco127686, w_eco127687, w_eco127688, w_eco127689, w_eco127690, w_eco127691, w_eco127692, w_eco127693, w_eco127694, w_eco127695, w_eco127696, w_eco127697, w_eco127698, w_eco127699, w_eco127700, w_eco127701, w_eco127702, w_eco127703, w_eco127704, w_eco127705, w_eco127706, w_eco127707, w_eco127708, w_eco127709, w_eco127710, w_eco127711, w_eco127712, w_eco127713, w_eco127714, w_eco127715, w_eco127716, w_eco127717, w_eco127718, w_eco127719, w_eco127720, w_eco127721, w_eco127722, w_eco127723, w_eco127724, w_eco127725, w_eco127726, w_eco127727, w_eco127728, w_eco127729, w_eco127730, w_eco127731, w_eco127732, w_eco127733, w_eco127734, w_eco127735, w_eco127736, w_eco127737, w_eco127738, w_eco127739, w_eco127740, w_eco127741, w_eco127742, w_eco127743, w_eco127744, w_eco127745, w_eco127746, w_eco127747, w_eco127748, w_eco127749, w_eco127750, w_eco127751, w_eco127752, w_eco127753, w_eco127754, w_eco127755, w_eco127756, w_eco127757, w_eco127758, w_eco127759, w_eco127760, w_eco127761, w_eco127762, w_eco127763, w_eco127764, w_eco127765, w_eco127766, w_eco127767, w_eco127768, w_eco127769, w_eco127770, w_eco127771, w_eco127772, w_eco127773, w_eco127774, w_eco127775, w_eco127776, w_eco127777, w_eco127778, w_eco127779, w_eco127780, w_eco127781, w_eco127782, w_eco127783, w_eco127784, w_eco127785, w_eco127786, w_eco127787, w_eco127788, w_eco127789, w_eco127790, w_eco127791, w_eco127792, w_eco127793, w_eco127794, w_eco127795, w_eco127796, w_eco127797, w_eco127798, w_eco127799, w_eco127800, w_eco127801, w_eco127802, w_eco127803, w_eco127804, w_eco127805, w_eco127806, w_eco127807, w_eco127808, w_eco127809, w_eco127810, w_eco127811, w_eco127812, w_eco127813, w_eco127814, w_eco127815, w_eco127816, w_eco127817, w_eco127818, w_eco127819, w_eco127820, w_eco127821, w_eco127822, w_eco127823, w_eco127824, w_eco127825, w_eco127826, w_eco127827, w_eco127828, w_eco127829, w_eco127830, w_eco127831, w_eco127832, w_eco127833, w_eco127834, w_eco127835, w_eco127836, w_eco127837, w_eco127838, w_eco127839, w_eco127840, w_eco127841, w_eco127842, w_eco127843, w_eco127844, w_eco127845, w_eco127846, w_eco127847, w_eco127848, w_eco127849, w_eco127850, w_eco127851, w_eco127852, w_eco127853, w_eco127854, w_eco127855, w_eco127856, w_eco127857, w_eco127858, w_eco127859, w_eco127860, w_eco127861, w_eco127862, w_eco127863, w_eco127864, w_eco127865, w_eco127866, w_eco127867, w_eco127868, w_eco127869, w_eco127870, w_eco127871, w_eco127872, w_eco127873, w_eco127874, w_eco127875, w_eco127876, w_eco127877, w_eco127878, w_eco127879, w_eco127880, w_eco127881, w_eco127882, w_eco127883, w_eco127884, w_eco127885, w_eco127886, w_eco127887, w_eco127888, w_eco127889, w_eco127890, w_eco127891, w_eco127892, w_eco127893, w_eco127894, w_eco127895, w_eco127896, w_eco127897, w_eco127898, w_eco127899, w_eco127900, w_eco127901, w_eco127902, w_eco127903, w_eco127904, w_eco127905, w_eco127906, w_eco127907, w_eco127908, w_eco127909, w_eco127910, w_eco127911, w_eco127912, w_eco127913, w_eco127914, w_eco127915, w_eco127916, w_eco127917, w_eco127918, w_eco127919, w_eco127920, w_eco127921, w_eco127922, w_eco127923, w_eco127924, w_eco127925, w_eco127926, w_eco127927, w_eco127928, w_eco127929, w_eco127930, w_eco127931, w_eco127932, w_eco127933, w_eco127934, w_eco127935, w_eco127936, w_eco127937, w_eco127938, w_eco127939, w_eco127940, w_eco127941, w_eco127942, w_eco127943, w_eco127944, w_eco127945, w_eco127946, w_eco127947, w_eco127948, w_eco127949, w_eco127950, w_eco127951, w_eco127952, w_eco127953, w_eco127954, w_eco127955, w_eco127956, w_eco127957, w_eco127958, w_eco127959, w_eco127960, w_eco127961, w_eco127962, w_eco127963, w_eco127964, w_eco127965, w_eco127966, w_eco127967, w_eco127968, w_eco127969, w_eco127970, w_eco127971, w_eco127972, w_eco127973, w_eco127974, w_eco127975, w_eco127976, w_eco127977, w_eco127978, w_eco127979, w_eco127980, w_eco127981, w_eco127982, w_eco127983, w_eco127984, w_eco127985, w_eco127986, w_eco127987, w_eco127988, w_eco127989, w_eco127990, w_eco127991, w_eco127992, w_eco127993, w_eco127994, w_eco127995, w_eco127996, w_eco127997, w_eco127998, w_eco127999, w_eco128000, w_eco128001, w_eco128002, w_eco128003, w_eco128004, w_eco128005, w_eco128006, w_eco128007, w_eco128008, w_eco128009, w_eco128010, w_eco128011, w_eco128012, w_eco128013, w_eco128014, w_eco128015, w_eco128016, w_eco128017, w_eco128018, w_eco128019, w_eco128020, w_eco128021, w_eco128022, w_eco128023, w_eco128024, w_eco128025, w_eco128026, w_eco128027, w_eco128028, w_eco128029, w_eco128030, w_eco128031, w_eco128032, w_eco128033, w_eco128034, w_eco128035, w_eco128036, w_eco128037, w_eco128038, w_eco128039, w_eco128040, w_eco128041, w_eco128042, w_eco128043, w_eco128044, w_eco128045, w_eco128046, w_eco128047, w_eco128048, w_eco128049, w_eco128050, w_eco128051, w_eco128052, w_eco128053, w_eco128054, w_eco128055, w_eco128056, w_eco128057, w_eco128058, w_eco128059, w_eco128060, w_eco128061, w_eco128062, w_eco128063, w_eco128064, w_eco128065, w_eco128066, w_eco128067, w_eco128068, w_eco128069, w_eco128070, w_eco128071, w_eco128072, w_eco128073, w_eco128074, w_eco128075, w_eco128076, w_eco128077, w_eco128078, w_eco128079, w_eco128080, w_eco128081, w_eco128082, w_eco128083, w_eco128084, w_eco128085, w_eco128086, w_eco128087, w_eco128088, w_eco128089, w_eco128090, w_eco128091, w_eco128092, w_eco128093, w_eco128094, w_eco128095, w_eco128096, w_eco128097, w_eco128098, w_eco128099, w_eco128100, w_eco128101, w_eco128102, w_eco128103, w_eco128104, w_eco128105, w_eco128106, w_eco128107, w_eco128108, w_eco128109, w_eco128110, w_eco128111, w_eco128112, w_eco128113, w_eco128114, w_eco128115, w_eco128116, w_eco128117, w_eco128118, w_eco128119, w_eco128120, w_eco128121, w_eco128122, w_eco128123, w_eco128124, w_eco128125, w_eco128126, w_eco128127, w_eco128128, w_eco128129, w_eco128130, w_eco128131, w_eco128132, w_eco128133, w_eco128134, w_eco128135, w_eco128136, w_eco128137, w_eco128138, w_eco128139, w_eco128140, w_eco128141, w_eco128142, w_eco128143, w_eco128144, w_eco128145, w_eco128146, w_eco128147, w_eco128148, w_eco128149, w_eco128150, w_eco128151, w_eco128152, w_eco128153, w_eco128154, w_eco128155, w_eco128156, w_eco128157, w_eco128158, w_eco128159, w_eco128160, w_eco128161, w_eco128162, w_eco128163, w_eco128164, w_eco128165, w_eco128166, w_eco128167, w_eco128168, w_eco128169, w_eco128170, w_eco128171, w_eco128172, w_eco128173, w_eco128174, w_eco128175, w_eco128176, w_eco128177, w_eco128178, w_eco128179, w_eco128180, w_eco128181, w_eco128182, w_eco128183, w_eco128184, w_eco128185, w_eco128186, w_eco128187, w_eco128188, w_eco128189, w_eco128190, w_eco128191, w_eco128192, w_eco128193, w_eco128194, w_eco128195, w_eco128196, w_eco128197, w_eco128198, w_eco128199, w_eco128200, w_eco128201, w_eco128202, w_eco128203, w_eco128204, w_eco128205, w_eco128206, w_eco128207, w_eco128208, w_eco128209, w_eco128210, w_eco128211, w_eco128212, w_eco128213, w_eco128214, w_eco128215, w_eco128216, w_eco128217, w_eco128218, w_eco128219, w_eco128220, w_eco128221, w_eco128222, w_eco128223, w_eco128224, w_eco128225, w_eco128226, w_eco128227, w_eco128228, w_eco128229, w_eco128230, w_eco128231, w_eco128232, w_eco128233, w_eco128234, w_eco128235, w_eco128236, w_eco128237, w_eco128238, w_eco128239, w_eco128240, w_eco128241, w_eco128242, w_eco128243, w_eco128244, w_eco128245, w_eco128246, w_eco128247, w_eco128248, w_eco128249, w_eco128250, w_eco128251, w_eco128252, w_eco128253, w_eco128254, w_eco128255, w_eco128256, w_eco128257, w_eco128258, w_eco128259, w_eco128260, w_eco128261, w_eco128262, w_eco128263, w_eco128264, w_eco128265, w_eco128266, w_eco128267, w_eco128268, w_eco128269, w_eco128270, w_eco128271, w_eco128272, w_eco128273, w_eco128274, w_eco128275, w_eco128276, w_eco128277, w_eco128278, w_eco128279, w_eco128280, w_eco128281, w_eco128282, w_eco128283, w_eco128284, w_eco128285, w_eco128286, w_eco128287, w_eco128288, w_eco128289, w_eco128290, w_eco128291, w_eco128292, w_eco128293, w_eco128294, w_eco128295, w_eco128296, w_eco128297, w_eco128298, w_eco128299, w_eco128300, w_eco128301, w_eco128302, w_eco128303, w_eco128304, w_eco128305, w_eco128306, w_eco128307, w_eco128308, w_eco128309, w_eco128310, w_eco128311, w_eco128312, w_eco128313, w_eco128314, w_eco128315, w_eco128316, w_eco128317, w_eco128318, w_eco128319, w_eco128320, w_eco128321, w_eco128322, w_eco128323, w_eco128324, w_eco128325, w_eco128326, w_eco128327, w_eco128328, w_eco128329, w_eco128330, w_eco128331, w_eco128332, w_eco128333, w_eco128334, w_eco128335, w_eco128336, w_eco128337, w_eco128338, w_eco128339, w_eco128340, w_eco128341, w_eco128342, w_eco128343, w_eco128344, w_eco128345, w_eco128346, w_eco128347, w_eco128348, w_eco128349, w_eco128350, w_eco128351, w_eco128352, w_eco128353, w_eco128354, w_eco128355, w_eco128356, w_eco128357, w_eco128358, w_eco128359, w_eco128360, w_eco128361, w_eco128362, w_eco128363, w_eco128364, w_eco128365, w_eco128366, w_eco128367, w_eco128368, w_eco128369, w_eco128370, w_eco128371, w_eco128372, w_eco128373, w_eco128374, w_eco128375, w_eco128376, w_eco128377, w_eco128378, w_eco128379, w_eco128380, w_eco128381, w_eco128382, w_eco128383, w_eco128384, w_eco128385, w_eco128386, w_eco128387, w_eco128388, w_eco128389, w_eco128390, w_eco128391, w_eco128392, w_eco128393, w_eco128394, w_eco128395, w_eco128396, w_eco128397, w_eco128398, w_eco128399, w_eco128400, w_eco128401, w_eco128402, w_eco128403, w_eco128404, w_eco128405, w_eco128406, w_eco128407, w_eco128408, w_eco128409, w_eco128410, w_eco128411, w_eco128412, w_eco128413, w_eco128414, w_eco128415, w_eco128416, w_eco128417, w_eco128418, w_eco128419, w_eco128420, w_eco128421, w_eco128422, w_eco128423, w_eco128424, w_eco128425, w_eco128426, w_eco128427, w_eco128428, w_eco128429, w_eco128430, w_eco128431, w_eco128432, w_eco128433, w_eco128434, w_eco128435, w_eco128436, w_eco128437, w_eco128438, w_eco128439, w_eco128440, w_eco128441, w_eco128442, w_eco128443, w_eco128444, w_eco128445, w_eco128446, w_eco128447, w_eco128448, w_eco128449, w_eco128450, w_eco128451, w_eco128452, w_eco128453, w_eco128454, w_eco128455, w_eco128456, w_eco128457, w_eco128458, w_eco128459, w_eco128460, w_eco128461, w_eco128462, w_eco128463, w_eco128464, w_eco128465, w_eco128466, w_eco128467, w_eco128468, w_eco128469, w_eco128470, w_eco128471, w_eco128472, w_eco128473, w_eco128474, w_eco128475, w_eco128476, w_eco128477, w_eco128478, w_eco128479, w_eco128480, w_eco128481, w_eco128482, w_eco128483, w_eco128484, w_eco128485, w_eco128486, w_eco128487, w_eco128488, w_eco128489, w_eco128490, w_eco128491, w_eco128492, w_eco128493, w_eco128494, w_eco128495, w_eco128496, w_eco128497, w_eco128498, w_eco128499, w_eco128500, w_eco128501, w_eco128502, w_eco128503, w_eco128504, w_eco128505, w_eco128506, w_eco128507, w_eco128508, w_eco128509, w_eco128510, w_eco128511, w_eco128512, w_eco128513, w_eco128514, w_eco128515, w_eco128516, w_eco128517, w_eco128518, w_eco128519, w_eco128520, w_eco128521, w_eco128522, w_eco128523, w_eco128524, w_eco128525, w_eco128526, w_eco128527, w_eco128528, w_eco128529, w_eco128530, w_eco128531, w_eco128532, w_eco128533, w_eco128534, w_eco128535, w_eco128536, w_eco128537, w_eco128538, w_eco128539, w_eco128540, w_eco128541, w_eco128542, w_eco128543, w_eco128544, w_eco128545, w_eco128546, w_eco128547, w_eco128548, w_eco128549, w_eco128550, w_eco128551, w_eco128552, w_eco128553, w_eco128554, w_eco128555, w_eco128556, w_eco128557, w_eco128558, w_eco128559, w_eco128560, w_eco128561, w_eco128562, w_eco128563, w_eco128564, w_eco128565, w_eco128566, w_eco128567, w_eco128568, w_eco128569, w_eco128570, w_eco128571, w_eco128572, w_eco128573, w_eco128574, w_eco128575, w_eco128576, w_eco128577, w_eco128578, w_eco128579, w_eco128580, w_eco128581, w_eco128582, w_eco128583, w_eco128584, w_eco128585, w_eco128586, w_eco128587, w_eco128588, w_eco128589, w_eco128590, w_eco128591, w_eco128592, w_eco128593, w_eco128594, w_eco128595, w_eco128596, w_eco128597, w_eco128598, w_eco128599, w_eco128600, w_eco128601, w_eco128602, w_eco128603, w_eco128604, w_eco128605, w_eco128606, w_eco128607, w_eco128608, w_eco128609, w_eco128610, w_eco128611, w_eco128612, w_eco128613, w_eco128614, w_eco128615, w_eco128616, w_eco128617, w_eco128618, w_eco128619, w_eco128620, w_eco128621, w_eco128622, w_eco128623, w_eco128624, w_eco128625, w_eco128626, w_eco128627, w_eco128628, w_eco128629, w_eco128630, w_eco128631, w_eco128632, w_eco128633, w_eco128634, w_eco128635, w_eco128636, w_eco128637, w_eco128638, w_eco128639, w_eco128640, w_eco128641, w_eco128642, w_eco128643, w_eco128644, w_eco128645, w_eco128646, w_eco128647, w_eco128648, w_eco128649, w_eco128650, w_eco128651, w_eco128652, w_eco128653, w_eco128654, w_eco128655, w_eco128656, w_eco128657, w_eco128658, w_eco128659, w_eco128660, w_eco128661, w_eco128662, w_eco128663, w_eco128664, w_eco128665, w_eco128666, w_eco128667, w_eco128668, w_eco128669, w_eco128670, w_eco128671, w_eco128672, w_eco128673, w_eco128674, w_eco128675, w_eco128676, w_eco128677, w_eco128678, w_eco128679, w_eco128680, w_eco128681, w_eco128682, w_eco128683, w_eco128684, w_eco128685, w_eco128686, w_eco128687, w_eco128688, w_eco128689, w_eco128690, w_eco128691, w_eco128692, w_eco128693, w_eco128694, w_eco128695, w_eco128696, w_eco128697, w_eco128698, w_eco128699, w_eco128700, w_eco128701, w_eco128702, w_eco128703, w_eco128704, w_eco128705, w_eco128706, w_eco128707, w_eco128708, w_eco128709, w_eco128710, w_eco128711, w_eco128712, w_eco128713, w_eco128714, w_eco128715, w_eco128716, w_eco128717, w_eco128718, w_eco128719, w_eco128720, w_eco128721, w_eco128722, w_eco128723, w_eco128724, w_eco128725, w_eco128726, w_eco128727, w_eco128728, w_eco128729, w_eco128730, w_eco128731, w_eco128732, w_eco128733, w_eco128734, w_eco128735, w_eco128736, w_eco128737, w_eco128738, w_eco128739, w_eco128740, w_eco128741, w_eco128742, w_eco128743, w_eco128744, w_eco128745, w_eco128746, w_eco128747, w_eco128748, w_eco128749, w_eco128750, w_eco128751, w_eco128752, w_eco128753, w_eco128754, w_eco128755, w_eco128756, w_eco128757, w_eco128758, w_eco128759, w_eco128760, w_eco128761, w_eco128762, w_eco128763, w_eco128764, w_eco128765, w_eco128766, w_eco128767, w_eco128768, w_eco128769, w_eco128770, w_eco128771, w_eco128772, w_eco128773, w_eco128774, w_eco128775, w_eco128776, w_eco128777, w_eco128778, w_eco128779, w_eco128780, w_eco128781, w_eco128782, w_eco128783, w_eco128784, w_eco128785, w_eco128786, w_eco128787, w_eco128788, w_eco128789, w_eco128790, w_eco128791, w_eco128792, w_eco128793, w_eco128794, w_eco128795, w_eco128796, w_eco128797, w_eco128798, w_eco128799, w_eco128800, w_eco128801, w_eco128802, w_eco128803, w_eco128804, w_eco128805, w_eco128806, w_eco128807, w_eco128808, w_eco128809, w_eco128810, w_eco128811, w_eco128812, w_eco128813, w_eco128814, w_eco128815, w_eco128816, w_eco128817, w_eco128818, w_eco128819, w_eco128820, w_eco128821, w_eco128822, w_eco128823, w_eco128824, w_eco128825, w_eco128826, w_eco128827, w_eco128828, w_eco128829, w_eco128830, w_eco128831, w_eco128832, w_eco128833, w_eco128834, w_eco128835, w_eco128836, w_eco128837, w_eco128838, w_eco128839, w_eco128840, w_eco128841, w_eco128842, w_eco128843, w_eco128844, w_eco128845, w_eco128846, w_eco128847, w_eco128848, w_eco128849, w_eco128850, w_eco128851, w_eco128852, w_eco128853, w_eco128854, w_eco128855, w_eco128856, w_eco128857, w_eco128858, w_eco128859, w_eco128860, w_eco128861, w_eco128862, w_eco128863, w_eco128864, w_eco128865, w_eco128866, w_eco128867, w_eco128868, w_eco128869, w_eco128870, w_eco128871, w_eco128872, w_eco128873, w_eco128874, w_eco128875, w_eco128876, w_eco128877, w_eco128878, w_eco128879, w_eco128880, w_eco128881, w_eco128882, w_eco128883, w_eco128884, w_eco128885, w_eco128886, w_eco128887, w_eco128888, w_eco128889, w_eco128890, w_eco128891, w_eco128892, w_eco128893, w_eco128894, w_eco128895, w_eco128896, w_eco128897, w_eco128898, w_eco128899, w_eco128900, w_eco128901, w_eco128902, w_eco128903, w_eco128904, w_eco128905, w_eco128906, w_eco128907, w_eco128908, w_eco128909, w_eco128910, w_eco128911, w_eco128912, w_eco128913, w_eco128914, w_eco128915, w_eco128916, w_eco128917, w_eco128918, w_eco128919, w_eco128920, w_eco128921, w_eco128922, w_eco128923, w_eco128924, w_eco128925, w_eco128926, w_eco128927, w_eco128928, w_eco128929, w_eco128930, w_eco128931, w_eco128932, w_eco128933, w_eco128934, w_eco128935, w_eco128936, w_eco128937, w_eco128938, w_eco128939, w_eco128940, w_eco128941, w_eco128942, w_eco128943, w_eco128944, w_eco128945, w_eco128946, w_eco128947, w_eco128948, w_eco128949, w_eco128950, w_eco128951, w_eco128952, w_eco128953, w_eco128954, w_eco128955, w_eco128956, w_eco128957, w_eco128958, w_eco128959, w_eco128960, w_eco128961, w_eco128962, w_eco128963, w_eco128964, w_eco128965, w_eco128966, w_eco128967, w_eco128968, w_eco128969, w_eco128970, w_eco128971, w_eco128972, w_eco128973, w_eco128974, w_eco128975, w_eco128976, w_eco128977, w_eco128978, w_eco128979, w_eco128980, w_eco128981, w_eco128982, w_eco128983, w_eco128984, w_eco128985, w_eco128986, w_eco128987, w_eco128988, w_eco128989, w_eco128990, w_eco128991, w_eco128992, w_eco128993, w_eco128994, w_eco128995, w_eco128996, w_eco128997, w_eco128998, w_eco128999, w_eco129000, w_eco129001, w_eco129002, w_eco129003, w_eco129004, w_eco129005, w_eco129006, w_eco129007, w_eco129008, w_eco129009, w_eco129010, w_eco129011, w_eco129012, w_eco129013, w_eco129014, w_eco129015, w_eco129016, w_eco129017, w_eco129018, w_eco129019, w_eco129020, w_eco129021, w_eco129022, w_eco129023, w_eco129024, w_eco129025, w_eco129026, w_eco129027, w_eco129028, w_eco129029, w_eco129030, w_eco129031, w_eco129032, w_eco129033, w_eco129034, w_eco129035, w_eco129036, w_eco129037, w_eco129038, w_eco129039, w_eco129040, w_eco129041, w_eco129042, w_eco129043, w_eco129044, w_eco129045, w_eco129046, w_eco129047, w_eco129048, w_eco129049, w_eco129050, w_eco129051, w_eco129052, w_eco129053, w_eco129054, w_eco129055, w_eco129056, w_eco129057, w_eco129058, w_eco129059, w_eco129060, w_eco129061, w_eco129062, w_eco129063, w_eco129064, w_eco129065, w_eco129066, w_eco129067, w_eco129068, w_eco129069, w_eco129070, w_eco129071, w_eco129072, w_eco129073, w_eco129074, w_eco129075, w_eco129076, w_eco129077, w_eco129078, w_eco129079, w_eco129080, w_eco129081, w_eco129082, w_eco129083, w_eco129084, w_eco129085, w_eco129086, w_eco129087, w_eco129088, w_eco129089, w_eco129090, w_eco129091, w_eco129092, w_eco129093, w_eco129094, w_eco129095, w_eco129096, w_eco129097, w_eco129098, w_eco129099, w_eco129100, w_eco129101, w_eco129102, w_eco129103, w_eco129104, w_eco129105, w_eco129106, w_eco129107, w_eco129108, w_eco129109, w_eco129110, w_eco129111, w_eco129112, w_eco129113, w_eco129114, w_eco129115, w_eco129116, w_eco129117, w_eco129118, w_eco129119, w_eco129120, w_eco129121, w_eco129122, w_eco129123, w_eco129124, w_eco129125, w_eco129126, w_eco129127, w_eco129128, w_eco129129, w_eco129130, w_eco129131, w_eco129132, w_eco129133, w_eco129134, w_eco129135, w_eco129136, w_eco129137, w_eco129138, w_eco129139, w_eco129140, w_eco129141, w_eco129142, w_eco129143, w_eco129144, w_eco129145, w_eco129146, w_eco129147, w_eco129148, w_eco129149, w_eco129150, w_eco129151, w_eco129152, w_eco129153, w_eco129154, w_eco129155, w_eco129156, w_eco129157, w_eco129158, w_eco129159, w_eco129160, w_eco129161, w_eco129162, w_eco129163, w_eco129164, w_eco129165, w_eco129166, w_eco129167, w_eco129168, w_eco129169, w_eco129170, w_eco129171, w_eco129172, w_eco129173, w_eco129174, w_eco129175, w_eco129176, w_eco129177, w_eco129178, w_eco129179, w_eco129180, w_eco129181, w_eco129182, w_eco129183, w_eco129184, w_eco129185, w_eco129186, w_eco129187, w_eco129188, w_eco129189, w_eco129190, w_eco129191, w_eco129192, w_eco129193, w_eco129194, w_eco129195, w_eco129196, w_eco129197, w_eco129198, w_eco129199, w_eco129200, w_eco129201, w_eco129202, w_eco129203, w_eco129204, w_eco129205, w_eco129206, w_eco129207, w_eco129208, w_eco129209, w_eco129210, w_eco129211, w_eco129212, w_eco129213, w_eco129214, w_eco129215, w_eco129216, w_eco129217, w_eco129218, w_eco129219, w_eco129220, w_eco129221, w_eco129222, w_eco129223, w_eco129224, w_eco129225, w_eco129226, w_eco129227, w_eco129228, w_eco129229, w_eco129230, w_eco129231, w_eco129232, w_eco129233, w_eco129234, w_eco129235, w_eco129236, w_eco129237, w_eco129238, w_eco129239, w_eco129240, w_eco129241, w_eco129242, w_eco129243, w_eco129244, w_eco129245, w_eco129246, w_eco129247, w_eco129248, w_eco129249, w_eco129250, w_eco129251, w_eco129252, w_eco129253, w_eco129254, w_eco129255, w_eco129256, w_eco129257, w_eco129258, w_eco129259, w_eco129260, w_eco129261, w_eco129262, w_eco129263, w_eco129264, w_eco129265, w_eco129266, w_eco129267, w_eco129268, w_eco129269, w_eco129270, w_eco129271, w_eco129272, w_eco129273, w_eco129274, w_eco129275, w_eco129276, w_eco129277, w_eco129278, w_eco129279, w_eco129280, w_eco129281, w_eco129282, w_eco129283, w_eco129284, w_eco129285, w_eco129286, w_eco129287, w_eco129288, w_eco129289, w_eco129290, w_eco129291, w_eco129292, w_eco129293, w_eco129294, w_eco129295, w_eco129296, w_eco129297, w_eco129298, w_eco129299, w_eco129300, w_eco129301, w_eco129302, w_eco129303, w_eco129304, w_eco129305, w_eco129306, w_eco129307, w_eco129308, w_eco129309, w_eco129310, w_eco129311, w_eco129312, w_eco129313, w_eco129314, w_eco129315, w_eco129316, w_eco129317, w_eco129318, w_eco129319, w_eco129320, w_eco129321, w_eco129322, w_eco129323, w_eco129324, w_eco129325, w_eco129326, w_eco129327, w_eco129328, w_eco129329, w_eco129330, w_eco129331, w_eco129332, w_eco129333, w_eco129334, w_eco129335, w_eco129336, w_eco129337, w_eco129338, w_eco129339, w_eco129340, w_eco129341, w_eco129342, w_eco129343, w_eco129344, w_eco129345, w_eco129346, w_eco129347, w_eco129348, w_eco129349, w_eco129350, w_eco129351, w_eco129352, w_eco129353, w_eco129354, w_eco129355, w_eco129356, w_eco129357, w_eco129358, w_eco129359, w_eco129360, w_eco129361, w_eco129362, w_eco129363, w_eco129364, w_eco129365, w_eco129366, w_eco129367, w_eco129368, w_eco129369, w_eco129370, w_eco129371, w_eco129372, w_eco129373, w_eco129374, w_eco129375, w_eco129376, w_eco129377, w_eco129378, w_eco129379, w_eco129380, w_eco129381, w_eco129382, w_eco129383, w_eco129384, w_eco129385, w_eco129386, w_eco129387, w_eco129388, w_eco129389, w_eco129390, w_eco129391, w_eco129392, w_eco129393, w_eco129394, w_eco129395, w_eco129396, w_eco129397, w_eco129398, w_eco129399, w_eco129400, w_eco129401, w_eco129402, w_eco129403, w_eco129404, w_eco129405, w_eco129406, w_eco129407, w_eco129408, w_eco129409, w_eco129410, w_eco129411, w_eco129412, w_eco129413, w_eco129414, w_eco129415, w_eco129416, w_eco129417, w_eco129418, w_eco129419, w_eco129420, w_eco129421, w_eco129422, w_eco129423, w_eco129424, w_eco129425, w_eco129426, w_eco129427, w_eco129428, w_eco129429, w_eco129430, w_eco129431, w_eco129432, w_eco129433, w_eco129434, w_eco129435, w_eco129436, w_eco129437, w_eco129438, w_eco129439, w_eco129440, w_eco129441, w_eco129442, w_eco129443, w_eco129444, w_eco129445, w_eco129446, w_eco129447, w_eco129448, w_eco129449, w_eco129450, w_eco129451, w_eco129452, w_eco129453, w_eco129454, w_eco129455, w_eco129456, w_eco129457, w_eco129458, w_eco129459, w_eco129460, w_eco129461, w_eco129462, w_eco129463, w_eco129464, w_eco129465, w_eco129466, w_eco129467, w_eco129468, w_eco129469, w_eco129470, w_eco129471, w_eco129472, w_eco129473, w_eco129474, w_eco129475, w_eco129476, w_eco129477, w_eco129478, w_eco129479, w_eco129480, w_eco129481, w_eco129482, w_eco129483, w_eco129484, w_eco129485, w_eco129486, w_eco129487, w_eco129488, w_eco129489, w_eco129490, w_eco129491, w_eco129492, w_eco129493, w_eco129494, w_eco129495, w_eco129496, w_eco129497, w_eco129498, w_eco129499, w_eco129500, w_eco129501, w_eco129502, w_eco129503, w_eco129504, w_eco129505, w_eco129506, w_eco129507, w_eco129508, w_eco129509, w_eco129510, w_eco129511, w_eco129512, w_eco129513, w_eco129514, w_eco129515, w_eco129516, w_eco129517, w_eco129518, w_eco129519, w_eco129520, w_eco129521, w_eco129522, w_eco129523, w_eco129524, w_eco129525, w_eco129526, w_eco129527, w_eco129528, w_eco129529, w_eco129530, w_eco129531, w_eco129532, w_eco129533, w_eco129534, w_eco129535, w_eco129536, w_eco129537, w_eco129538, w_eco129539, w_eco129540, w_eco129541, w_eco129542, w_eco129543, w_eco129544, w_eco129545, w_eco129546, w_eco129547, w_eco129548, w_eco129549, w_eco129550, w_eco129551, w_eco129552, w_eco129553, w_eco129554, w_eco129555, w_eco129556, w_eco129557, w_eco129558, w_eco129559, w_eco129560, w_eco129561, w_eco129562, w_eco129563, w_eco129564, w_eco129565, w_eco129566, w_eco129567, w_eco129568, w_eco129569, w_eco129570, w_eco129571, w_eco129572, w_eco129573, w_eco129574, w_eco129575, w_eco129576, w_eco129577, w_eco129578, w_eco129579, w_eco129580, w_eco129581, w_eco129582, w_eco129583, w_eco129584, w_eco129585, w_eco129586, w_eco129587, w_eco129588, w_eco129589, w_eco129590, w_eco129591, w_eco129592, w_eco129593, w_eco129594, w_eco129595, w_eco129596, w_eco129597, w_eco129598, w_eco129599, w_eco129600, w_eco129601, w_eco129602, w_eco129603, w_eco129604, w_eco129605, w_eco129606, w_eco129607, w_eco129608, w_eco129609, w_eco129610, w_eco129611, w_eco129612, w_eco129613, w_eco129614, w_eco129615, w_eco129616, w_eco129617, w_eco129618, w_eco129619, w_eco129620, w_eco129621, w_eco129622, w_eco129623, w_eco129624, w_eco129625, w_eco129626, w_eco129627, w_eco129628, w_eco129629, w_eco129630, w_eco129631, w_eco129632, w_eco129633, w_eco129634, w_eco129635, w_eco129636, w_eco129637, w_eco129638, w_eco129639, w_eco129640, w_eco129641, w_eco129642, w_eco129643, w_eco129644, w_eco129645, w_eco129646, w_eco129647, w_eco129648, w_eco129649, w_eco129650, w_eco129651, w_eco129652, w_eco129653, w_eco129654, w_eco129655, w_eco129656, w_eco129657, w_eco129658, w_eco129659, w_eco129660, w_eco129661, w_eco129662, w_eco129663, w_eco129664, w_eco129665, w_eco129666, w_eco129667, w_eco129668, w_eco129669, w_eco129670, w_eco129671, w_eco129672, w_eco129673, w_eco129674, w_eco129675, w_eco129676, w_eco129677, w_eco129678, w_eco129679, w_eco129680, w_eco129681, w_eco129682, w_eco129683, w_eco129684, w_eco129685, w_eco129686, w_eco129687, w_eco129688, w_eco129689, w_eco129690, w_eco129691, w_eco129692, w_eco129693, w_eco129694, w_eco129695, w_eco129696, w_eco129697, w_eco129698, w_eco129699, w_eco129700, w_eco129701, w_eco129702, w_eco129703, w_eco129704, w_eco129705, w_eco129706, w_eco129707, w_eco129708, w_eco129709, w_eco129710, w_eco129711, w_eco129712, w_eco129713, w_eco129714, w_eco129715, w_eco129716, w_eco129717, w_eco129718, w_eco129719, w_eco129720, w_eco129721, w_eco129722, w_eco129723, w_eco129724, w_eco129725, w_eco129726, w_eco129727, w_eco129728, w_eco129729, w_eco129730, w_eco129731, w_eco129732, w_eco129733, w_eco129734, w_eco129735, w_eco129736, w_eco129737, w_eco129738, w_eco129739, w_eco129740, w_eco129741, w_eco129742, w_eco129743, w_eco129744, w_eco129745, w_eco129746, w_eco129747, w_eco129748, w_eco129749, w_eco129750, w_eco129751, w_eco129752, w_eco129753, w_eco129754, w_eco129755, w_eco129756, w_eco129757, w_eco129758, w_eco129759, w_eco129760, w_eco129761, w_eco129762, w_eco129763, w_eco129764, w_eco129765, w_eco129766, w_eco129767, w_eco129768, w_eco129769, w_eco129770, w_eco129771, w_eco129772, w_eco129773, w_eco129774, w_eco129775, w_eco129776, w_eco129777, w_eco129778, w_eco129779, w_eco129780, w_eco129781, w_eco129782, w_eco129783, w_eco129784, w_eco129785, w_eco129786, w_eco129787, w_eco129788, w_eco129789, w_eco129790, w_eco129791, w_eco129792, w_eco129793, w_eco129794, w_eco129795, w_eco129796, w_eco129797, w_eco129798, w_eco129799, w_eco129800, w_eco129801, w_eco129802, w_eco129803, w_eco129804, w_eco129805, w_eco129806, w_eco129807, w_eco129808, w_eco129809, w_eco129810, w_eco129811, w_eco129812, w_eco129813, w_eco129814, w_eco129815, w_eco129816, w_eco129817, w_eco129818, w_eco129819, w_eco129820, w_eco129821, w_eco129822, w_eco129823, w_eco129824, w_eco129825, w_eco129826, w_eco129827, w_eco129828, w_eco129829, w_eco129830, w_eco129831, w_eco129832, w_eco129833, w_eco129834, w_eco129835, w_eco129836, w_eco129837, w_eco129838, w_eco129839, w_eco129840, w_eco129841, w_eco129842, w_eco129843, w_eco129844, w_eco129845, w_eco129846, w_eco129847, w_eco129848, w_eco129849, w_eco129850, w_eco129851, w_eco129852, w_eco129853, w_eco129854, w_eco129855, w_eco129856, w_eco129857, w_eco129858, w_eco129859, w_eco129860, w_eco129861, w_eco129862, w_eco129863, w_eco129864, w_eco129865, w_eco129866, w_eco129867, w_eco129868, w_eco129869, w_eco129870, w_eco129871, w_eco129872, w_eco129873, w_eco129874, w_eco129875, w_eco129876, w_eco129877, w_eco129878, w_eco129879, w_eco129880, w_eco129881, w_eco129882, w_eco129883, w_eco129884, w_eco129885, w_eco129886, w_eco129887, w_eco129888, w_eco129889, w_eco129890, w_eco129891, w_eco129892, w_eco129893, w_eco129894, w_eco129895, w_eco129896, w_eco129897, w_eco129898, w_eco129899, w_eco129900, w_eco129901, w_eco129902, w_eco129903, w_eco129904, w_eco129905, w_eco129906, w_eco129907, w_eco129908, w_eco129909, w_eco129910, w_eco129911, w_eco129912, w_eco129913, w_eco129914, w_eco129915, w_eco129916, w_eco129917, w_eco129918, w_eco129919, w_eco129920, w_eco129921, w_eco129922, w_eco129923, w_eco129924, w_eco129925, w_eco129926, w_eco129927, w_eco129928, w_eco129929, w_eco129930, w_eco129931, w_eco129932, w_eco129933, w_eco129934, w_eco129935, w_eco129936, w_eco129937, w_eco129938, w_eco129939, w_eco129940, w_eco129941, w_eco129942, w_eco129943, w_eco129944, w_eco129945, w_eco129946, w_eco129947, w_eco129948, w_eco129949, w_eco129950, w_eco129951, w_eco129952, w_eco129953, w_eco129954, w_eco129955, w_eco129956, w_eco129957, w_eco129958, w_eco129959, w_eco129960, w_eco129961, w_eco129962, w_eco129963, w_eco129964, w_eco129965, w_eco129966, w_eco129967, w_eco129968, w_eco129969, w_eco129970, w_eco129971, w_eco129972, w_eco129973, w_eco129974, w_eco129975, w_eco129976, w_eco129977, w_eco129978, w_eco129979, w_eco129980, w_eco129981, w_eco129982, w_eco129983, w_eco129984, w_eco129985, w_eco129986, w_eco129987, w_eco129988, w_eco129989, w_eco129990, w_eco129991, w_eco129992, w_eco129993, w_eco129994, w_eco129995, w_eco129996, w_eco129997, w_eco129998, w_eco129999, w_eco130000, w_eco130001, w_eco130002, w_eco130003, w_eco130004, w_eco130005, w_eco130006, w_eco130007, w_eco130008, w_eco130009, w_eco130010, w_eco130011, w_eco130012, w_eco130013, w_eco130014, w_eco130015, w_eco130016, w_eco130017, w_eco130018, w_eco130019, w_eco130020, w_eco130021, w_eco130022, w_eco130023, w_eco130024, w_eco130025, w_eco130026, w_eco130027, w_eco130028, w_eco130029, w_eco130030, w_eco130031, w_eco130032, w_eco130033, w_eco130034, w_eco130035, w_eco130036, w_eco130037, w_eco130038, w_eco130039, w_eco130040, w_eco130041, w_eco130042, w_eco130043, w_eco130044, w_eco130045, w_eco130046, w_eco130047, w_eco130048, w_eco130049, w_eco130050, w_eco130051, w_eco130052, w_eco130053, w_eco130054, w_eco130055, w_eco130056, w_eco130057, w_eco130058, w_eco130059, w_eco130060, w_eco130061, w_eco130062, w_eco130063, w_eco130064, w_eco130065, w_eco130066, w_eco130067, w_eco130068, w_eco130069, w_eco130070, w_eco130071, w_eco130072, w_eco130073, w_eco130074, w_eco130075, w_eco130076, w_eco130077, w_eco130078, w_eco130079, w_eco130080, w_eco130081, w_eco130082, w_eco130083, w_eco130084, w_eco130085, w_eco130086, w_eco130087, w_eco130088, w_eco130089, w_eco130090, w_eco130091, w_eco130092, w_eco130093, w_eco130094, w_eco130095, w_eco130096, w_eco130097, w_eco130098, w_eco130099, w_eco130100, w_eco130101, w_eco130102, w_eco130103, w_eco130104, w_eco130105, w_eco130106, w_eco130107, w_eco130108, w_eco130109, w_eco130110, w_eco130111, w_eco130112, w_eco130113, w_eco130114, w_eco130115, w_eco130116, w_eco130117, w_eco130118, w_eco130119, w_eco130120, w_eco130121, w_eco130122, w_eco130123, w_eco130124, w_eco130125, w_eco130126, w_eco130127, w_eco130128, w_eco130129, w_eco130130, w_eco130131, w_eco130132, w_eco130133, w_eco130134, w_eco130135, w_eco130136, w_eco130137, w_eco130138, w_eco130139, w_eco130140, w_eco130141, w_eco130142, w_eco130143, w_eco130144, w_eco130145, w_eco130146, w_eco130147, w_eco130148, w_eco130149, w_eco130150, w_eco130151, w_eco130152, w_eco130153, w_eco130154, w_eco130155, w_eco130156, w_eco130157, w_eco130158, w_eco130159, w_eco130160, w_eco130161, w_eco130162, w_eco130163, w_eco130164, w_eco130165, w_eco130166, w_eco130167, w_eco130168, w_eco130169, w_eco130170, w_eco130171, w_eco130172, w_eco130173, w_eco130174, w_eco130175, w_eco130176, w_eco130177, w_eco130178, w_eco130179, w_eco130180, w_eco130181, w_eco130182, w_eco130183, w_eco130184, w_eco130185, w_eco130186, w_eco130187, w_eco130188, w_eco130189, w_eco130190, w_eco130191, w_eco130192, w_eco130193, w_eco130194, w_eco130195, w_eco130196, w_eco130197, w_eco130198, w_eco130199, w_eco130200, w_eco130201, w_eco130202, w_eco130203, w_eco130204, w_eco130205, w_eco130206, w_eco130207, w_eco130208, w_eco130209, w_eco130210, w_eco130211, w_eco130212, w_eco130213, w_eco130214, w_eco130215, w_eco130216, w_eco130217, w_eco130218, w_eco130219, w_eco130220, w_eco130221, w_eco130222, w_eco130223, w_eco130224, w_eco130225, w_eco130226, w_eco130227, w_eco130228, w_eco130229, w_eco130230, w_eco130231, w_eco130232, w_eco130233, w_eco130234, w_eco130235, w_eco130236, w_eco130237, w_eco130238, w_eco130239, w_eco130240, w_eco130241, w_eco130242, w_eco130243, w_eco130244, w_eco130245, w_eco130246, w_eco130247, w_eco130248, w_eco130249, w_eco130250, w_eco130251, w_eco130252, w_eco130253, w_eco130254, w_eco130255, w_eco130256, w_eco130257, w_eco130258, w_eco130259, w_eco130260, w_eco130261, w_eco130262, w_eco130263, w_eco130264, w_eco130265, w_eco130266, w_eco130267, w_eco130268, w_eco130269, w_eco130270, w_eco130271, w_eco130272, w_eco130273, w_eco130274, w_eco130275, w_eco130276, w_eco130277, w_eco130278, w_eco130279, w_eco130280, w_eco130281, w_eco130282, w_eco130283, w_eco130284, w_eco130285, w_eco130286, w_eco130287, w_eco130288, w_eco130289, w_eco130290, w_eco130291, w_eco130292, w_eco130293, w_eco130294, w_eco130295, w_eco130296, w_eco130297, w_eco130298, w_eco130299, w_eco130300, w_eco130301, w_eco130302, w_eco130303, w_eco130304, w_eco130305, w_eco130306, w_eco130307, w_eco130308, w_eco130309, w_eco130310, w_eco130311, w_eco130312, w_eco130313, w_eco130314, w_eco130315, w_eco130316, w_eco130317, w_eco130318, w_eco130319, w_eco130320, w_eco130321, w_eco130322, w_eco130323, w_eco130324, w_eco130325, w_eco130326, w_eco130327, w_eco130328, w_eco130329, w_eco130330, w_eco130331, w_eco130332, w_eco130333, w_eco130334, w_eco130335, w_eco130336, w_eco130337, w_eco130338, w_eco130339, w_eco130340, w_eco130341, w_eco130342, w_eco130343, w_eco130344, w_eco130345, w_eco130346, w_eco130347, w_eco130348, w_eco130349, w_eco130350, w_eco130351, w_eco130352, w_eco130353, w_eco130354, w_eco130355, w_eco130356, w_eco130357, w_eco130358, w_eco130359, w_eco130360, w_eco130361, w_eco130362, w_eco130363, w_eco130364, w_eco130365, w_eco130366, w_eco130367, w_eco130368, w_eco130369, w_eco130370, w_eco130371, w_eco130372, w_eco130373, w_eco130374, w_eco130375, w_eco130376, w_eco130377, w_eco130378, w_eco130379, w_eco130380, w_eco130381, w_eco130382, w_eco130383, w_eco130384, w_eco130385, w_eco130386, w_eco130387, w_eco130388, w_eco130389, w_eco130390, w_eco130391, w_eco130392, w_eco130393, w_eco130394, w_eco130395, w_eco130396, w_eco130397, w_eco130398, w_eco130399, w_eco130400, w_eco130401, w_eco130402, w_eco130403, w_eco130404, w_eco130405, w_eco130406, w_eco130407, w_eco130408, w_eco130409, w_eco130410, w_eco130411, w_eco130412, w_eco130413, w_eco130414, w_eco130415, w_eco130416, w_eco130417, w_eco130418, w_eco130419, w_eco130420, w_eco130421, w_eco130422, w_eco130423, w_eco130424, w_eco130425, w_eco130426, w_eco130427, w_eco130428, w_eco130429, w_eco130430, w_eco130431, w_eco130432, w_eco130433, w_eco130434, w_eco130435, w_eco130436, w_eco130437, w_eco130438, w_eco130439, w_eco130440, w_eco130441, w_eco130442, w_eco130443, w_eco130444, w_eco130445, w_eco130446, w_eco130447, w_eco130448, w_eco130449, w_eco130450, w_eco130451, w_eco130452, w_eco130453, w_eco130454, w_eco130455, w_eco130456, w_eco130457, w_eco130458, w_eco130459, w_eco130460, w_eco130461, w_eco130462, w_eco130463, w_eco130464, w_eco130465, w_eco130466, w_eco130467, w_eco130468, w_eco130469, w_eco130470, w_eco130471, w_eco130472, w_eco130473, w_eco130474, w_eco130475, w_eco130476, w_eco130477, w_eco130478, w_eco130479, w_eco130480, w_eco130481, w_eco130482, w_eco130483, w_eco130484, w_eco130485, w_eco130486, w_eco130487, w_eco130488, w_eco130489, w_eco130490, w_eco130491, w_eco130492, w_eco130493, w_eco130494, w_eco130495, w_eco130496, w_eco130497, w_eco130498, w_eco130499, w_eco130500, w_eco130501, w_eco130502, w_eco130503, w_eco130504, w_eco130505, w_eco130506, w_eco130507, w_eco130508, w_eco130509, w_eco130510, w_eco130511, w_eco130512, w_eco130513, w_eco130514, w_eco130515, w_eco130516, w_eco130517, w_eco130518, w_eco130519, w_eco130520, w_eco130521, w_eco130522, w_eco130523, w_eco130524, w_eco130525, w_eco130526, w_eco130527, w_eco130528, w_eco130529, w_eco130530, w_eco130531, w_eco130532, w_eco130533, w_eco130534, w_eco130535, w_eco130536, w_eco130537, w_eco130538, w_eco130539, w_eco130540, w_eco130541, w_eco130542, w_eco130543, w_eco130544, w_eco130545, w_eco130546, w_eco130547, w_eco130548, w_eco130549, w_eco130550, w_eco130551, w_eco130552, w_eco130553, w_eco130554, w_eco130555, w_eco130556, w_eco130557, w_eco130558, w_eco130559, w_eco130560, w_eco130561, w_eco130562, w_eco130563, w_eco130564, w_eco130565, w_eco130566, w_eco130567, w_eco130568, w_eco130569, w_eco130570, w_eco130571, w_eco130572, w_eco130573, w_eco130574, w_eco130575, w_eco130576, w_eco130577, w_eco130578, w_eco130579, w_eco130580, w_eco130581, w_eco130582, w_eco130583, w_eco130584, w_eco130585, w_eco130586, w_eco130587, w_eco130588, w_eco130589, w_eco130590, w_eco130591, w_eco130592, w_eco130593, w_eco130594, w_eco130595, w_eco130596, w_eco130597, w_eco130598, w_eco130599, w_eco130600, w_eco130601, w_eco130602, w_eco130603, w_eco130604, w_eco130605, w_eco130606, w_eco130607, w_eco130608, w_eco130609, w_eco130610, w_eco130611, w_eco130612, w_eco130613, w_eco130614, w_eco130615, w_eco130616, w_eco130617, w_eco130618, w_eco130619, w_eco130620, w_eco130621, w_eco130622, w_eco130623, w_eco130624, w_eco130625, w_eco130626, w_eco130627, w_eco130628, w_eco130629, w_eco130630, w_eco130631, w_eco130632, w_eco130633, w_eco130634, w_eco130635, w_eco130636, w_eco130637, w_eco130638, w_eco130639, w_eco130640, w_eco130641, w_eco130642, w_eco130643, w_eco130644, w_eco130645, w_eco130646, w_eco130647, w_eco130648, w_eco130649, w_eco130650, w_eco130651, w_eco130652, w_eco130653, w_eco130654, w_eco130655, w_eco130656, w_eco130657, w_eco130658, w_eco130659, w_eco130660, w_eco130661, w_eco130662, w_eco130663, w_eco130664, w_eco130665, w_eco130666, w_eco130667, w_eco130668, w_eco130669, w_eco130670, w_eco130671, w_eco130672, w_eco130673, w_eco130674, w_eco130675, w_eco130676, w_eco130677, w_eco130678, w_eco130679, w_eco130680, w_eco130681, w_eco130682, w_eco130683, w_eco130684, w_eco130685, w_eco130686, w_eco130687, w_eco130688, w_eco130689, w_eco130690, w_eco130691, w_eco130692, w_eco130693, w_eco130694, w_eco130695, w_eco130696, w_eco130697, w_eco130698, w_eco130699, w_eco130700, w_eco130701, w_eco130702, w_eco130703, w_eco130704, w_eco130705, w_eco130706, w_eco130707, w_eco130708, w_eco130709, w_eco130710, w_eco130711, w_eco130712, w_eco130713, w_eco130714, w_eco130715, w_eco130716, w_eco130717, w_eco130718, w_eco130719, w_eco130720, w_eco130721, w_eco130722, w_eco130723, w_eco130724, w_eco130725, w_eco130726, w_eco130727, w_eco130728, w_eco130729, w_eco130730, w_eco130731, w_eco130732, w_eco130733, w_eco130734, w_eco130735, w_eco130736, w_eco130737, w_eco130738, w_eco130739, w_eco130740, w_eco130741, w_eco130742, w_eco130743, w_eco130744, w_eco130745, w_eco130746, w_eco130747, w_eco130748, w_eco130749, w_eco130750, w_eco130751, w_eco130752, w_eco130753, w_eco130754, w_eco130755, w_eco130756, w_eco130757, w_eco130758, w_eco130759, w_eco130760, w_eco130761, w_eco130762, w_eco130763, w_eco130764, w_eco130765, w_eco130766, w_eco130767, w_eco130768, w_eco130769, w_eco130770, w_eco130771, w_eco130772, w_eco130773, w_eco130774, w_eco130775, w_eco130776, w_eco130777, w_eco130778, w_eco130779, w_eco130780, w_eco130781, w_eco130782, w_eco130783, w_eco130784, w_eco130785, w_eco130786, w_eco130787, w_eco130788, w_eco130789, w_eco130790, w_eco130791, w_eco130792, w_eco130793, w_eco130794, w_eco130795, w_eco130796, w_eco130797, w_eco130798, w_eco130799, w_eco130800, w_eco130801, w_eco130802, w_eco130803, w_eco130804, w_eco130805, w_eco130806, w_eco130807, w_eco130808, w_eco130809, w_eco130810, w_eco130811, w_eco130812, w_eco130813, w_eco130814, w_eco130815, w_eco130816, w_eco130817, w_eco130818, w_eco130819, w_eco130820, w_eco130821, w_eco130822, w_eco130823, w_eco130824, w_eco130825, w_eco130826, w_eco130827, w_eco130828, w_eco130829, w_eco130830, w_eco130831, w_eco130832, w_eco130833, w_eco130834, w_eco130835, w_eco130836, w_eco130837, w_eco130838, w_eco130839, w_eco130840, w_eco130841, w_eco130842, w_eco130843, w_eco130844, w_eco130845, w_eco130846, w_eco130847, w_eco130848, w_eco130849, w_eco130850, w_eco130851, w_eco130852, w_eco130853, w_eco130854, w_eco130855, w_eco130856, w_eco130857, w_eco130858, w_eco130859, w_eco130860, w_eco130861, w_eco130862, w_eco130863, w_eco130864, w_eco130865, w_eco130866, w_eco130867, w_eco130868, w_eco130869, w_eco130870, w_eco130871, w_eco130872, w_eco130873, w_eco130874, w_eco130875, w_eco130876, w_eco130877, w_eco130878, w_eco130879, w_eco130880, w_eco130881, w_eco130882, w_eco130883, w_eco130884, w_eco130885, w_eco130886, w_eco130887, w_eco130888, w_eco130889, w_eco130890, w_eco130891, w_eco130892, w_eco130893, w_eco130894, w_eco130895, w_eco130896, w_eco130897, w_eco130898, w_eco130899, w_eco130900, w_eco130901, w_eco130902, w_eco130903, w_eco130904, w_eco130905, w_eco130906, w_eco130907, w_eco130908, w_eco130909, w_eco130910, w_eco130911, w_eco130912, w_eco130913, w_eco130914, w_eco130915, w_eco130916, w_eco130917, w_eco130918, w_eco130919, w_eco130920, w_eco130921, w_eco130922, w_eco130923, w_eco130924, w_eco130925, w_eco130926, w_eco130927, w_eco130928, w_eco130929, w_eco130930, w_eco130931, w_eco130932, w_eco130933, w_eco130934, w_eco130935, w_eco130936, w_eco130937, w_eco130938, w_eco130939, w_eco130940, w_eco130941, w_eco130942, w_eco130943, w_eco130944, w_eco130945, w_eco130946, w_eco130947, w_eco130948, w_eco130949, w_eco130950, w_eco130951, w_eco130952, w_eco130953, w_eco130954, w_eco130955, w_eco130956, w_eco130957, w_eco130958, w_eco130959, w_eco130960, w_eco130961, w_eco130962, w_eco130963, w_eco130964, w_eco130965, w_eco130966, w_eco130967, w_eco130968, w_eco130969, w_eco130970, w_eco130971, w_eco130972, w_eco130973, w_eco130974, w_eco130975, w_eco130976, w_eco130977, w_eco130978, w_eco130979, w_eco130980, w_eco130981, w_eco130982, w_eco130983, w_eco130984, w_eco130985, w_eco130986, w_eco130987, w_eco130988, w_eco130989, w_eco130990, w_eco130991, w_eco130992, w_eco130993, w_eco130994, w_eco130995, w_eco130996, w_eco130997, w_eco130998, w_eco130999, w_eco131000, w_eco131001, w_eco131002, w_eco131003, w_eco131004, w_eco131005, w_eco131006, w_eco131007, w_eco131008, w_eco131009, w_eco131010, w_eco131011, w_eco131012, w_eco131013, w_eco131014, w_eco131015, w_eco131016, w_eco131017, w_eco131018, w_eco131019, w_eco131020, w_eco131021, w_eco131022, w_eco131023, w_eco131024, w_eco131025, w_eco131026, w_eco131027, w_eco131028, w_eco131029, w_eco131030, w_eco131031, w_eco131032, w_eco131033, w_eco131034, w_eco131035, w_eco131036, w_eco131037, w_eco131038, w_eco131039, w_eco131040, w_eco131041, w_eco131042, w_eco131043, w_eco131044, w_eco131045, w_eco131046, w_eco131047, w_eco131048, w_eco131049, w_eco131050, w_eco131051, w_eco131052, w_eco131053, w_eco131054, w_eco131055, w_eco131056, w_eco131057, w_eco131058, w_eco131059, w_eco131060, w_eco131061, w_eco131062, w_eco131063, w_eco131064, w_eco131065, w_eco131066, w_eco131067, w_eco131068, w_eco131069, w_eco131070, w_eco131071, w_eco131072, w_eco131073, w_eco131074, w_eco131075, w_eco131076, w_eco131077, w_eco131078, w_eco131079, w_eco131080, w_eco131081, w_eco131082, w_eco131083, w_eco131084, w_eco131085, w_eco131086, w_eco131087, w_eco131088, w_eco131089, w_eco131090, w_eco131091, w_eco131092, w_eco131093, w_eco131094, w_eco131095, w_eco131096, w_eco131097, w_eco131098, w_eco131099, w_eco131100, w_eco131101, w_eco131102, w_eco131103, w_eco131104, w_eco131105, w_eco131106, w_eco131107, w_eco131108, w_eco131109, w_eco131110, w_eco131111, w_eco131112, w_eco131113, w_eco131114, w_eco131115, w_eco131116, w_eco131117, w_eco131118, w_eco131119, w_eco131120, w_eco131121, w_eco131122, w_eco131123, w_eco131124, w_eco131125, w_eco131126, w_eco131127, w_eco131128, w_eco131129, w_eco131130, w_eco131131, w_eco131132, w_eco131133, w_eco131134, w_eco131135, w_eco131136, w_eco131137, w_eco131138, w_eco131139, w_eco131140, w_eco131141, w_eco131142, w_eco131143, w_eco131144, w_eco131145, w_eco131146, w_eco131147, w_eco131148, w_eco131149, w_eco131150, w_eco131151, w_eco131152, w_eco131153, w_eco131154, w_eco131155, w_eco131156, w_eco131157, w_eco131158, w_eco131159, w_eco131160, w_eco131161, w_eco131162, w_eco131163, w_eco131164, w_eco131165, w_eco131166, w_eco131167, w_eco131168, w_eco131169, w_eco131170, w_eco131171, w_eco131172, w_eco131173, w_eco131174, w_eco131175, w_eco131176, w_eco131177, w_eco131178, w_eco131179, w_eco131180, w_eco131181, w_eco131182, w_eco131183, w_eco131184, w_eco131185, w_eco131186, w_eco131187, w_eco131188, w_eco131189, w_eco131190, w_eco131191, w_eco131192, w_eco131193, w_eco131194, w_eco131195, w_eco131196, w_eco131197, w_eco131198, w_eco131199, w_eco131200, w_eco131201, w_eco131202, w_eco131203, w_eco131204, w_eco131205, w_eco131206, w_eco131207, w_eco131208, w_eco131209, w_eco131210, w_eco131211, w_eco131212, w_eco131213, w_eco131214, w_eco131215, w_eco131216, w_eco131217, w_eco131218, w_eco131219, w_eco131220, w_eco131221, w_eco131222, w_eco131223, w_eco131224, w_eco131225, w_eco131226, w_eco131227, w_eco131228, w_eco131229, w_eco131230, w_eco131231, w_eco131232, w_eco131233, w_eco131234, w_eco131235, w_eco131236, w_eco131237, w_eco131238, w_eco131239, w_eco131240, w_eco131241, w_eco131242, w_eco131243, w_eco131244, w_eco131245, w_eco131246, w_eco131247, w_eco131248, w_eco131249, w_eco131250, w_eco131251, w_eco131252, w_eco131253, w_eco131254, w_eco131255, w_eco131256, w_eco131257, w_eco131258, w_eco131259, w_eco131260, w_eco131261, w_eco131262, w_eco131263, w_eco131264, w_eco131265, w_eco131266, w_eco131267, w_eco131268, w_eco131269, w_eco131270, w_eco131271, w_eco131272, w_eco131273, w_eco131274, w_eco131275, w_eco131276, w_eco131277, w_eco131278, w_eco131279, w_eco131280, w_eco131281, w_eco131282, w_eco131283, w_eco131284, w_eco131285, w_eco131286, w_eco131287, w_eco131288, w_eco131289, w_eco131290, w_eco131291, w_eco131292, w_eco131293, w_eco131294, w_eco131295, w_eco131296, w_eco131297, w_eco131298, w_eco131299, w_eco131300, w_eco131301, w_eco131302, w_eco131303, w_eco131304, w_eco131305, w_eco131306, w_eco131307, w_eco131308, w_eco131309, w_eco131310, w_eco131311, w_eco131312, w_eco131313, w_eco131314, w_eco131315, w_eco131316, w_eco131317, w_eco131318, w_eco131319, w_eco131320, w_eco131321, w_eco131322, w_eco131323, w_eco131324, w_eco131325, w_eco131326, w_eco131327, w_eco131328, w_eco131329, w_eco131330, w_eco131331, w_eco131332, w_eco131333, w_eco131334, w_eco131335, w_eco131336, w_eco131337, w_eco131338, w_eco131339, w_eco131340, w_eco131341, w_eco131342, w_eco131343, w_eco131344, w_eco131345, w_eco131346, w_eco131347, w_eco131348, w_eco131349, w_eco131350, w_eco131351, w_eco131352, w_eco131353, w_eco131354, w_eco131355, w_eco131356, w_eco131357, w_eco131358, w_eco131359, w_eco131360, w_eco131361, w_eco131362, w_eco131363, w_eco131364, w_eco131365, w_eco131366, w_eco131367, w_eco131368, w_eco131369, w_eco131370, w_eco131371, w_eco131372, w_eco131373, w_eco131374, w_eco131375, w_eco131376, w_eco131377, w_eco131378, w_eco131379, w_eco131380, w_eco131381, w_eco131382, w_eco131383, w_eco131384, w_eco131385, w_eco131386, w_eco131387, w_eco131388, w_eco131389, w_eco131390, w_eco131391, w_eco131392, w_eco131393, w_eco131394, w_eco131395, w_eco131396, w_eco131397, w_eco131398, w_eco131399, w_eco131400, w_eco131401, w_eco131402, w_eco131403, w_eco131404, w_eco131405, w_eco131406, w_eco131407, w_eco131408, w_eco131409, w_eco131410, w_eco131411, w_eco131412, w_eco131413, w_eco131414, w_eco131415, w_eco131416, w_eco131417, w_eco131418, w_eco131419, w_eco131420, w_eco131421, w_eco131422, w_eco131423, w_eco131424, w_eco131425, w_eco131426, w_eco131427, w_eco131428, w_eco131429, w_eco131430, w_eco131431, w_eco131432, w_eco131433, w_eco131434, w_eco131435, w_eco131436, w_eco131437, w_eco131438, w_eco131439, w_eco131440, w_eco131441, w_eco131442, w_eco131443, w_eco131444, w_eco131445, w_eco131446, w_eco131447, w_eco131448, w_eco131449, w_eco131450, w_eco131451, w_eco131452, w_eco131453, w_eco131454, w_eco131455, w_eco131456, w_eco131457, w_eco131458, w_eco131459, w_eco131460, w_eco131461, w_eco131462, w_eco131463, w_eco131464, w_eco131465, w_eco131466, w_eco131467, w_eco131468, w_eco131469, w_eco131470, w_eco131471, w_eco131472, w_eco131473, w_eco131474, w_eco131475, w_eco131476, w_eco131477, w_eco131478, w_eco131479, w_eco131480, w_eco131481, w_eco131482, w_eco131483, w_eco131484, w_eco131485, w_eco131486, w_eco131487, w_eco131488, w_eco131489, w_eco131490, w_eco131491, w_eco131492, w_eco131493, w_eco131494, w_eco131495, w_eco131496, w_eco131497, w_eco131498, w_eco131499, w_eco131500, w_eco131501, w_eco131502, w_eco131503, w_eco131504, w_eco131505, w_eco131506, w_eco131507, w_eco131508, w_eco131509, w_eco131510, w_eco131511, w_eco131512, w_eco131513, w_eco131514, w_eco131515, w_eco131516, w_eco131517, w_eco131518, w_eco131519, w_eco131520, w_eco131521, w_eco131522, w_eco131523, w_eco131524, w_eco131525, w_eco131526, w_eco131527, w_eco131528, w_eco131529, w_eco131530, w_eco131531, w_eco131532, w_eco131533, w_eco131534, w_eco131535, w_eco131536, w_eco131537, w_eco131538, w_eco131539, w_eco131540, w_eco131541, w_eco131542, w_eco131543, w_eco131544, w_eco131545, w_eco131546, w_eco131547, w_eco131548, w_eco131549, w_eco131550, w_eco131551, w_eco131552, w_eco131553, w_eco131554, w_eco131555, w_eco131556, w_eco131557, w_eco131558, w_eco131559, w_eco131560, w_eco131561, w_eco131562, w_eco131563, w_eco131564, w_eco131565, w_eco131566, w_eco131567, w_eco131568, w_eco131569, w_eco131570, w_eco131571, w_eco131572, w_eco131573, w_eco131574, w_eco131575, w_eco131576, w_eco131577, w_eco131578, w_eco131579, w_eco131580, w_eco131581, w_eco131582, w_eco131583, w_eco131584, w_eco131585, w_eco131586, w_eco131587, w_eco131588, w_eco131589, w_eco131590, w_eco131591, w_eco131592, w_eco131593, w_eco131594, w_eco131595, w_eco131596, w_eco131597, w_eco131598, w_eco131599, w_eco131600, w_eco131601, w_eco131602, w_eco131603, w_eco131604, w_eco131605, w_eco131606, w_eco131607, w_eco131608, w_eco131609, w_eco131610, w_eco131611, w_eco131612, w_eco131613, w_eco131614, w_eco131615, w_eco131616, w_eco131617, w_eco131618, w_eco131619, w_eco131620, w_eco131621, w_eco131622, w_eco131623, w_eco131624, w_eco131625, w_eco131626, w_eco131627, w_eco131628, w_eco131629, w_eco131630, w_eco131631, w_eco131632, w_eco131633, w_eco131634, w_eco131635, w_eco131636, w_eco131637, w_eco131638, w_eco131639, w_eco131640, w_eco131641, w_eco131642, w_eco131643, w_eco131644, w_eco131645, w_eco131646, w_eco131647, w_eco131648, w_eco131649, w_eco131650, w_eco131651, w_eco131652, w_eco131653, w_eco131654, w_eco131655, w_eco131656, w_eco131657, w_eco131658, w_eco131659, w_eco131660, w_eco131661, w_eco131662, w_eco131663, w_eco131664, w_eco131665, w_eco131666, w_eco131667, w_eco131668, w_eco131669, w_eco131670, w_eco131671, w_eco131672, w_eco131673, w_eco131674, w_eco131675, w_eco131676, w_eco131677, w_eco131678, w_eco131679, w_eco131680, w_eco131681, w_eco131682, w_eco131683, w_eco131684, w_eco131685, w_eco131686, w_eco131687, w_eco131688, w_eco131689, w_eco131690, w_eco131691, w_eco131692, w_eco131693, w_eco131694, w_eco131695, w_eco131696, w_eco131697, w_eco131698, w_eco131699, w_eco131700, w_eco131701, w_eco131702, w_eco131703, w_eco131704, w_eco131705, w_eco131706, w_eco131707, w_eco131708, w_eco131709, w_eco131710, w_eco131711, w_eco131712, w_eco131713, w_eco131714, w_eco131715, w_eco131716, w_eco131717, w_eco131718, w_eco131719, w_eco131720, w_eco131721, w_eco131722, w_eco131723, w_eco131724, w_eco131725, w_eco131726, w_eco131727, w_eco131728, w_eco131729, w_eco131730, w_eco131731, w_eco131732, w_eco131733, w_eco131734, w_eco131735, w_eco131736, w_eco131737, w_eco131738, w_eco131739, w_eco131740, w_eco131741, w_eco131742, w_eco131743, w_eco131744, w_eco131745, w_eco131746, w_eco131747, w_eco131748, w_eco131749, w_eco131750, w_eco131751, w_eco131752, w_eco131753, w_eco131754, w_eco131755, w_eco131756, w_eco131757, w_eco131758, w_eco131759, w_eco131760, w_eco131761, w_eco131762, w_eco131763, w_eco131764, w_eco131765, w_eco131766, w_eco131767, w_eco131768, w_eco131769, w_eco131770, w_eco131771, w_eco131772, w_eco131773, w_eco131774, w_eco131775, w_eco131776, w_eco131777, w_eco131778, w_eco131779, w_eco131780, w_eco131781, w_eco131782, w_eco131783, w_eco131784, w_eco131785, w_eco131786, w_eco131787, w_eco131788, w_eco131789, w_eco131790, w_eco131791, w_eco131792, w_eco131793, w_eco131794, w_eco131795, w_eco131796, w_eco131797, w_eco131798, w_eco131799, w_eco131800, w_eco131801, w_eco131802, w_eco131803, w_eco131804, w_eco131805, w_eco131806, w_eco131807, w_eco131808, w_eco131809, w_eco131810, w_eco131811, w_eco131812, w_eco131813, w_eco131814, w_eco131815, w_eco131816, w_eco131817, w_eco131818, w_eco131819, w_eco131820, w_eco131821, w_eco131822, w_eco131823, w_eco131824, w_eco131825, w_eco131826, w_eco131827, w_eco131828, w_eco131829, w_eco131830, w_eco131831, w_eco131832, w_eco131833, w_eco131834, w_eco131835, w_eco131836, w_eco131837, w_eco131838, w_eco131839, w_eco131840, w_eco131841, w_eco131842, w_eco131843, w_eco131844, w_eco131845, w_eco131846, w_eco131847, w_eco131848, w_eco131849, w_eco131850, w_eco131851, w_eco131852, w_eco131853, w_eco131854, w_eco131855, w_eco131856, w_eco131857, w_eco131858, w_eco131859, w_eco131860, w_eco131861, w_eco131862, w_eco131863, w_eco131864, w_eco131865, w_eco131866, w_eco131867, w_eco131868, w_eco131869, w_eco131870, w_eco131871, w_eco131872, w_eco131873, w_eco131874, w_eco131875, w_eco131876, w_eco131877, w_eco131878, w_eco131879, w_eco131880, w_eco131881, w_eco131882, w_eco131883, w_eco131884, w_eco131885, w_eco131886, w_eco131887, w_eco131888, w_eco131889, w_eco131890, w_eco131891, w_eco131892, w_eco131893, w_eco131894, w_eco131895, w_eco131896, w_eco131897, w_eco131898, w_eco131899, w_eco131900, w_eco131901, w_eco131902, w_eco131903, w_eco131904, w_eco131905, w_eco131906, w_eco131907, w_eco131908, w_eco131909, w_eco131910, w_eco131911, w_eco131912, w_eco131913, w_eco131914, w_eco131915, w_eco131916, w_eco131917, w_eco131918, w_eco131919, w_eco131920, w_eco131921, w_eco131922, w_eco131923, w_eco131924, w_eco131925, w_eco131926, w_eco131927, w_eco131928, w_eco131929, w_eco131930, w_eco131931, w_eco131932, w_eco131933, w_eco131934, w_eco131935, w_eco131936, w_eco131937, w_eco131938, w_eco131939, w_eco131940, w_eco131941, w_eco131942, w_eco131943, w_eco131944, w_eco131945, w_eco131946, w_eco131947, w_eco131948, w_eco131949, w_eco131950, w_eco131951, w_eco131952, w_eco131953, w_eco131954, w_eco131955, w_eco131956, w_eco131957, w_eco131958, w_eco131959, w_eco131960, w_eco131961, w_eco131962, w_eco131963, w_eco131964, w_eco131965, w_eco131966, w_eco131967, w_eco131968, w_eco131969, w_eco131970, w_eco131971, w_eco131972, w_eco131973, w_eco131974, w_eco131975, w_eco131976, w_eco131977, w_eco131978, w_eco131979, w_eco131980, w_eco131981, w_eco131982, w_eco131983, w_eco131984, w_eco131985, w_eco131986, w_eco131987, w_eco131988, w_eco131989, w_eco131990, w_eco131991, w_eco131992, w_eco131993, w_eco131994, w_eco131995, w_eco131996, w_eco131997, w_eco131998, w_eco131999, w_eco132000, w_eco132001, w_eco132002, w_eco132003, w_eco132004, w_eco132005, w_eco132006, w_eco132007, w_eco132008, w_eco132009, w_eco132010, w_eco132011, w_eco132012, w_eco132013, w_eco132014, w_eco132015, w_eco132016, w_eco132017, w_eco132018, w_eco132019, w_eco132020, w_eco132021, w_eco132022, w_eco132023, w_eco132024, w_eco132025, w_eco132026, w_eco132027, w_eco132028, w_eco132029, w_eco132030, w_eco132031, w_eco132032, w_eco132033, w_eco132034, w_eco132035, w_eco132036, w_eco132037, w_eco132038, w_eco132039, w_eco132040, w_eco132041, w_eco132042, w_eco132043, w_eco132044, w_eco132045, w_eco132046, w_eco132047, w_eco132048, w_eco132049, w_eco132050, w_eco132051, w_eco132052, w_eco132053, w_eco132054, w_eco132055, w_eco132056, w_eco132057, w_eco132058, w_eco132059, w_eco132060, w_eco132061, w_eco132062, w_eco132063, w_eco132064, w_eco132065, w_eco132066, w_eco132067, w_eco132068, w_eco132069, w_eco132070, w_eco132071, w_eco132072, w_eco132073, w_eco132074, w_eco132075, w_eco132076, w_eco132077, w_eco132078, w_eco132079, w_eco132080, w_eco132081, w_eco132082, w_eco132083, w_eco132084, w_eco132085, w_eco132086, w_eco132087, w_eco132088, w_eco132089, w_eco132090, w_eco132091, w_eco132092, w_eco132093, w_eco132094, w_eco132095, w_eco132096, w_eco132097, w_eco132098, w_eco132099, w_eco132100, w_eco132101, w_eco132102, w_eco132103, w_eco132104, w_eco132105, w_eco132106, w_eco132107, w_eco132108, w_eco132109, w_eco132110, w_eco132111, w_eco132112, w_eco132113, w_eco132114, w_eco132115, w_eco132116, w_eco132117, w_eco132118, w_eco132119, w_eco132120, w_eco132121, w_eco132122, w_eco132123, w_eco132124, w_eco132125, w_eco132126, w_eco132127, w_eco132128, w_eco132129, w_eco132130, w_eco132131, w_eco132132, w_eco132133, w_eco132134, w_eco132135, w_eco132136, w_eco132137, w_eco132138, w_eco132139, w_eco132140, w_eco132141, w_eco132142, w_eco132143, w_eco132144, w_eco132145, w_eco132146, w_eco132147, w_eco132148, w_eco132149, w_eco132150, w_eco132151, w_eco132152, w_eco132153, w_eco132154, w_eco132155, w_eco132156, w_eco132157, w_eco132158, w_eco132159, w_eco132160, w_eco132161, w_eco132162, w_eco132163, w_eco132164, w_eco132165, w_eco132166, w_eco132167, w_eco132168, w_eco132169, w_eco132170, w_eco132171, w_eco132172, w_eco132173, w_eco132174, w_eco132175, w_eco132176, w_eco132177, w_eco132178, w_eco132179, w_eco132180, w_eco132181, w_eco132182, w_eco132183, w_eco132184, w_eco132185, w_eco132186, w_eco132187, w_eco132188, w_eco132189, w_eco132190, w_eco132191, w_eco132192, w_eco132193, w_eco132194, w_eco132195, w_eco132196, w_eco132197, w_eco132198, w_eco132199, w_eco132200, w_eco132201, w_eco132202, w_eco132203, w_eco132204, w_eco132205, w_eco132206, w_eco132207, w_eco132208, w_eco132209, w_eco132210, w_eco132211, w_eco132212, w_eco132213, w_eco132214, w_eco132215, w_eco132216, w_eco132217, w_eco132218, w_eco132219, w_eco132220, w_eco132221, w_eco132222, w_eco132223, w_eco132224, w_eco132225, w_eco132226, w_eco132227, w_eco132228, w_eco132229, w_eco132230, w_eco132231, w_eco132232, w_eco132233, w_eco132234, w_eco132235, w_eco132236, w_eco132237, w_eco132238, w_eco132239, w_eco132240, w_eco132241, w_eco132242, w_eco132243, w_eco132244, w_eco132245, w_eco132246, w_eco132247, w_eco132248, w_eco132249, w_eco132250, w_eco132251, w_eco132252, w_eco132253, w_eco132254, w_eco132255, w_eco132256, w_eco132257, w_eco132258, w_eco132259, w_eco132260, w_eco132261, w_eco132262, w_eco132263, w_eco132264, w_eco132265, w_eco132266, w_eco132267, w_eco132268, w_eco132269, w_eco132270, w_eco132271, w_eco132272, w_eco132273, w_eco132274, w_eco132275, w_eco132276, w_eco132277, w_eco132278, w_eco132279, w_eco132280, w_eco132281, w_eco132282, w_eco132283, w_eco132284, w_eco132285, w_eco132286, w_eco132287, w_eco132288, w_eco132289, w_eco132290, w_eco132291, w_eco132292, w_eco132293, w_eco132294, w_eco132295, w_eco132296, w_eco132297, w_eco132298, w_eco132299, w_eco132300, w_eco132301, w_eco132302, w_eco132303, w_eco132304, w_eco132305, w_eco132306, w_eco132307, w_eco132308, w_eco132309, w_eco132310, w_eco132311, w_eco132312, w_eco132313, w_eco132314, w_eco132315, w_eco132316, w_eco132317, w_eco132318, w_eco132319, w_eco132320, w_eco132321, w_eco132322, w_eco132323, w_eco132324, w_eco132325, w_eco132326, w_eco132327, w_eco132328, w_eco132329, w_eco132330, w_eco132331, w_eco132332, w_eco132333, w_eco132334, w_eco132335, w_eco132336, w_eco132337, w_eco132338, w_eco132339, w_eco132340, w_eco132341, w_eco132342, w_eco132343, w_eco132344, w_eco132345, w_eco132346, w_eco132347, w_eco132348, w_eco132349, w_eco132350, w_eco132351, w_eco132352, w_eco132353, w_eco132354, w_eco132355, w_eco132356, w_eco132357, w_eco132358, w_eco132359, w_eco132360, w_eco132361, w_eco132362, w_eco132363, w_eco132364, w_eco132365, w_eco132366, w_eco132367, w_eco132368, w_eco132369, w_eco132370, w_eco132371, w_eco132372, w_eco132373, w_eco132374, w_eco132375, w_eco132376, w_eco132377, w_eco132378, w_eco132379, w_eco132380, w_eco132381, w_eco132382, w_eco132383, w_eco132384, w_eco132385, w_eco132386, w_eco132387, w_eco132388, w_eco132389, w_eco132390, w_eco132391, w_eco132392, w_eco132393, w_eco132394, w_eco132395, w_eco132396, w_eco132397, w_eco132398, w_eco132399, w_eco132400, w_eco132401, w_eco132402, w_eco132403, w_eco132404, w_eco132405, w_eco132406, w_eco132407, w_eco132408, w_eco132409, w_eco132410, w_eco132411, w_eco132412, w_eco132413, w_eco132414, w_eco132415, w_eco132416, w_eco132417, w_eco132418, w_eco132419, w_eco132420, w_eco132421, w_eco132422, w_eco132423, w_eco132424, w_eco132425, w_eco132426, w_eco132427, w_eco132428, w_eco132429, w_eco132430, w_eco132431, w_eco132432, w_eco132433, w_eco132434, w_eco132435, w_eco132436, w_eco132437, w_eco132438, w_eco132439, w_eco132440, w_eco132441, w_eco132442, w_eco132443, w_eco132444, w_eco132445, w_eco132446, w_eco132447, w_eco132448, w_eco132449, w_eco132450, w_eco132451, w_eco132452, w_eco132453, w_eco132454, w_eco132455, w_eco132456, w_eco132457, w_eco132458, w_eco132459, w_eco132460, w_eco132461, w_eco132462, w_eco132463, w_eco132464, w_eco132465, w_eco132466, w_eco132467, w_eco132468, w_eco132469, w_eco132470, w_eco132471, w_eco132472, w_eco132473, w_eco132474, w_eco132475, w_eco132476, w_eco132477, w_eco132478, w_eco132479, w_eco132480, w_eco132481, w_eco132482, w_eco132483, w_eco132484, w_eco132485, w_eco132486, w_eco132487, w_eco132488, w_eco132489, w_eco132490, w_eco132491, w_eco132492, w_eco132493, w_eco132494, w_eco132495, w_eco132496, w_eco132497, w_eco132498, w_eco132499, w_eco132500, w_eco132501, w_eco132502, w_eco132503, w_eco132504, w_eco132505, w_eco132506, w_eco132507, w_eco132508, w_eco132509, w_eco132510, w_eco132511, w_eco132512, w_eco132513, w_eco132514, w_eco132515, w_eco132516, w_eco132517, w_eco132518, w_eco132519, w_eco132520, w_eco132521, w_eco132522, w_eco132523, w_eco132524, w_eco132525, w_eco132526, w_eco132527, w_eco132528, w_eco132529, w_eco132530, w_eco132531, w_eco132532, w_eco132533, w_eco132534, w_eco132535, w_eco132536, w_eco132537, w_eco132538, w_eco132539, w_eco132540, w_eco132541, w_eco132542, w_eco132543, w_eco132544, w_eco132545, w_eco132546, w_eco132547, w_eco132548, w_eco132549, w_eco132550, w_eco132551, w_eco132552, w_eco132553, w_eco132554, w_eco132555, w_eco132556, w_eco132557, w_eco132558, w_eco132559, w_eco132560, w_eco132561, w_eco132562, w_eco132563, w_eco132564, w_eco132565, w_eco132566, w_eco132567, w_eco132568, w_eco132569, w_eco132570, w_eco132571, w_eco132572, w_eco132573, w_eco132574, w_eco132575, w_eco132576, w_eco132577, w_eco132578, w_eco132579, w_eco132580, w_eco132581, w_eco132582, w_eco132583, w_eco132584, w_eco132585, w_eco132586, w_eco132587, w_eco132588, w_eco132589, w_eco132590, w_eco132591, w_eco132592, w_eco132593, w_eco132594, w_eco132595, w_eco132596, w_eco132597, w_eco132598, w_eco132599, w_eco132600, w_eco132601, w_eco132602, w_eco132603, w_eco132604, w_eco132605, w_eco132606, w_eco132607, w_eco132608, w_eco132609, w_eco132610, w_eco132611, w_eco132612, w_eco132613, w_eco132614, w_eco132615, w_eco132616, w_eco132617, w_eco132618, w_eco132619, w_eco132620, w_eco132621, w_eco132622, w_eco132623, w_eco132624, w_eco132625, w_eco132626, w_eco132627, w_eco132628, w_eco132629, w_eco132630, w_eco132631, w_eco132632, w_eco132633, w_eco132634, w_eco132635, w_eco132636, w_eco132637, w_eco132638, w_eco132639, w_eco132640, w_eco132641, w_eco132642, w_eco132643, w_eco132644, w_eco132645, w_eco132646, w_eco132647, w_eco132648, w_eco132649, w_eco132650, w_eco132651, w_eco132652, w_eco132653, w_eco132654, w_eco132655, w_eco132656, w_eco132657, w_eco132658, w_eco132659, w_eco132660, w_eco132661, w_eco132662, w_eco132663, w_eco132664, w_eco132665, w_eco132666, w_eco132667, w_eco132668, w_eco132669, w_eco132670, w_eco132671, w_eco132672, w_eco132673, w_eco132674, w_eco132675, w_eco132676, w_eco132677, w_eco132678, w_eco132679, w_eco132680, w_eco132681, w_eco132682, w_eco132683, w_eco132684, w_eco132685, w_eco132686, w_eco132687, w_eco132688, w_eco132689, w_eco132690, w_eco132691, w_eco132692, w_eco132693, w_eco132694, w_eco132695, w_eco132696, w_eco132697, w_eco132698, w_eco132699, w_eco132700, w_eco132701, w_eco132702, w_eco132703, w_eco132704, w_eco132705, w_eco132706, w_eco132707, w_eco132708, w_eco132709, w_eco132710, w_eco132711, w_eco132712, w_eco132713, w_eco132714, w_eco132715, w_eco132716, w_eco132717, w_eco132718, w_eco132719, w_eco132720, w_eco132721, w_eco132722, w_eco132723, w_eco132724, w_eco132725, w_eco132726, w_eco132727, w_eco132728, w_eco132729, w_eco132730, w_eco132731, w_eco132732, w_eco132733, w_eco132734, w_eco132735, w_eco132736, w_eco132737, w_eco132738, w_eco132739, w_eco132740, w_eco132741, w_eco132742, w_eco132743, w_eco132744, w_eco132745, w_eco132746, w_eco132747, w_eco132748, w_eco132749, w_eco132750, w_eco132751, w_eco132752, w_eco132753, w_eco132754, w_eco132755, w_eco132756, w_eco132757, w_eco132758, w_eco132759, w_eco132760, w_eco132761, w_eco132762, w_eco132763, w_eco132764, w_eco132765, w_eco132766, w_eco132767, w_eco132768, w_eco132769, w_eco132770, w_eco132771, w_eco132772, w_eco132773, w_eco132774, w_eco132775, w_eco132776, w_eco132777, w_eco132778, w_eco132779, w_eco132780, w_eco132781, w_eco132782, w_eco132783, w_eco132784, w_eco132785, w_eco132786, w_eco132787, w_eco132788, w_eco132789, w_eco132790, w_eco132791, w_eco132792, w_eco132793, w_eco132794, w_eco132795, w_eco132796, w_eco132797, w_eco132798, w_eco132799, w_eco132800, w_eco132801, w_eco132802, w_eco132803, w_eco132804, w_eco132805, w_eco132806, w_eco132807, w_eco132808, w_eco132809, w_eco132810, w_eco132811, w_eco132812, w_eco132813, w_eco132814, w_eco132815, w_eco132816, w_eco132817, w_eco132818, w_eco132819, w_eco132820, w_eco132821, w_eco132822, w_eco132823, w_eco132824, w_eco132825, w_eco132826, w_eco132827, w_eco132828, w_eco132829, w_eco132830, w_eco132831, w_eco132832, w_eco132833, w_eco132834, w_eco132835, w_eco132836, w_eco132837, w_eco132838, w_eco132839, w_eco132840, w_eco132841, w_eco132842, w_eco132843, w_eco132844, w_eco132845, w_eco132846, w_eco132847, w_eco132848, w_eco132849, w_eco132850, w_eco132851, w_eco132852, w_eco132853, w_eco132854, w_eco132855, w_eco132856, w_eco132857, w_eco132858, w_eco132859, w_eco132860, w_eco132861, w_eco132862, w_eco132863, w_eco132864, w_eco132865, w_eco132866, w_eco132867, w_eco132868, w_eco132869, w_eco132870, w_eco132871, w_eco132872, w_eco132873, w_eco132874, w_eco132875, w_eco132876, w_eco132877, w_eco132878, w_eco132879, w_eco132880, w_eco132881, w_eco132882, w_eco132883, w_eco132884, w_eco132885, w_eco132886, w_eco132887, w_eco132888, w_eco132889, w_eco132890, w_eco132891, w_eco132892, w_eco132893, w_eco132894, w_eco132895, w_eco132896, w_eco132897, w_eco132898, w_eco132899, w_eco132900, w_eco132901, w_eco132902, w_eco132903, w_eco132904, w_eco132905, w_eco132906, w_eco132907, w_eco132908, w_eco132909, w_eco132910, w_eco132911, w_eco132912, w_eco132913, w_eco132914, w_eco132915, w_eco132916, w_eco132917, w_eco132918, w_eco132919, w_eco132920, w_eco132921, w_eco132922, w_eco132923, w_eco132924, w_eco132925, w_eco132926, w_eco132927, w_eco132928, w_eco132929, w_eco132930, w_eco132931, w_eco132932, w_eco132933, w_eco132934, w_eco132935, w_eco132936, w_eco132937, w_eco132938, w_eco132939, w_eco132940, w_eco132941, w_eco132942, w_eco132943, w_eco132944, w_eco132945, w_eco132946, w_eco132947, w_eco132948, w_eco132949, w_eco132950, w_eco132951, w_eco132952, w_eco132953, w_eco132954, w_eco132955, w_eco132956, w_eco132957, w_eco132958, w_eco132959, w_eco132960, w_eco132961, w_eco132962, w_eco132963, w_eco132964, w_eco132965, w_eco132966, w_eco132967, w_eco132968, w_eco132969, w_eco132970, w_eco132971, w_eco132972, w_eco132973, w_eco132974, w_eco132975, w_eco132976, w_eco132977, w_eco132978, w_eco132979, w_eco132980, w_eco132981, w_eco132982, w_eco132983, w_eco132984, w_eco132985, w_eco132986, w_eco132987, w_eco132988, w_eco132989, w_eco132990, w_eco132991, w_eco132992, w_eco132993, w_eco132994, w_eco132995, w_eco132996, w_eco132997, w_eco132998, w_eco132999, w_eco133000, w_eco133001, w_eco133002, w_eco133003, w_eco133004, w_eco133005, w_eco133006, w_eco133007, w_eco133008, w_eco133009, w_eco133010, w_eco133011, w_eco133012, w_eco133013, w_eco133014, w_eco133015, w_eco133016, w_eco133017, w_eco133018, w_eco133019, w_eco133020, w_eco133021, w_eco133022, w_eco133023, w_eco133024, w_eco133025, w_eco133026, w_eco133027, w_eco133028, w_eco133029, w_eco133030, w_eco133031, w_eco133032, w_eco133033, w_eco133034, w_eco133035, w_eco133036, w_eco133037, w_eco133038, w_eco133039, w_eco133040, w_eco133041, w_eco133042, w_eco133043, w_eco133044, w_eco133045, w_eco133046, w_eco133047, w_eco133048, w_eco133049, w_eco133050, w_eco133051, w_eco133052, w_eco133053, w_eco133054, w_eco133055, w_eco133056, w_eco133057, w_eco133058, w_eco133059, w_eco133060, w_eco133061, w_eco133062, w_eco133063, w_eco133064, w_eco133065, w_eco133066, w_eco133067, w_eco133068, w_eco133069, w_eco133070, w_eco133071, w_eco133072, w_eco133073, w_eco133074, w_eco133075, w_eco133076, w_eco133077, w_eco133078, w_eco133079, w_eco133080, w_eco133081, w_eco133082, w_eco133083, w_eco133084, w_eco133085, w_eco133086, w_eco133087, w_eco133088, w_eco133089, w_eco133090, w_eco133091, w_eco133092, w_eco133093, w_eco133094, w_eco133095, w_eco133096, w_eco133097, w_eco133098, w_eco133099, w_eco133100, w_eco133101, w_eco133102, w_eco133103, w_eco133104, w_eco133105, w_eco133106, w_eco133107, w_eco133108, w_eco133109, w_eco133110, w_eco133111, w_eco133112, w_eco133113, w_eco133114, w_eco133115, w_eco133116, w_eco133117, w_eco133118, w_eco133119, w_eco133120, w_eco133121, w_eco133122, w_eco133123, w_eco133124, w_eco133125, w_eco133126, w_eco133127, w_eco133128, w_eco133129, w_eco133130, w_eco133131, w_eco133132, w_eco133133, w_eco133134, w_eco133135, w_eco133136, w_eco133137, w_eco133138, w_eco133139, w_eco133140, w_eco133141, w_eco133142, w_eco133143, w_eco133144, w_eco133145, w_eco133146, w_eco133147, w_eco133148, w_eco133149, w_eco133150, w_eco133151, w_eco133152, w_eco133153, w_eco133154, w_eco133155, w_eco133156, w_eco133157, w_eco133158, w_eco133159, w_eco133160, w_eco133161, w_eco133162, w_eco133163, w_eco133164, w_eco133165, w_eco133166, w_eco133167, w_eco133168, w_eco133169, w_eco133170, w_eco133171, w_eco133172, w_eco133173, w_eco133174, w_eco133175, w_eco133176, w_eco133177, w_eco133178, w_eco133179, w_eco133180, w_eco133181, w_eco133182, w_eco133183, w_eco133184, w_eco133185, w_eco133186, w_eco133187, w_eco133188, w_eco133189, w_eco133190, w_eco133191, w_eco133192, w_eco133193, w_eco133194, w_eco133195, w_eco133196, w_eco133197, w_eco133198, w_eco133199, w_eco133200, w_eco133201, w_eco133202, w_eco133203, w_eco133204, w_eco133205, w_eco133206, w_eco133207, w_eco133208, w_eco133209, w_eco133210, w_eco133211, w_eco133212, w_eco133213, w_eco133214, w_eco133215, w_eco133216, w_eco133217, w_eco133218, w_eco133219, w_eco133220, w_eco133221, w_eco133222, w_eco133223, w_eco133224, w_eco133225, w_eco133226, w_eco133227, w_eco133228, w_eco133229, w_eco133230, w_eco133231, w_eco133232, w_eco133233, w_eco133234, w_eco133235, w_eco133236, w_eco133237, w_eco133238, w_eco133239, w_eco133240, w_eco133241, w_eco133242, w_eco133243, w_eco133244, w_eco133245, w_eco133246, w_eco133247, w_eco133248, w_eco133249, w_eco133250, w_eco133251, w_eco133252, w_eco133253, w_eco133254, w_eco133255, w_eco133256, w_eco133257, w_eco133258, w_eco133259, w_eco133260, w_eco133261, w_eco133262, w_eco133263, w_eco133264, w_eco133265, w_eco133266, w_eco133267, w_eco133268, w_eco133269, w_eco133270, w_eco133271, w_eco133272, w_eco133273, w_eco133274, w_eco133275, w_eco133276, w_eco133277, w_eco133278, w_eco133279, w_eco133280, w_eco133281, w_eco133282, w_eco133283, w_eco133284, w_eco133285, w_eco133286, w_eco133287, w_eco133288, w_eco133289, w_eco133290, w_eco133291, w_eco133292, w_eco133293, w_eco133294, w_eco133295, w_eco133296, w_eco133297, w_eco133298, w_eco133299, w_eco133300, w_eco133301, w_eco133302, w_eco133303, w_eco133304, w_eco133305, w_eco133306, w_eco133307, w_eco133308, w_eco133309, w_eco133310, w_eco133311, w_eco133312, w_eco133313, w_eco133314, w_eco133315, w_eco133316, w_eco133317, w_eco133318, w_eco133319, w_eco133320, w_eco133321, w_eco133322, w_eco133323, w_eco133324, w_eco133325, w_eco133326, w_eco133327, w_eco133328, w_eco133329, w_eco133330, w_eco133331, w_eco133332, w_eco133333, w_eco133334, w_eco133335, w_eco133336, w_eco133337, w_eco133338, w_eco133339, w_eco133340, w_eco133341, w_eco133342, w_eco133343, w_eco133344, w_eco133345, w_eco133346, w_eco133347, w_eco133348, w_eco133349, w_eco133350, w_eco133351, w_eco133352, w_eco133353, w_eco133354, w_eco133355, w_eco133356, w_eco133357, w_eco133358, w_eco133359, w_eco133360, w_eco133361, w_eco133362, w_eco133363, w_eco133364, w_eco133365, w_eco133366, w_eco133367, w_eco133368, w_eco133369, w_eco133370, w_eco133371, w_eco133372, w_eco133373, w_eco133374, w_eco133375, w_eco133376, w_eco133377, w_eco133378, w_eco133379, w_eco133380, w_eco133381, w_eco133382, w_eco133383, w_eco133384, w_eco133385, w_eco133386, w_eco133387, w_eco133388, w_eco133389, w_eco133390, w_eco133391, w_eco133392, w_eco133393, w_eco133394, w_eco133395, w_eco133396, w_eco133397, w_eco133398, w_eco133399, w_eco133400, w_eco133401, w_eco133402, w_eco133403, w_eco133404, w_eco133405, w_eco133406, w_eco133407, w_eco133408, w_eco133409, w_eco133410, w_eco133411, w_eco133412, w_eco133413, w_eco133414, w_eco133415, w_eco133416, w_eco133417, w_eco133418, w_eco133419, w_eco133420, w_eco133421, w_eco133422, w_eco133423, w_eco133424, w_eco133425, w_eco133426, w_eco133427, w_eco133428, w_eco133429, w_eco133430, w_eco133431, w_eco133432, w_eco133433, w_eco133434, w_eco133435, w_eco133436, w_eco133437, w_eco133438, w_eco133439, w_eco133440, w_eco133441, w_eco133442, w_eco133443, w_eco133444, w_eco133445, w_eco133446, w_eco133447, w_eco133448, w_eco133449, w_eco133450, w_eco133451, w_eco133452, w_eco133453, w_eco133454, w_eco133455, w_eco133456, w_eco133457, w_eco133458, w_eco133459, w_eco133460, w_eco133461, w_eco133462, w_eco133463, w_eco133464, w_eco133465, w_eco133466, w_eco133467, w_eco133468, w_eco133469, w_eco133470, w_eco133471, w_eco133472, w_eco133473, w_eco133474, w_eco133475, w_eco133476, w_eco133477, w_eco133478, w_eco133479, w_eco133480, w_eco133481, w_eco133482, w_eco133483, w_eco133484, w_eco133485, w_eco133486, w_eco133487, w_eco133488, w_eco133489, w_eco133490, w_eco133491, w_eco133492, w_eco133493, w_eco133494, w_eco133495, w_eco133496, w_eco133497, w_eco133498, w_eco133499, w_eco133500, w_eco133501, w_eco133502, w_eco133503, w_eco133504, w_eco133505, w_eco133506, w_eco133507, w_eco133508, w_eco133509, w_eco133510, w_eco133511, w_eco133512, w_eco133513, w_eco133514, w_eco133515, w_eco133516, w_eco133517, w_eco133518, w_eco133519, w_eco133520, w_eco133521, w_eco133522, w_eco133523, w_eco133524, w_eco133525, w_eco133526, w_eco133527, w_eco133528, w_eco133529, w_eco133530, w_eco133531, w_eco133532, w_eco133533, w_eco133534, w_eco133535, w_eco133536, w_eco133537, w_eco133538, w_eco133539, w_eco133540, w_eco133541, w_eco133542, w_eco133543, w_eco133544, w_eco133545, w_eco133546, w_eco133547, w_eco133548, w_eco133549, w_eco133550, w_eco133551, w_eco133552, w_eco133553, w_eco133554, w_eco133555, w_eco133556, w_eco133557, w_eco133558, w_eco133559, w_eco133560, w_eco133561, w_eco133562, w_eco133563, w_eco133564, w_eco133565, w_eco133566, w_eco133567, w_eco133568, w_eco133569, w_eco133570, w_eco133571, w_eco133572, w_eco133573, w_eco133574, w_eco133575, w_eco133576, w_eco133577, w_eco133578, w_eco133579, w_eco133580, w_eco133581, w_eco133582, w_eco133583, w_eco133584, w_eco133585, w_eco133586, w_eco133587, w_eco133588, w_eco133589, w_eco133590, w_eco133591, w_eco133592, w_eco133593, w_eco133594, w_eco133595, w_eco133596, w_eco133597, w_eco133598, w_eco133599, w_eco133600, w_eco133601, w_eco133602, w_eco133603, w_eco133604, w_eco133605, w_eco133606, w_eco133607, w_eco133608, w_eco133609, w_eco133610, w_eco133611, w_eco133612, w_eco133613, w_eco133614, w_eco133615, w_eco133616, w_eco133617, w_eco133618, w_eco133619, w_eco133620, w_eco133621, w_eco133622, w_eco133623, w_eco133624, w_eco133625, w_eco133626, w_eco133627, w_eco133628, w_eco133629, w_eco133630, w_eco133631, w_eco133632, w_eco133633, w_eco133634, w_eco133635, w_eco133636, w_eco133637, w_eco133638, w_eco133639, w_eco133640, w_eco133641, w_eco133642, w_eco133643, w_eco133644, w_eco133645, w_eco133646, w_eco133647, w_eco133648, w_eco133649, w_eco133650, w_eco133651, w_eco133652, w_eco133653, w_eco133654, w_eco133655, w_eco133656, w_eco133657, w_eco133658, w_eco133659, w_eco133660, w_eco133661, w_eco133662, w_eco133663, w_eco133664, w_eco133665, w_eco133666, w_eco133667, w_eco133668, w_eco133669, w_eco133670, w_eco133671, w_eco133672, w_eco133673, w_eco133674, w_eco133675, w_eco133676, w_eco133677, w_eco133678, w_eco133679, w_eco133680, w_eco133681, w_eco133682, w_eco133683, w_eco133684, w_eco133685, w_eco133686, w_eco133687, w_eco133688, w_eco133689, w_eco133690, w_eco133691, w_eco133692, w_eco133693, w_eco133694, w_eco133695, w_eco133696, w_eco133697, w_eco133698, w_eco133699, w_eco133700, w_eco133701, w_eco133702, w_eco133703, w_eco133704, w_eco133705, w_eco133706, w_eco133707, w_eco133708, w_eco133709, w_eco133710, w_eco133711, w_eco133712, w_eco133713, w_eco133714, w_eco133715, w_eco133716, w_eco133717, w_eco133718, w_eco133719, w_eco133720, w_eco133721, w_eco133722, w_eco133723, w_eco133724, w_eco133725, w_eco133726, w_eco133727, w_eco133728, w_eco133729, w_eco133730, w_eco133731, w_eco133732, w_eco133733, w_eco133734, w_eco133735, w_eco133736, w_eco133737, w_eco133738, w_eco133739, w_eco133740, w_eco133741, w_eco133742, w_eco133743, w_eco133744, w_eco133745, w_eco133746, w_eco133747, w_eco133748, w_eco133749, w_eco133750, w_eco133751, w_eco133752, w_eco133753, w_eco133754, w_eco133755, w_eco133756, w_eco133757, w_eco133758, w_eco133759, w_eco133760, w_eco133761, w_eco133762, w_eco133763, w_eco133764, w_eco133765, w_eco133766, w_eco133767, w_eco133768, w_eco133769, w_eco133770, w_eco133771, w_eco133772, w_eco133773, w_eco133774, w_eco133775, w_eco133776, w_eco133777, w_eco133778, w_eco133779, w_eco133780, w_eco133781, w_eco133782, w_eco133783, w_eco133784, w_eco133785, w_eco133786, w_eco133787, w_eco133788, w_eco133789, w_eco133790, w_eco133791, w_eco133792, w_eco133793, w_eco133794, w_eco133795, w_eco133796, w_eco133797, w_eco133798, w_eco133799, w_eco133800, w_eco133801, w_eco133802, w_eco133803, w_eco133804, w_eco133805, w_eco133806, w_eco133807, w_eco133808, w_eco133809, w_eco133810, w_eco133811, w_eco133812, w_eco133813, w_eco133814, w_eco133815, w_eco133816, w_eco133817, w_eco133818, w_eco133819, w_eco133820, w_eco133821, w_eco133822, w_eco133823, w_eco133824, w_eco133825, w_eco133826, w_eco133827, w_eco133828, w_eco133829, w_eco133830, w_eco133831, w_eco133832, w_eco133833, w_eco133834, w_eco133835, w_eco133836, w_eco133837, w_eco133838, w_eco133839, w_eco133840, w_eco133841, w_eco133842, w_eco133843, w_eco133844, w_eco133845, w_eco133846, w_eco133847, w_eco133848, w_eco133849, w_eco133850, w_eco133851, w_eco133852, w_eco133853, w_eco133854, w_eco133855, w_eco133856, w_eco133857, w_eco133858, w_eco133859, w_eco133860, w_eco133861, w_eco133862, w_eco133863, w_eco133864, w_eco133865, w_eco133866, w_eco133867, w_eco133868, w_eco133869, w_eco133870, w_eco133871, w_eco133872, w_eco133873, w_eco133874, w_eco133875, w_eco133876, w_eco133877, w_eco133878, w_eco133879, w_eco133880, w_eco133881, w_eco133882, w_eco133883, w_eco133884, w_eco133885, w_eco133886, w_eco133887, w_eco133888, w_eco133889, w_eco133890, w_eco133891, w_eco133892, w_eco133893, w_eco133894, w_eco133895, w_eco133896, w_eco133897, w_eco133898, w_eco133899, w_eco133900, w_eco133901, w_eco133902, w_eco133903, w_eco133904, w_eco133905, w_eco133906, w_eco133907, w_eco133908, w_eco133909, w_eco133910, w_eco133911, w_eco133912, w_eco133913, w_eco133914, w_eco133915, w_eco133916, w_eco133917, w_eco133918, w_eco133919, w_eco133920, w_eco133921, w_eco133922, w_eco133923, w_eco133924, w_eco133925, w_eco133926, w_eco133927, w_eco133928, w_eco133929, w_eco133930, w_eco133931, w_eco133932, w_eco133933, w_eco133934, w_eco133935, w_eco133936, w_eco133937, w_eco133938, w_eco133939, w_eco133940, w_eco133941, w_eco133942, w_eco133943, w_eco133944, w_eco133945, w_eco133946, w_eco133947, w_eco133948, w_eco133949, w_eco133950, w_eco133951, w_eco133952, w_eco133953, w_eco133954, w_eco133955, w_eco133956, w_eco133957, w_eco133958, w_eco133959, w_eco133960, w_eco133961, w_eco133962, w_eco133963, w_eco133964, w_eco133965, w_eco133966, w_eco133967, w_eco133968, w_eco133969, w_eco133970, w_eco133971, w_eco133972, w_eco133973, w_eco133974, w_eco133975, w_eco133976, w_eco133977, w_eco133978, w_eco133979, w_eco133980, w_eco133981, w_eco133982, w_eco133983, w_eco133984, w_eco133985, w_eco133986, w_eco133987, w_eco133988, w_eco133989, w_eco133990, w_eco133991, w_eco133992, w_eco133993, w_eco133994, w_eco133995, w_eco133996, w_eco133997, w_eco133998, w_eco133999, w_eco134000, w_eco134001, w_eco134002, w_eco134003, w_eco134004, w_eco134005, w_eco134006, w_eco134007, w_eco134008, w_eco134009, w_eco134010, w_eco134011, w_eco134012, w_eco134013, w_eco134014, w_eco134015, w_eco134016, w_eco134017, w_eco134018, w_eco134019, w_eco134020, w_eco134021, w_eco134022, w_eco134023, w_eco134024, w_eco134025, w_eco134026, w_eco134027, w_eco134028, w_eco134029, w_eco134030, w_eco134031, w_eco134032, w_eco134033, w_eco134034, w_eco134035, w_eco134036, w_eco134037, w_eco134038, w_eco134039, w_eco134040, w_eco134041, w_eco134042, w_eco134043, w_eco134044, w_eco134045, w_eco134046, w_eco134047, w_eco134048, w_eco134049, w_eco134050, w_eco134051, w_eco134052, w_eco134053, w_eco134054, w_eco134055, w_eco134056, w_eco134057, w_eco134058, w_eco134059, w_eco134060, w_eco134061, w_eco134062, w_eco134063, w_eco134064, w_eco134065, w_eco134066, w_eco134067, w_eco134068, w_eco134069, w_eco134070, w_eco134071, w_eco134072, w_eco134073, w_eco134074, w_eco134075, w_eco134076, w_eco134077, w_eco134078, w_eco134079, w_eco134080, w_eco134081, w_eco134082, w_eco134083, w_eco134084, w_eco134085, w_eco134086, w_eco134087, w_eco134088, w_eco134089, w_eco134090, w_eco134091, w_eco134092, w_eco134093, w_eco134094, w_eco134095, w_eco134096, w_eco134097, w_eco134098, w_eco134099, w_eco134100, w_eco134101, w_eco134102, w_eco134103, w_eco134104, w_eco134105, w_eco134106, w_eco134107, w_eco134108, w_eco134109, w_eco134110, w_eco134111, w_eco134112, w_eco134113, w_eco134114, w_eco134115, w_eco134116, w_eco134117, w_eco134118, w_eco134119, w_eco134120, w_eco134121, w_eco134122, w_eco134123, w_eco134124, w_eco134125, w_eco134126, w_eco134127, w_eco134128, w_eco134129, w_eco134130, w_eco134131, w_eco134132, w_eco134133, w_eco134134, w_eco134135, w_eco134136, w_eco134137, w_eco134138, w_eco134139, w_eco134140, w_eco134141, w_eco134142, w_eco134143, w_eco134144, w_eco134145, w_eco134146, w_eco134147, w_eco134148, w_eco134149, w_eco134150, w_eco134151, w_eco134152, w_eco134153, w_eco134154, w_eco134155, w_eco134156, w_eco134157, w_eco134158, w_eco134159, w_eco134160, w_eco134161, w_eco134162, w_eco134163, w_eco134164, w_eco134165, w_eco134166, w_eco134167, w_eco134168, w_eco134169, w_eco134170, w_eco134171, w_eco134172, w_eco134173, w_eco134174, w_eco134175, w_eco134176, w_eco134177, w_eco134178, w_eco134179, w_eco134180, w_eco134181, w_eco134182, w_eco134183, w_eco134184, w_eco134185, w_eco134186, w_eco134187, w_eco134188, w_eco134189, w_eco134190, w_eco134191, w_eco134192, w_eco134193, w_eco134194, w_eco134195, w_eco134196, w_eco134197, w_eco134198, w_eco134199, w_eco134200, w_eco134201, w_eco134202, w_eco134203, w_eco134204, w_eco134205, w_eco134206, w_eco134207, w_eco134208, w_eco134209, w_eco134210, w_eco134211, w_eco134212, w_eco134213, w_eco134214, w_eco134215, w_eco134216, w_eco134217, w_eco134218, w_eco134219, w_eco134220, w_eco134221, w_eco134222, w_eco134223, w_eco134224, w_eco134225, w_eco134226, w_eco134227, w_eco134228, w_eco134229, w_eco134230, w_eco134231, w_eco134232, w_eco134233, w_eco134234, w_eco134235, w_eco134236, w_eco134237, w_eco134238, w_eco134239, w_eco134240, w_eco134241, w_eco134242, w_eco134243, w_eco134244, w_eco134245, w_eco134246, w_eco134247, w_eco134248, w_eco134249, w_eco134250, w_eco134251, w_eco134252, w_eco134253, w_eco134254, w_eco134255, w_eco134256, w_eco134257, w_eco134258, w_eco134259, w_eco134260, w_eco134261, w_eco134262, w_eco134263, w_eco134264, w_eco134265, w_eco134266, w_eco134267, w_eco134268, w_eco134269, w_eco134270, w_eco134271, w_eco134272, w_eco134273, w_eco134274, w_eco134275, w_eco134276, w_eco134277, w_eco134278, w_eco134279, w_eco134280, w_eco134281, w_eco134282, w_eco134283, w_eco134284, w_eco134285, w_eco134286, w_eco134287, w_eco134288, w_eco134289, w_eco134290, w_eco134291, w_eco134292, w_eco134293, w_eco134294, w_eco134295, w_eco134296, w_eco134297, w_eco134298, w_eco134299, w_eco134300, w_eco134301, w_eco134302, w_eco134303, w_eco134304, w_eco134305, w_eco134306, w_eco134307, w_eco134308, w_eco134309, w_eco134310, w_eco134311, w_eco134312, w_eco134313, w_eco134314, w_eco134315, w_eco134316, w_eco134317, w_eco134318, w_eco134319, w_eco134320, w_eco134321, w_eco134322, w_eco134323, w_eco134324, w_eco134325, w_eco134326, w_eco134327, w_eco134328, w_eco134329, w_eco134330, w_eco134331, w_eco134332, w_eco134333, w_eco134334, w_eco134335, w_eco134336, w_eco134337, w_eco134338, w_eco134339, w_eco134340, w_eco134341, w_eco134342, w_eco134343, w_eco134344, w_eco134345, w_eco134346, w_eco134347, w_eco134348, w_eco134349, w_eco134350, w_eco134351, w_eco134352, w_eco134353, w_eco134354, w_eco134355, w_eco134356, w_eco134357, w_eco134358, w_eco134359, w_eco134360, w_eco134361, w_eco134362, w_eco134363, w_eco134364, w_eco134365, w_eco134366, w_eco134367, w_eco134368, w_eco134369, w_eco134370, w_eco134371, w_eco134372, w_eco134373, w_eco134374, w_eco134375, w_eco134376, w_eco134377, w_eco134378, w_eco134379, w_eco134380, w_eco134381, w_eco134382, w_eco134383, w_eco134384, w_eco134385, w_eco134386, w_eco134387, w_eco134388, w_eco134389, w_eco134390, w_eco134391, w_eco134392, w_eco134393, w_eco134394, w_eco134395, w_eco134396, w_eco134397, w_eco134398, w_eco134399, w_eco134400, w_eco134401, w_eco134402, w_eco134403, w_eco134404, w_eco134405, w_eco134406, w_eco134407, w_eco134408, w_eco134409, w_eco134410, w_eco134411, w_eco134412, w_eco134413, w_eco134414, w_eco134415, w_eco134416, w_eco134417, w_eco134418, w_eco134419, w_eco134420, w_eco134421, w_eco134422, w_eco134423, w_eco134424, w_eco134425, w_eco134426, w_eco134427, w_eco134428, w_eco134429, w_eco134430, w_eco134431, w_eco134432, w_eco134433, w_eco134434, w_eco134435, w_eco134436, w_eco134437, w_eco134438, w_eco134439, w_eco134440, w_eco134441, w_eco134442, w_eco134443, w_eco134444, w_eco134445, w_eco134446, w_eco134447, w_eco134448, w_eco134449, w_eco134450, w_eco134451, w_eco134452, w_eco134453, w_eco134454, w_eco134455, w_eco134456, w_eco134457, w_eco134458, w_eco134459, w_eco134460, w_eco134461, w_eco134462, w_eco134463, w_eco134464, w_eco134465, w_eco134466, w_eco134467, w_eco134468, w_eco134469, w_eco134470, w_eco134471, w_eco134472, w_eco134473, w_eco134474, w_eco134475, w_eco134476, w_eco134477, w_eco134478, w_eco134479, w_eco134480, w_eco134481, w_eco134482, w_eco134483, w_eco134484, w_eco134485, w_eco134486, w_eco134487, w_eco134488, w_eco134489, w_eco134490, w_eco134491, w_eco134492, w_eco134493, w_eco134494, w_eco134495, w_eco134496, w_eco134497, w_eco134498, w_eco134499, w_eco134500, w_eco134501, w_eco134502, w_eco134503, w_eco134504, w_eco134505, w_eco134506, w_eco134507, w_eco134508, w_eco134509, w_eco134510, w_eco134511, w_eco134512, w_eco134513, w_eco134514, w_eco134515, w_eco134516, w_eco134517, w_eco134518, w_eco134519, w_eco134520, w_eco134521, w_eco134522, w_eco134523, w_eco134524, w_eco134525, w_eco134526, w_eco134527, w_eco134528, w_eco134529, w_eco134530, w_eco134531, w_eco134532, w_eco134533, w_eco134534, w_eco134535, w_eco134536, w_eco134537, w_eco134538, w_eco134539, w_eco134540, w_eco134541, w_eco134542, w_eco134543, w_eco134544, w_eco134545, w_eco134546, w_eco134547, w_eco134548, w_eco134549, w_eco134550, w_eco134551, w_eco134552, w_eco134553, w_eco134554, w_eco134555, w_eco134556, w_eco134557, w_eco134558, w_eco134559, w_eco134560, w_eco134561, w_eco134562, w_eco134563, w_eco134564, w_eco134565, w_eco134566, w_eco134567, w_eco134568, w_eco134569, w_eco134570, w_eco134571, w_eco134572, w_eco134573, w_eco134574, w_eco134575, w_eco134576, w_eco134577, w_eco134578, w_eco134579, w_eco134580, w_eco134581, w_eco134582, w_eco134583, w_eco134584, w_eco134585, w_eco134586, w_eco134587, w_eco134588, w_eco134589, w_eco134590, w_eco134591, w_eco134592, w_eco134593, w_eco134594, w_eco134595, w_eco134596, w_eco134597, w_eco134598, w_eco134599, w_eco134600, w_eco134601, w_eco134602, w_eco134603, w_eco134604, w_eco134605, w_eco134606, w_eco134607, w_eco134608, w_eco134609, w_eco134610, w_eco134611, w_eco134612, w_eco134613, w_eco134614, w_eco134615, w_eco134616, w_eco134617, w_eco134618, w_eco134619, w_eco134620, w_eco134621, w_eco134622, w_eco134623, w_eco134624, w_eco134625, w_eco134626, w_eco134627, w_eco134628, w_eco134629, w_eco134630, w_eco134631, w_eco134632, w_eco134633, w_eco134634, w_eco134635, w_eco134636, w_eco134637, w_eco134638, w_eco134639, w_eco134640, w_eco134641, w_eco134642, w_eco134643, w_eco134644, w_eco134645, w_eco134646, w_eco134647, w_eco134648, w_eco134649, w_eco134650, w_eco134651, w_eco134652, w_eco134653, w_eco134654, w_eco134655, w_eco134656, w_eco134657, w_eco134658, w_eco134659, w_eco134660, w_eco134661, w_eco134662, w_eco134663, w_eco134664, w_eco134665, w_eco134666, w_eco134667, w_eco134668, w_eco134669, w_eco134670, w_eco134671, w_eco134672, w_eco134673, w_eco134674, w_eco134675, w_eco134676, w_eco134677, w_eco134678, w_eco134679, w_eco134680, w_eco134681, w_eco134682, w_eco134683, w_eco134684, w_eco134685, w_eco134686, w_eco134687, w_eco134688, w_eco134689, w_eco134690, w_eco134691, w_eco134692, w_eco134693, w_eco134694, w_eco134695, w_eco134696, w_eco134697, w_eco134698, w_eco134699, w_eco134700, w_eco134701, w_eco134702, w_eco134703, w_eco134704, w_eco134705, w_eco134706, w_eco134707, w_eco134708, w_eco134709, w_eco134710, w_eco134711, w_eco134712, w_eco134713, w_eco134714, w_eco134715, w_eco134716, w_eco134717, w_eco134718, w_eco134719, w_eco134720, w_eco134721, w_eco134722, w_eco134723, w_eco134724, w_eco134725, w_eco134726, w_eco134727, w_eco134728, w_eco134729, w_eco134730, w_eco134731, w_eco134732, w_eco134733, w_eco134734, w_eco134735, w_eco134736, w_eco134737, w_eco134738, w_eco134739, w_eco134740, w_eco134741, w_eco134742, w_eco134743, w_eco134744, w_eco134745, w_eco134746, w_eco134747, w_eco134748, w_eco134749, w_eco134750, w_eco134751, w_eco134752, w_eco134753, w_eco134754, w_eco134755, w_eco134756, w_eco134757, w_eco134758, w_eco134759, w_eco134760, w_eco134761, w_eco134762, w_eco134763, w_eco134764, w_eco134765, w_eco134766, w_eco134767, w_eco134768, w_eco134769, w_eco134770, w_eco134771, w_eco134772, w_eco134773, w_eco134774, w_eco134775, w_eco134776, w_eco134777, w_eco134778, w_eco134779, w_eco134780, w_eco134781, w_eco134782, w_eco134783, w_eco134784, w_eco134785, w_eco134786, w_eco134787, w_eco134788, w_eco134789, w_eco134790, w_eco134791, w_eco134792, w_eco134793, w_eco134794, w_eco134795, w_eco134796, w_eco134797, w_eco134798, w_eco134799, w_eco134800, w_eco134801, w_eco134802, w_eco134803, w_eco134804, w_eco134805, w_eco134806, w_eco134807, w_eco134808, w_eco134809, w_eco134810, w_eco134811, w_eco134812, w_eco134813, w_eco134814, w_eco134815, w_eco134816, w_eco134817, w_eco134818, w_eco134819, w_eco134820, w_eco134821, w_eco134822, w_eco134823, w_eco134824, w_eco134825, w_eco134826, w_eco134827, w_eco134828, w_eco134829, w_eco134830, w_eco134831, w_eco134832, w_eco134833, w_eco134834, w_eco134835, w_eco134836, w_eco134837, w_eco134838, w_eco134839, w_eco134840, w_eco134841, w_eco134842, w_eco134843, w_eco134844, w_eco134845, w_eco134846, w_eco134847, w_eco134848, w_eco134849, w_eco134850, w_eco134851, w_eco134852, w_eco134853, w_eco134854, w_eco134855, w_eco134856, w_eco134857, w_eco134858, w_eco134859, w_eco134860, w_eco134861, w_eco134862, w_eco134863, w_eco134864, w_eco134865, w_eco134866, w_eco134867, w_eco134868, w_eco134869, w_eco134870, w_eco134871, w_eco134872, w_eco134873, w_eco134874, w_eco134875, w_eco134876, w_eco134877, w_eco134878, w_eco134879, w_eco134880, w_eco134881, w_eco134882, w_eco134883, w_eco134884, w_eco134885, w_eco134886, w_eco134887, w_eco134888, w_eco134889, w_eco134890, w_eco134891, w_eco134892, w_eco134893, w_eco134894, w_eco134895, w_eco134896, w_eco134897, w_eco134898, w_eco134899, w_eco134900, w_eco134901, w_eco134902, w_eco134903, w_eco134904, w_eco134905, w_eco134906, w_eco134907, w_eco134908, w_eco134909, w_eco134910, w_eco134911, w_eco134912, w_eco134913, w_eco134914, w_eco134915, w_eco134916, w_eco134917, w_eco134918, w_eco134919, w_eco134920, w_eco134921, w_eco134922, w_eco134923, w_eco134924, w_eco134925, w_eco134926, w_eco134927, w_eco134928, w_eco134929, w_eco134930, w_eco134931, w_eco134932, w_eco134933, w_eco134934, w_eco134935, w_eco134936, w_eco134937, w_eco134938, w_eco134939, w_eco134940, w_eco134941, w_eco134942, w_eco134943, w_eco134944, w_eco134945, w_eco134946, w_eco134947, w_eco134948, w_eco134949, w_eco134950, w_eco134951, w_eco134952, w_eco134953, w_eco134954, w_eco134955, w_eco134956, w_eco134957, w_eco134958, w_eco134959, w_eco134960, w_eco134961, w_eco134962, w_eco134963, w_eco134964, w_eco134965, w_eco134966, w_eco134967, w_eco134968, w_eco134969, w_eco134970, w_eco134971, w_eco134972, w_eco134973, w_eco134974, w_eco134975, w_eco134976, w_eco134977, w_eco134978, w_eco134979, w_eco134980, w_eco134981, w_eco134982, w_eco134983, w_eco134984, w_eco134985, w_eco134986, w_eco134987, w_eco134988, w_eco134989, w_eco134990, w_eco134991, w_eco134992, w_eco134993, w_eco134994, w_eco134995, w_eco134996, w_eco134997, w_eco134998, w_eco134999, w_eco135000, w_eco135001, w_eco135002, w_eco135003, w_eco135004, w_eco135005, w_eco135006, w_eco135007, w_eco135008, w_eco135009, w_eco135010, w_eco135011, w_eco135012, w_eco135013, w_eco135014, w_eco135015, w_eco135016, w_eco135017, w_eco135018, w_eco135019, w_eco135020, w_eco135021, w_eco135022, w_eco135023, w_eco135024, w_eco135025, w_eco135026, w_eco135027, w_eco135028, w_eco135029, w_eco135030, w_eco135031, w_eco135032, w_eco135033, w_eco135034, w_eco135035, w_eco135036, w_eco135037, w_eco135038, w_eco135039, w_eco135040, w_eco135041, w_eco135042, w_eco135043, w_eco135044, w_eco135045, w_eco135046, w_eco135047, w_eco135048, w_eco135049, w_eco135050, w_eco135051, w_eco135052, w_eco135053, w_eco135054, w_eco135055, w_eco135056, w_eco135057, w_eco135058, w_eco135059, w_eco135060, w_eco135061, w_eco135062, w_eco135063, w_eco135064, w_eco135065, w_eco135066, w_eco135067, w_eco135068, w_eco135069, w_eco135070, w_eco135071, w_eco135072, w_eco135073, w_eco135074, w_eco135075, w_eco135076, w_eco135077, w_eco135078, w_eco135079, w_eco135080, w_eco135081, w_eco135082, w_eco135083, w_eco135084, w_eco135085, w_eco135086, w_eco135087, w_eco135088, w_eco135089, w_eco135090, w_eco135091, w_eco135092, w_eco135093, w_eco135094, w_eco135095, w_eco135096, w_eco135097, w_eco135098, w_eco135099, w_eco135100, w_eco135101, w_eco135102, w_eco135103, w_eco135104, w_eco135105, w_eco135106, w_eco135107, w_eco135108, w_eco135109, w_eco135110, w_eco135111, w_eco135112, w_eco135113, w_eco135114, w_eco135115, w_eco135116, w_eco135117, w_eco135118, w_eco135119, w_eco135120, w_eco135121, w_eco135122, w_eco135123, w_eco135124, w_eco135125, w_eco135126, w_eco135127, w_eco135128, w_eco135129, w_eco135130, w_eco135131, w_eco135132, w_eco135133, w_eco135134, w_eco135135, w_eco135136, w_eco135137, w_eco135138, w_eco135139, w_eco135140, w_eco135141, w_eco135142, w_eco135143, w_eco135144, w_eco135145, w_eco135146, w_eco135147, w_eco135148, w_eco135149, w_eco135150, w_eco135151, w_eco135152, w_eco135153, w_eco135154, w_eco135155, w_eco135156, w_eco135157, w_eco135158, w_eco135159, w_eco135160, w_eco135161, w_eco135162, w_eco135163, w_eco135164, w_eco135165, w_eco135166, w_eco135167, w_eco135168, w_eco135169, w_eco135170, w_eco135171, w_eco135172, w_eco135173, w_eco135174, w_eco135175, w_eco135176, w_eco135177, w_eco135178, w_eco135179, w_eco135180, w_eco135181, w_eco135182, w_eco135183, w_eco135184, w_eco135185, w_eco135186, w_eco135187, w_eco135188, w_eco135189, w_eco135190, w_eco135191, w_eco135192, w_eco135193, w_eco135194, w_eco135195, w_eco135196, w_eco135197, w_eco135198, w_eco135199, w_eco135200, w_eco135201, w_eco135202, w_eco135203, w_eco135204, w_eco135205, w_eco135206, w_eco135207, w_eco135208, w_eco135209, w_eco135210, w_eco135211, w_eco135212, w_eco135213, w_eco135214, w_eco135215, w_eco135216, w_eco135217, w_eco135218, w_eco135219, w_eco135220, w_eco135221, w_eco135222, w_eco135223, w_eco135224, w_eco135225, w_eco135226, w_eco135227, w_eco135228, w_eco135229, w_eco135230, w_eco135231, w_eco135232, w_eco135233, w_eco135234, w_eco135235, w_eco135236, w_eco135237, w_eco135238, w_eco135239, w_eco135240, w_eco135241, w_eco135242, w_eco135243, w_eco135244, w_eco135245, w_eco135246, w_eco135247, w_eco135248, w_eco135249, w_eco135250, w_eco135251, w_eco135252, w_eco135253, w_eco135254, w_eco135255, w_eco135256, w_eco135257, w_eco135258, w_eco135259, w_eco135260, w_eco135261, w_eco135262, w_eco135263, w_eco135264, w_eco135265, w_eco135266, w_eco135267, w_eco135268, w_eco135269, w_eco135270, w_eco135271, w_eco135272, w_eco135273, w_eco135274, w_eco135275, w_eco135276, w_eco135277, w_eco135278, w_eco135279, w_eco135280, w_eco135281, w_eco135282, w_eco135283, w_eco135284, w_eco135285, w_eco135286, w_eco135287, w_eco135288, w_eco135289, w_eco135290, w_eco135291, w_eco135292, w_eco135293, w_eco135294, w_eco135295, w_eco135296, w_eco135297, w_eco135298, w_eco135299, w_eco135300, w_eco135301, w_eco135302, w_eco135303, w_eco135304, w_eco135305, w_eco135306, w_eco135307, w_eco135308, w_eco135309, w_eco135310, w_eco135311, w_eco135312, w_eco135313, w_eco135314, w_eco135315, w_eco135316, w_eco135317, w_eco135318, w_eco135319, w_eco135320, w_eco135321, w_eco135322, w_eco135323, w_eco135324, w_eco135325, w_eco135326, w_eco135327, w_eco135328, w_eco135329, w_eco135330, w_eco135331, w_eco135332, w_eco135333, w_eco135334, w_eco135335, w_eco135336, w_eco135337, w_eco135338, w_eco135339, w_eco135340, w_eco135341, w_eco135342, w_eco135343, w_eco135344, w_eco135345, w_eco135346, w_eco135347, w_eco135348, w_eco135349, w_eco135350, w_eco135351, w_eco135352, w_eco135353, w_eco135354, w_eco135355, w_eco135356, w_eco135357, w_eco135358, w_eco135359, w_eco135360, w_eco135361, w_eco135362, w_eco135363, w_eco135364, w_eco135365, w_eco135366, w_eco135367, w_eco135368, w_eco135369, w_eco135370, w_eco135371, w_eco135372, w_eco135373, w_eco135374, w_eco135375, w_eco135376, w_eco135377, w_eco135378, w_eco135379, w_eco135380, w_eco135381, w_eco135382, w_eco135383, w_eco135384, w_eco135385, w_eco135386, w_eco135387, w_eco135388, w_eco135389, w_eco135390, w_eco135391, w_eco135392, w_eco135393, w_eco135394, w_eco135395, w_eco135396, w_eco135397, w_eco135398, w_eco135399, w_eco135400, w_eco135401, w_eco135402, w_eco135403, w_eco135404, w_eco135405, w_eco135406, w_eco135407, w_eco135408, w_eco135409, w_eco135410, w_eco135411, w_eco135412, w_eco135413, w_eco135414, w_eco135415, w_eco135416, w_eco135417, w_eco135418, w_eco135419, w_eco135420, w_eco135421, w_eco135422, w_eco135423, w_eco135424, w_eco135425, w_eco135426, w_eco135427, w_eco135428, w_eco135429, w_eco135430, w_eco135431, w_eco135432, w_eco135433, w_eco135434, w_eco135435, w_eco135436, w_eco135437, w_eco135438, w_eco135439, w_eco135440, w_eco135441, w_eco135442, w_eco135443, w_eco135444, w_eco135445, w_eco135446, w_eco135447, w_eco135448, w_eco135449, w_eco135450, w_eco135451, w_eco135452, w_eco135453, w_eco135454, w_eco135455, w_eco135456, w_eco135457, w_eco135458, w_eco135459, w_eco135460, w_eco135461, w_eco135462, w_eco135463, w_eco135464, w_eco135465, w_eco135466, w_eco135467, w_eco135468, w_eco135469, w_eco135470, w_eco135471, w_eco135472, w_eco135473, w_eco135474, w_eco135475, w_eco135476, w_eco135477, w_eco135478, w_eco135479, w_eco135480, w_eco135481, w_eco135482, w_eco135483, w_eco135484, w_eco135485, w_eco135486, w_eco135487, w_eco135488, w_eco135489, w_eco135490, w_eco135491, w_eco135492, w_eco135493, w_eco135494, w_eco135495, w_eco135496, w_eco135497, w_eco135498, w_eco135499, w_eco135500, w_eco135501, w_eco135502, w_eco135503, w_eco135504, w_eco135505, w_eco135506, w_eco135507, w_eco135508, w_eco135509, w_eco135510, w_eco135511, w_eco135512, w_eco135513, w_eco135514, w_eco135515, w_eco135516, w_eco135517, w_eco135518, w_eco135519, w_eco135520, w_eco135521, w_eco135522, w_eco135523, w_eco135524, w_eco135525, w_eco135526, w_eco135527, w_eco135528, w_eco135529, w_eco135530, w_eco135531, w_eco135532, w_eco135533, w_eco135534, w_eco135535, w_eco135536, w_eco135537, w_eco135538, w_eco135539, w_eco135540, w_eco135541, w_eco135542, w_eco135543, w_eco135544, w_eco135545, w_eco135546, w_eco135547, w_eco135548, w_eco135549, w_eco135550, w_eco135551, w_eco135552, w_eco135553, w_eco135554, w_eco135555, w_eco135556, w_eco135557, w_eco135558, w_eco135559, w_eco135560, w_eco135561, w_eco135562, w_eco135563, w_eco135564, w_eco135565, w_eco135566, w_eco135567, w_eco135568, w_eco135569, w_eco135570, w_eco135571, w_eco135572, w_eco135573, w_eco135574, w_eco135575, w_eco135576, w_eco135577, w_eco135578, w_eco135579, w_eco135580, w_eco135581, w_eco135582, w_eco135583, w_eco135584, w_eco135585, w_eco135586, w_eco135587, w_eco135588, w_eco135589, w_eco135590, w_eco135591, w_eco135592, w_eco135593, w_eco135594, w_eco135595, w_eco135596, w_eco135597, w_eco135598, w_eco135599, w_eco135600, w_eco135601, w_eco135602, w_eco135603, w_eco135604, w_eco135605, w_eco135606, w_eco135607, w_eco135608, w_eco135609, w_eco135610, w_eco135611, w_eco135612, w_eco135613, w_eco135614, w_eco135615, w_eco135616, w_eco135617, w_eco135618, w_eco135619, w_eco135620, w_eco135621, w_eco135622, w_eco135623, w_eco135624, w_eco135625, w_eco135626, w_eco135627, w_eco135628, w_eco135629, w_eco135630, w_eco135631, w_eco135632, w_eco135633, w_eco135634, w_eco135635, w_eco135636, w_eco135637, w_eco135638, w_eco135639, w_eco135640, w_eco135641, w_eco135642, w_eco135643, w_eco135644, w_eco135645, w_eco135646, w_eco135647, w_eco135648, w_eco135649, w_eco135650, w_eco135651, w_eco135652, w_eco135653, w_eco135654, w_eco135655, w_eco135656, w_eco135657, w_eco135658, w_eco135659, w_eco135660, w_eco135661, w_eco135662, w_eco135663, w_eco135664, w_eco135665, w_eco135666, w_eco135667, w_eco135668, w_eco135669, w_eco135670, w_eco135671, w_eco135672, w_eco135673, w_eco135674, w_eco135675, w_eco135676, w_eco135677, w_eco135678, w_eco135679, w_eco135680, w_eco135681, w_eco135682, w_eco135683, w_eco135684, w_eco135685, w_eco135686, w_eco135687, w_eco135688, w_eco135689, w_eco135690, w_eco135691, w_eco135692, w_eco135693, w_eco135694, w_eco135695, w_eco135696, w_eco135697, w_eco135698, w_eco135699, w_eco135700, w_eco135701, w_eco135702, w_eco135703, w_eco135704, w_eco135705, w_eco135706, w_eco135707, w_eco135708, w_eco135709, w_eco135710, w_eco135711, w_eco135712, w_eco135713, w_eco135714, w_eco135715, w_eco135716, w_eco135717, w_eco135718, w_eco135719, w_eco135720, w_eco135721, w_eco135722, w_eco135723, w_eco135724, w_eco135725, w_eco135726, w_eco135727, w_eco135728, w_eco135729, w_eco135730, w_eco135731, w_eco135732, w_eco135733, w_eco135734, w_eco135735, w_eco135736, w_eco135737, w_eco135738, w_eco135739, w_eco135740, w_eco135741, w_eco135742, w_eco135743, w_eco135744, w_eco135745, w_eco135746, w_eco135747, w_eco135748, w_eco135749, w_eco135750, w_eco135751, w_eco135752, w_eco135753, w_eco135754, w_eco135755, w_eco135756, w_eco135757, w_eco135758, w_eco135759, w_eco135760, w_eco135761, w_eco135762, w_eco135763, w_eco135764, w_eco135765, w_eco135766, w_eco135767, w_eco135768, w_eco135769, w_eco135770, w_eco135771, w_eco135772, w_eco135773, w_eco135774, w_eco135775, w_eco135776, w_eco135777, w_eco135778, w_eco135779, w_eco135780, w_eco135781, w_eco135782, w_eco135783, w_eco135784, w_eco135785, w_eco135786, w_eco135787, w_eco135788, w_eco135789, w_eco135790, w_eco135791, w_eco135792, w_eco135793, w_eco135794, w_eco135795, w_eco135796, w_eco135797, w_eco135798, w_eco135799, w_eco135800, w_eco135801, w_eco135802, w_eco135803, w_eco135804, w_eco135805, w_eco135806, w_eco135807, w_eco135808, w_eco135809, w_eco135810, w_eco135811, w_eco135812, w_eco135813, w_eco135814, w_eco135815, w_eco135816, w_eco135817, w_eco135818, w_eco135819, w_eco135820, w_eco135821, w_eco135822, w_eco135823, w_eco135824, w_eco135825, w_eco135826, w_eco135827, w_eco135828, w_eco135829, w_eco135830, w_eco135831, w_eco135832, w_eco135833, w_eco135834, w_eco135835, w_eco135836, w_eco135837, w_eco135838, w_eco135839, w_eco135840, w_eco135841, w_eco135842, w_eco135843, w_eco135844, w_eco135845, w_eco135846, w_eco135847, w_eco135848, w_eco135849, w_eco135850, w_eco135851, w_eco135852, w_eco135853, w_eco135854, w_eco135855, w_eco135856, w_eco135857, w_eco135858, w_eco135859, w_eco135860, w_eco135861, w_eco135862, w_eco135863, w_eco135864, w_eco135865, w_eco135866, w_eco135867, w_eco135868, w_eco135869, w_eco135870, w_eco135871, w_eco135872, w_eco135873, w_eco135874, w_eco135875, w_eco135876, w_eco135877, w_eco135878, w_eco135879, w_eco135880, w_eco135881, w_eco135882, w_eco135883, w_eco135884, w_eco135885, w_eco135886, w_eco135887, w_eco135888, w_eco135889, w_eco135890, w_eco135891, w_eco135892, w_eco135893, w_eco135894, w_eco135895, w_eco135896, w_eco135897, w_eco135898, w_eco135899, w_eco135900, w_eco135901, w_eco135902, w_eco135903, w_eco135904, w_eco135905, w_eco135906, w_eco135907, w_eco135908, w_eco135909, w_eco135910, w_eco135911, w_eco135912, w_eco135913, w_eco135914, w_eco135915, w_eco135916, w_eco135917, w_eco135918, w_eco135919, w_eco135920, w_eco135921, w_eco135922, w_eco135923, w_eco135924, w_eco135925, w_eco135926, w_eco135927, w_eco135928, w_eco135929, w_eco135930, w_eco135931, w_eco135932, w_eco135933, w_eco135934, w_eco135935, w_eco135936, w_eco135937, w_eco135938, w_eco135939, w_eco135940, w_eco135941, w_eco135942, w_eco135943, w_eco135944, w_eco135945, w_eco135946, w_eco135947, w_eco135948, w_eco135949, w_eco135950, w_eco135951, w_eco135952, w_eco135953, w_eco135954, w_eco135955, w_eco135956, w_eco135957, w_eco135958, w_eco135959, w_eco135960, w_eco135961, w_eco135962, w_eco135963, w_eco135964, w_eco135965, w_eco135966, w_eco135967, w_eco135968, w_eco135969, w_eco135970, w_eco135971, w_eco135972, w_eco135973, w_eco135974, w_eco135975, w_eco135976, w_eco135977, w_eco135978, w_eco135979, w_eco135980, w_eco135981, w_eco135982, w_eco135983, w_eco135984, w_eco135985, w_eco135986, w_eco135987, w_eco135988, w_eco135989, w_eco135990, w_eco135991, w_eco135992, w_eco135993, w_eco135994, w_eco135995, w_eco135996, w_eco135997, w_eco135998, w_eco135999, w_eco136000, w_eco136001, w_eco136002, w_eco136003, w_eco136004, w_eco136005, w_eco136006, w_eco136007, w_eco136008, w_eco136009, w_eco136010, w_eco136011, w_eco136012, w_eco136013, w_eco136014, w_eco136015, w_eco136016, w_eco136017, w_eco136018, w_eco136019, w_eco136020, w_eco136021, w_eco136022, w_eco136023, w_eco136024, w_eco136025, w_eco136026, w_eco136027, w_eco136028, w_eco136029, w_eco136030, w_eco136031, w_eco136032, w_eco136033, w_eco136034, w_eco136035, w_eco136036, w_eco136037, w_eco136038, w_eco136039, w_eco136040, w_eco136041, w_eco136042, w_eco136043, w_eco136044, w_eco136045, w_eco136046, w_eco136047, w_eco136048, w_eco136049, w_eco136050, w_eco136051, w_eco136052, w_eco136053, w_eco136054, w_eco136055, w_eco136056, w_eco136057, w_eco136058, w_eco136059, w_eco136060, w_eco136061, w_eco136062, w_eco136063, w_eco136064, w_eco136065, w_eco136066, w_eco136067, w_eco136068, w_eco136069, w_eco136070, w_eco136071, w_eco136072, w_eco136073, w_eco136074, w_eco136075, w_eco136076, w_eco136077, w_eco136078, w_eco136079, w_eco136080, w_eco136081, w_eco136082, w_eco136083, w_eco136084, w_eco136085, w_eco136086, w_eco136087, w_eco136088, w_eco136089, w_eco136090, w_eco136091, w_eco136092, w_eco136093, w_eco136094, w_eco136095, w_eco136096, w_eco136097, w_eco136098, w_eco136099, w_eco136100, w_eco136101, w_eco136102, w_eco136103, w_eco136104, w_eco136105, w_eco136106, w_eco136107, w_eco136108, w_eco136109, w_eco136110, w_eco136111, w_eco136112, w_eco136113, w_eco136114, w_eco136115, w_eco136116, w_eco136117, w_eco136118, w_eco136119, w_eco136120, w_eco136121, w_eco136122, w_eco136123, w_eco136124, w_eco136125, w_eco136126, w_eco136127, w_eco136128, w_eco136129, w_eco136130, w_eco136131, w_eco136132, w_eco136133, w_eco136134, w_eco136135, w_eco136136, w_eco136137, w_eco136138, w_eco136139, w_eco136140, w_eco136141, w_eco136142, w_eco136143, w_eco136144, w_eco136145, w_eco136146, w_eco136147, w_eco136148, w_eco136149, w_eco136150, w_eco136151, w_eco136152, w_eco136153, w_eco136154, w_eco136155, w_eco136156, w_eco136157, w_eco136158, w_eco136159, w_eco136160, w_eco136161, w_eco136162, w_eco136163, w_eco136164, w_eco136165, w_eco136166, w_eco136167, w_eco136168, w_eco136169, w_eco136170, w_eco136171, w_eco136172, w_eco136173, w_eco136174, w_eco136175, w_eco136176, w_eco136177, w_eco136178, w_eco136179, w_eco136180, w_eco136181, w_eco136182, w_eco136183, w_eco136184, w_eco136185, w_eco136186, w_eco136187, w_eco136188, w_eco136189, w_eco136190, w_eco136191, w_eco136192, w_eco136193, w_eco136194, w_eco136195, w_eco136196, w_eco136197, w_eco136198, w_eco136199, w_eco136200, w_eco136201, w_eco136202, w_eco136203, w_eco136204, w_eco136205, w_eco136206, w_eco136207, w_eco136208, w_eco136209, w_eco136210, w_eco136211, w_eco136212, w_eco136213, w_eco136214, w_eco136215, w_eco136216, w_eco136217, w_eco136218, w_eco136219, w_eco136220, w_eco136221, w_eco136222, w_eco136223, w_eco136224, w_eco136225, w_eco136226, w_eco136227, w_eco136228, w_eco136229, w_eco136230, w_eco136231, w_eco136232, w_eco136233, w_eco136234, w_eco136235, w_eco136236, w_eco136237, w_eco136238, w_eco136239, w_eco136240, w_eco136241, w_eco136242, w_eco136243, w_eco136244, w_eco136245, w_eco136246, w_eco136247, w_eco136248, w_eco136249, w_eco136250, w_eco136251, w_eco136252, w_eco136253, w_eco136254, w_eco136255, w_eco136256, w_eco136257, w_eco136258, w_eco136259, w_eco136260, w_eco136261, w_eco136262, w_eco136263, w_eco136264, w_eco136265, w_eco136266, w_eco136267, w_eco136268, w_eco136269, w_eco136270, w_eco136271, w_eco136272, w_eco136273, w_eco136274, w_eco136275, w_eco136276, w_eco136277, w_eco136278, w_eco136279, w_eco136280, w_eco136281, w_eco136282, w_eco136283, w_eco136284, w_eco136285, w_eco136286, w_eco136287, w_eco136288, w_eco136289, w_eco136290, w_eco136291, w_eco136292, w_eco136293, w_eco136294, w_eco136295, w_eco136296, w_eco136297, w_eco136298, w_eco136299, w_eco136300, w_eco136301, w_eco136302, w_eco136303, w_eco136304, w_eco136305, w_eco136306, w_eco136307, w_eco136308, w_eco136309, w_eco136310, w_eco136311, w_eco136312, w_eco136313, w_eco136314, w_eco136315, w_eco136316, w_eco136317, w_eco136318, w_eco136319, w_eco136320, w_eco136321, w_eco136322, w_eco136323, w_eco136324, w_eco136325, w_eco136326, w_eco136327, w_eco136328, w_eco136329, w_eco136330, w_eco136331, w_eco136332, w_eco136333, w_eco136334, w_eco136335, w_eco136336, w_eco136337, w_eco136338, w_eco136339, w_eco136340, w_eco136341, w_eco136342, w_eco136343, w_eco136344, w_eco136345, w_eco136346, w_eco136347, w_eco136348, w_eco136349, w_eco136350, w_eco136351, w_eco136352, w_eco136353, w_eco136354, w_eco136355, w_eco136356, w_eco136357, w_eco136358, w_eco136359, w_eco136360, w_eco136361, w_eco136362, w_eco136363, w_eco136364, w_eco136365, w_eco136366, w_eco136367, w_eco136368, w_eco136369, w_eco136370, w_eco136371, w_eco136372, w_eco136373, w_eco136374, w_eco136375, w_eco136376, w_eco136377, w_eco136378, w_eco136379, w_eco136380, w_eco136381, w_eco136382, w_eco136383, w_eco136384, w_eco136385, w_eco136386, w_eco136387, w_eco136388, w_eco136389, w_eco136390, w_eco136391, w_eco136392, w_eco136393, w_eco136394, w_eco136395, w_eco136396, w_eco136397, w_eco136398, w_eco136399, w_eco136400, w_eco136401, w_eco136402, w_eco136403, w_eco136404, w_eco136405, w_eco136406, w_eco136407, w_eco136408, w_eco136409, w_eco136410, w_eco136411, w_eco136412, w_eco136413, w_eco136414, w_eco136415, w_eco136416, w_eco136417, w_eco136418, w_eco136419, w_eco136420, w_eco136421, w_eco136422, w_eco136423, w_eco136424, w_eco136425, w_eco136426, w_eco136427, w_eco136428, w_eco136429, w_eco136430, w_eco136431, w_eco136432, w_eco136433, w_eco136434, w_eco136435, w_eco136436, w_eco136437, w_eco136438, w_eco136439, w_eco136440, w_eco136441, w_eco136442, w_eco136443, w_eco136444, w_eco136445, w_eco136446, w_eco136447, w_eco136448, w_eco136449, w_eco136450, w_eco136451, w_eco136452, w_eco136453, w_eco136454, w_eco136455, w_eco136456, w_eco136457, w_eco136458, w_eco136459, w_eco136460, w_eco136461, w_eco136462, w_eco136463, w_eco136464, w_eco136465, w_eco136466, w_eco136467, w_eco136468, w_eco136469, w_eco136470, w_eco136471, w_eco136472, w_eco136473, w_eco136474, w_eco136475, w_eco136476, w_eco136477, w_eco136478, w_eco136479, w_eco136480, w_eco136481, w_eco136482, w_eco136483, w_eco136484, w_eco136485, w_eco136486, w_eco136487, w_eco136488, w_eco136489, w_eco136490, w_eco136491, w_eco136492, w_eco136493, w_eco136494, w_eco136495, w_eco136496, w_eco136497, w_eco136498, w_eco136499, w_eco136500, w_eco136501, w_eco136502, w_eco136503, w_eco136504, w_eco136505, w_eco136506, w_eco136507, w_eco136508, w_eco136509, w_eco136510, w_eco136511, w_eco136512, w_eco136513, w_eco136514, w_eco136515, w_eco136516, w_eco136517, w_eco136518, w_eco136519, w_eco136520, w_eco136521, w_eco136522, w_eco136523, w_eco136524, w_eco136525, w_eco136526, w_eco136527, w_eco136528, w_eco136529, w_eco136530, w_eco136531, w_eco136532, w_eco136533, w_eco136534, w_eco136535, w_eco136536, w_eco136537, w_eco136538, w_eco136539, w_eco136540, w_eco136541, w_eco136542, w_eco136543, w_eco136544, w_eco136545, w_eco136546, w_eco136547, w_eco136548, w_eco136549, w_eco136550, w_eco136551, w_eco136552, w_eco136553, w_eco136554, w_eco136555, w_eco136556, w_eco136557, w_eco136558, w_eco136559, w_eco136560, w_eco136561, w_eco136562, w_eco136563, w_eco136564, w_eco136565, w_eco136566, w_eco136567, w_eco136568, w_eco136569, w_eco136570, w_eco136571, w_eco136572, w_eco136573, w_eco136574, w_eco136575, w_eco136576, w_eco136577, w_eco136578, w_eco136579, w_eco136580, w_eco136581, w_eco136582, w_eco136583, w_eco136584, w_eco136585, w_eco136586, w_eco136587, w_eco136588, w_eco136589, w_eco136590, w_eco136591, w_eco136592, w_eco136593, w_eco136594, w_eco136595, w_eco136596, w_eco136597, w_eco136598, w_eco136599, w_eco136600, w_eco136601, w_eco136602, w_eco136603, w_eco136604, w_eco136605, w_eco136606, w_eco136607, w_eco136608, w_eco136609, w_eco136610, w_eco136611, w_eco136612, w_eco136613, w_eco136614, w_eco136615, w_eco136616, w_eco136617, w_eco136618, w_eco136619, w_eco136620, w_eco136621, w_eco136622, w_eco136623, w_eco136624, w_eco136625, w_eco136626, w_eco136627, w_eco136628, w_eco136629, w_eco136630, w_eco136631, w_eco136632, w_eco136633, w_eco136634, w_eco136635, w_eco136636, w_eco136637, w_eco136638, w_eco136639, w_eco136640, w_eco136641, w_eco136642, w_eco136643, w_eco136644, w_eco136645, w_eco136646, w_eco136647, w_eco136648, w_eco136649, w_eco136650, w_eco136651, w_eco136652, w_eco136653, w_eco136654, w_eco136655, w_eco136656, w_eco136657, w_eco136658, w_eco136659, w_eco136660, w_eco136661, w_eco136662, w_eco136663, w_eco136664, w_eco136665, w_eco136666, w_eco136667, w_eco136668, w_eco136669, w_eco136670, w_eco136671, w_eco136672, w_eco136673, w_eco136674, w_eco136675, w_eco136676, w_eco136677, w_eco136678, w_eco136679, w_eco136680, w_eco136681, w_eco136682, w_eco136683, w_eco136684, w_eco136685, w_eco136686, w_eco136687, w_eco136688, w_eco136689, w_eco136690, w_eco136691, w_eco136692, w_eco136693, w_eco136694, w_eco136695, w_eco136696, w_eco136697, w_eco136698, w_eco136699, w_eco136700, w_eco136701, w_eco136702, w_eco136703, w_eco136704, w_eco136705, w_eco136706, w_eco136707, w_eco136708, w_eco136709, w_eco136710, w_eco136711, w_eco136712, w_eco136713, w_eco136714, w_eco136715, w_eco136716, w_eco136717, w_eco136718, w_eco136719, w_eco136720, w_eco136721, w_eco136722, w_eco136723, w_eco136724, w_eco136725, w_eco136726, w_eco136727, w_eco136728, w_eco136729, w_eco136730, w_eco136731, w_eco136732, w_eco136733, w_eco136734, w_eco136735, w_eco136736, w_eco136737, w_eco136738, w_eco136739, w_eco136740, w_eco136741, w_eco136742, w_eco136743, w_eco136744, w_eco136745, w_eco136746, w_eco136747, w_eco136748, w_eco136749, w_eco136750, w_eco136751, w_eco136752, w_eco136753, w_eco136754, w_eco136755, w_eco136756, w_eco136757, w_eco136758, w_eco136759, w_eco136760, w_eco136761, w_eco136762, w_eco136763, w_eco136764, w_eco136765, w_eco136766, w_eco136767, w_eco136768, w_eco136769, w_eco136770, w_eco136771, w_eco136772, w_eco136773, w_eco136774, w_eco136775, w_eco136776, w_eco136777, w_eco136778, w_eco136779, w_eco136780, w_eco136781, w_eco136782, w_eco136783, w_eco136784, w_eco136785, w_eco136786, w_eco136787, w_eco136788, w_eco136789, w_eco136790, w_eco136791, w_eco136792, w_eco136793, w_eco136794, w_eco136795, w_eco136796, w_eco136797, w_eco136798, w_eco136799, w_eco136800, w_eco136801, w_eco136802, w_eco136803, w_eco136804, w_eco136805, w_eco136806, w_eco136807, w_eco136808, w_eco136809, w_eco136810, w_eco136811, w_eco136812, w_eco136813, w_eco136814, w_eco136815, w_eco136816, w_eco136817, w_eco136818, w_eco136819, w_eco136820, w_eco136821, w_eco136822, w_eco136823, w_eco136824, w_eco136825, w_eco136826, w_eco136827, w_eco136828, w_eco136829, w_eco136830, w_eco136831, w_eco136832, w_eco136833, w_eco136834, w_eco136835, w_eco136836, w_eco136837, w_eco136838, w_eco136839, w_eco136840, w_eco136841, w_eco136842, w_eco136843, w_eco136844, w_eco136845, w_eco136846, w_eco136847, w_eco136848, w_eco136849, w_eco136850, w_eco136851, w_eco136852, w_eco136853, w_eco136854, w_eco136855, w_eco136856, w_eco136857, w_eco136858, w_eco136859, w_eco136860, w_eco136861, w_eco136862, w_eco136863, w_eco136864, w_eco136865, w_eco136866, w_eco136867, w_eco136868, w_eco136869, w_eco136870, w_eco136871, w_eco136872, w_eco136873, w_eco136874, w_eco136875, w_eco136876, w_eco136877, w_eco136878, w_eco136879, w_eco136880, w_eco136881, w_eco136882, w_eco136883, w_eco136884, w_eco136885, w_eco136886, w_eco136887, w_eco136888, w_eco136889, w_eco136890, w_eco136891, w_eco136892, w_eco136893, w_eco136894, w_eco136895, w_eco136896, w_eco136897, w_eco136898, w_eco136899, w_eco136900, w_eco136901, w_eco136902, w_eco136903, w_eco136904, w_eco136905, w_eco136906, w_eco136907, w_eco136908, w_eco136909, w_eco136910, w_eco136911, w_eco136912, w_eco136913, w_eco136914, w_eco136915, w_eco136916, w_eco136917, w_eco136918, w_eco136919, w_eco136920, w_eco136921, w_eco136922, w_eco136923, w_eco136924, w_eco136925, w_eco136926, w_eco136927, w_eco136928, w_eco136929, w_eco136930, w_eco136931, w_eco136932, w_eco136933, w_eco136934, w_eco136935, w_eco136936, w_eco136937, w_eco136938, w_eco136939, w_eco136940, w_eco136941, w_eco136942, w_eco136943, w_eco136944, w_eco136945, w_eco136946, w_eco136947, w_eco136948, w_eco136949, w_eco136950, w_eco136951, w_eco136952, w_eco136953, w_eco136954, w_eco136955, w_eco136956, w_eco136957, w_eco136958, w_eco136959, w_eco136960, w_eco136961, w_eco136962, w_eco136963, w_eco136964, w_eco136965, w_eco136966, w_eco136967, w_eco136968, w_eco136969, w_eco136970, w_eco136971, w_eco136972, w_eco136973, w_eco136974, w_eco136975, w_eco136976, w_eco136977, w_eco136978, w_eco136979, w_eco136980, w_eco136981, w_eco136982, w_eco136983, w_eco136984, w_eco136985, w_eco136986, w_eco136987, w_eco136988, w_eco136989, w_eco136990, w_eco136991, w_eco136992, w_eco136993, w_eco136994, w_eco136995, w_eco136996, w_eco136997, w_eco136998, w_eco136999, w_eco137000, w_eco137001, w_eco137002, w_eco137003, w_eco137004, w_eco137005, w_eco137006, w_eco137007, w_eco137008, w_eco137009, w_eco137010, w_eco137011, w_eco137012, w_eco137013, w_eco137014, w_eco137015, w_eco137016, w_eco137017, w_eco137018, w_eco137019, w_eco137020, w_eco137021, w_eco137022, w_eco137023, w_eco137024, w_eco137025, w_eco137026, w_eco137027, w_eco137028, w_eco137029, w_eco137030, w_eco137031, w_eco137032, w_eco137033, w_eco137034, w_eco137035, w_eco137036, w_eco137037, w_eco137038, w_eco137039, w_eco137040, w_eco137041, w_eco137042, w_eco137043, w_eco137044, w_eco137045, w_eco137046, w_eco137047, w_eco137048, w_eco137049, w_eco137050, w_eco137051, w_eco137052, w_eco137053, w_eco137054, w_eco137055, w_eco137056, w_eco137057, w_eco137058, w_eco137059, w_eco137060, w_eco137061, w_eco137062, w_eco137063, w_eco137064, w_eco137065, w_eco137066, w_eco137067, w_eco137068, w_eco137069, w_eco137070, w_eco137071, w_eco137072, w_eco137073, w_eco137074, w_eco137075, w_eco137076, w_eco137077, w_eco137078, w_eco137079, w_eco137080, w_eco137081, w_eco137082, w_eco137083, w_eco137084, w_eco137085, w_eco137086, w_eco137087, w_eco137088, w_eco137089, w_eco137090, w_eco137091, w_eco137092, w_eco137093, w_eco137094, w_eco137095, w_eco137096, w_eco137097, w_eco137098, w_eco137099, w_eco137100, w_eco137101, w_eco137102, w_eco137103, w_eco137104, w_eco137105, w_eco137106, w_eco137107, w_eco137108, w_eco137109, w_eco137110, w_eco137111, w_eco137112, w_eco137113, w_eco137114, w_eco137115, w_eco137116, w_eco137117, w_eco137118, w_eco137119, w_eco137120, w_eco137121, w_eco137122, w_eco137123, w_eco137124, w_eco137125, w_eco137126, w_eco137127, w_eco137128, w_eco137129, w_eco137130, w_eco137131, w_eco137132, w_eco137133, w_eco137134, w_eco137135, w_eco137136, w_eco137137, w_eco137138, w_eco137139, w_eco137140, w_eco137141, w_eco137142, w_eco137143, w_eco137144, w_eco137145, w_eco137146, w_eco137147, w_eco137148, w_eco137149, w_eco137150, w_eco137151, w_eco137152, w_eco137153, w_eco137154, w_eco137155, w_eco137156, w_eco137157, w_eco137158, w_eco137159, w_eco137160, w_eco137161, w_eco137162, w_eco137163, w_eco137164, w_eco137165, w_eco137166, w_eco137167, w_eco137168, w_eco137169, w_eco137170, w_eco137171, w_eco137172, w_eco137173, w_eco137174, w_eco137175, w_eco137176, w_eco137177, w_eco137178, w_eco137179, w_eco137180, w_eco137181, w_eco137182, w_eco137183, w_eco137184, w_eco137185, w_eco137186, w_eco137187, w_eco137188, w_eco137189, w_eco137190, w_eco137191, w_eco137192, w_eco137193, w_eco137194, w_eco137195, w_eco137196, w_eco137197, w_eco137198, w_eco137199, w_eco137200, w_eco137201, w_eco137202, w_eco137203, w_eco137204, w_eco137205, w_eco137206, w_eco137207, w_eco137208, w_eco137209, w_eco137210, w_eco137211, w_eco137212, w_eco137213, w_eco137214, w_eco137215, w_eco137216, w_eco137217, w_eco137218, w_eco137219, w_eco137220, w_eco137221, w_eco137222, w_eco137223, w_eco137224, w_eco137225, w_eco137226, w_eco137227, w_eco137228, w_eco137229, w_eco137230, w_eco137231, w_eco137232, w_eco137233, w_eco137234, w_eco137235, w_eco137236, w_eco137237, w_eco137238, w_eco137239, w_eco137240, w_eco137241, w_eco137242, w_eco137243, w_eco137244, w_eco137245, w_eco137246, w_eco137247, w_eco137248, w_eco137249, w_eco137250, w_eco137251, w_eco137252, w_eco137253, w_eco137254, w_eco137255, w_eco137256, w_eco137257, w_eco137258, w_eco137259, w_eco137260, w_eco137261, w_eco137262, w_eco137263, w_eco137264, w_eco137265, w_eco137266, w_eco137267, w_eco137268, w_eco137269, w_eco137270, w_eco137271, w_eco137272, w_eco137273, w_eco137274, w_eco137275, w_eco137276, w_eco137277, w_eco137278, w_eco137279, w_eco137280, w_eco137281, w_eco137282, w_eco137283, w_eco137284, w_eco137285, w_eco137286, w_eco137287, w_eco137288, w_eco137289, w_eco137290, w_eco137291, w_eco137292, w_eco137293, w_eco137294, w_eco137295, w_eco137296, w_eco137297, w_eco137298, w_eco137299, w_eco137300, w_eco137301, w_eco137302, w_eco137303, w_eco137304, w_eco137305, w_eco137306, w_eco137307, w_eco137308, w_eco137309, w_eco137310, w_eco137311, w_eco137312, w_eco137313, w_eco137314, w_eco137315, w_eco137316, w_eco137317, w_eco137318, w_eco137319, w_eco137320, w_eco137321, w_eco137322, w_eco137323, w_eco137324, w_eco137325, w_eco137326, w_eco137327, w_eco137328, w_eco137329, w_eco137330, w_eco137331, w_eco137332, w_eco137333, w_eco137334, w_eco137335, w_eco137336, w_eco137337, w_eco137338, w_eco137339, w_eco137340, w_eco137341, w_eco137342, w_eco137343, w_eco137344, w_eco137345, w_eco137346, w_eco137347, w_eco137348, w_eco137349, w_eco137350, w_eco137351, w_eco137352, w_eco137353, w_eco137354, w_eco137355, w_eco137356, w_eco137357, w_eco137358, w_eco137359, w_eco137360, w_eco137361, w_eco137362, w_eco137363, w_eco137364, w_eco137365, w_eco137366, w_eco137367, w_eco137368, w_eco137369, w_eco137370, w_eco137371, w_eco137372, w_eco137373, w_eco137374, w_eco137375, w_eco137376, w_eco137377, w_eco137378, w_eco137379, w_eco137380, w_eco137381, w_eco137382, w_eco137383, w_eco137384, w_eco137385, w_eco137386, w_eco137387, w_eco137388, w_eco137389, w_eco137390, w_eco137391, w_eco137392, w_eco137393, w_eco137394, w_eco137395, w_eco137396, w_eco137397, w_eco137398, w_eco137399, w_eco137400, w_eco137401, w_eco137402, w_eco137403, w_eco137404, w_eco137405, w_eco137406, w_eco137407, w_eco137408, w_eco137409, w_eco137410, w_eco137411, w_eco137412, w_eco137413, w_eco137414, w_eco137415, w_eco137416, w_eco137417, w_eco137418, w_eco137419, w_eco137420, w_eco137421, w_eco137422, w_eco137423, w_eco137424, w_eco137425, w_eco137426, w_eco137427, w_eco137428, w_eco137429, w_eco137430, w_eco137431, w_eco137432, w_eco137433, w_eco137434, w_eco137435, w_eco137436, w_eco137437, w_eco137438, w_eco137439, w_eco137440, w_eco137441, w_eco137442, w_eco137443, w_eco137444, w_eco137445, w_eco137446, w_eco137447, w_eco137448, w_eco137449, w_eco137450, w_eco137451, w_eco137452, w_eco137453, w_eco137454, w_eco137455, w_eco137456, w_eco137457, w_eco137458, w_eco137459, w_eco137460, w_eco137461, w_eco137462, w_eco137463, w_eco137464, w_eco137465, w_eco137466, w_eco137467, w_eco137468, w_eco137469, w_eco137470, w_eco137471, w_eco137472, w_eco137473, w_eco137474, w_eco137475, w_eco137476, w_eco137477, w_eco137478, w_eco137479, w_eco137480, w_eco137481, w_eco137482, w_eco137483, w_eco137484, w_eco137485, w_eco137486, w_eco137487, w_eco137488, w_eco137489, w_eco137490, w_eco137491, w_eco137492, w_eco137493, w_eco137494, w_eco137495, w_eco137496, w_eco137497, w_eco137498, w_eco137499, w_eco137500, w_eco137501, w_eco137502, w_eco137503, w_eco137504, w_eco137505, w_eco137506, w_eco137507, w_eco137508, w_eco137509, w_eco137510, w_eco137511, w_eco137512, w_eco137513, w_eco137514, w_eco137515, w_eco137516, w_eco137517, w_eco137518, w_eco137519, w_eco137520, w_eco137521, w_eco137522, w_eco137523, w_eco137524, w_eco137525, w_eco137526, w_eco137527, w_eco137528, w_eco137529, w_eco137530, w_eco137531, w_eco137532, w_eco137533, w_eco137534, w_eco137535, w_eco137536, w_eco137537, w_eco137538, w_eco137539, w_eco137540, w_eco137541, w_eco137542, w_eco137543, w_eco137544, w_eco137545, w_eco137546, w_eco137547, w_eco137548, w_eco137549, w_eco137550, w_eco137551, w_eco137552, w_eco137553, w_eco137554, w_eco137555, w_eco137556, w_eco137557, w_eco137558, w_eco137559, w_eco137560, w_eco137561, w_eco137562, w_eco137563, w_eco137564, w_eco137565, w_eco137566, w_eco137567, w_eco137568, w_eco137569, w_eco137570, w_eco137571, w_eco137572, w_eco137573, w_eco137574, w_eco137575, w_eco137576, w_eco137577, w_eco137578, w_eco137579, w_eco137580, w_eco137581, w_eco137582, w_eco137583, w_eco137584, w_eco137585, w_eco137586, w_eco137587, w_eco137588, w_eco137589, w_eco137590, w_eco137591, w_eco137592, w_eco137593, w_eco137594, w_eco137595, w_eco137596, w_eco137597, w_eco137598, w_eco137599, w_eco137600, w_eco137601, w_eco137602, w_eco137603, w_eco137604, w_eco137605, w_eco137606, w_eco137607, w_eco137608, w_eco137609, w_eco137610, w_eco137611, w_eco137612, w_eco137613, w_eco137614, w_eco137615, w_eco137616, w_eco137617, w_eco137618, w_eco137619, w_eco137620, w_eco137621, w_eco137622, w_eco137623, w_eco137624, w_eco137625, w_eco137626, w_eco137627, w_eco137628, w_eco137629, w_eco137630, w_eco137631, w_eco137632, w_eco137633, w_eco137634, w_eco137635, w_eco137636, w_eco137637, w_eco137638, w_eco137639, w_eco137640, w_eco137641, w_eco137642, w_eco137643, w_eco137644, w_eco137645, w_eco137646, w_eco137647, w_eco137648, w_eco137649, w_eco137650, w_eco137651, w_eco137652, w_eco137653, w_eco137654, w_eco137655, w_eco137656, w_eco137657, w_eco137658, w_eco137659, w_eco137660, w_eco137661, w_eco137662, w_eco137663, w_eco137664, w_eco137665, w_eco137666, w_eco137667, w_eco137668, w_eco137669, w_eco137670, w_eco137671, w_eco137672, w_eco137673, w_eco137674, w_eco137675, w_eco137676, w_eco137677, w_eco137678, w_eco137679, w_eco137680, w_eco137681, w_eco137682, w_eco137683, w_eco137684, w_eco137685, w_eco137686, w_eco137687, w_eco137688, w_eco137689, w_eco137690, w_eco137691, w_eco137692, w_eco137693, w_eco137694, w_eco137695, w_eco137696, w_eco137697, w_eco137698, w_eco137699, w_eco137700, w_eco137701, w_eco137702, w_eco137703, w_eco137704, w_eco137705, w_eco137706, w_eco137707, w_eco137708, w_eco137709, w_eco137710, w_eco137711, w_eco137712, w_eco137713, w_eco137714, w_eco137715, w_eco137716, w_eco137717, w_eco137718, w_eco137719, w_eco137720, w_eco137721, w_eco137722, w_eco137723, w_eco137724, w_eco137725, w_eco137726, w_eco137727, w_eco137728, w_eco137729, w_eco137730, w_eco137731, w_eco137732, w_eco137733, w_eco137734, w_eco137735, w_eco137736, w_eco137737, w_eco137738, w_eco137739, w_eco137740, w_eco137741, w_eco137742, w_eco137743, w_eco137744, w_eco137745, w_eco137746, w_eco137747, w_eco137748, w_eco137749, w_eco137750, w_eco137751, w_eco137752, w_eco137753, w_eco137754, w_eco137755, w_eco137756, w_eco137757, w_eco137758, w_eco137759, w_eco137760, w_eco137761, w_eco137762, w_eco137763, w_eco137764, w_eco137765, w_eco137766, w_eco137767, w_eco137768, w_eco137769, w_eco137770, w_eco137771, w_eco137772, w_eco137773, w_eco137774, w_eco137775, w_eco137776, w_eco137777, w_eco137778, w_eco137779, w_eco137780, w_eco137781, w_eco137782, w_eco137783, w_eco137784, w_eco137785, w_eco137786, w_eco137787, w_eco137788, w_eco137789, w_eco137790, w_eco137791, w_eco137792, w_eco137793, w_eco137794, w_eco137795, w_eco137796, w_eco137797, w_eco137798, w_eco137799, w_eco137800, w_eco137801, w_eco137802, w_eco137803, w_eco137804, w_eco137805, w_eco137806, w_eco137807, w_eco137808, w_eco137809, w_eco137810, w_eco137811, w_eco137812, w_eco137813, w_eco137814, w_eco137815, w_eco137816, w_eco137817, w_eco137818, w_eco137819, w_eco137820, w_eco137821, w_eco137822, w_eco137823, w_eco137824, w_eco137825, w_eco137826, w_eco137827, w_eco137828, w_eco137829, w_eco137830, w_eco137831, w_eco137832, w_eco137833, w_eco137834, w_eco137835, w_eco137836, w_eco137837, w_eco137838, w_eco137839, w_eco137840, w_eco137841, w_eco137842, w_eco137843, w_eco137844, w_eco137845, w_eco137846, w_eco137847, w_eco137848, w_eco137849, w_eco137850, w_eco137851, w_eco137852, w_eco137853, w_eco137854, w_eco137855, w_eco137856, w_eco137857, w_eco137858, w_eco137859, w_eco137860, w_eco137861, w_eco137862, w_eco137863, w_eco137864, w_eco137865, w_eco137866, w_eco137867, w_eco137868, w_eco137869, w_eco137870, w_eco137871, w_eco137872, w_eco137873, w_eco137874, w_eco137875, w_eco137876, w_eco137877, w_eco137878, w_eco137879, w_eco137880, w_eco137881, w_eco137882, w_eco137883, w_eco137884, w_eco137885, w_eco137886, w_eco137887, w_eco137888, w_eco137889, w_eco137890, w_eco137891, w_eco137892, w_eco137893, w_eco137894, w_eco137895, w_eco137896, w_eco137897, w_eco137898, w_eco137899, w_eco137900, w_eco137901, w_eco137902, w_eco137903, w_eco137904, w_eco137905, w_eco137906, w_eco137907, w_eco137908, w_eco137909, w_eco137910, w_eco137911, w_eco137912, w_eco137913, w_eco137914, w_eco137915, w_eco137916, w_eco137917, w_eco137918, w_eco137919, w_eco137920, w_eco137921, w_eco137922, w_eco137923, w_eco137924, w_eco137925, w_eco137926, w_eco137927, w_eco137928, w_eco137929, w_eco137930, w_eco137931, w_eco137932, w_eco137933, w_eco137934, w_eco137935, w_eco137936, w_eco137937, w_eco137938, w_eco137939, w_eco137940, w_eco137941, w_eco137942, w_eco137943, w_eco137944, w_eco137945, w_eco137946, w_eco137947, w_eco137948, w_eco137949, w_eco137950, w_eco137951, w_eco137952, w_eco137953, w_eco137954, w_eco137955, w_eco137956, w_eco137957, w_eco137958, w_eco137959, w_eco137960, w_eco137961, w_eco137962, w_eco137963, w_eco137964, w_eco137965, w_eco137966, w_eco137967, w_eco137968, w_eco137969, w_eco137970, w_eco137971, w_eco137972, w_eco137973, w_eco137974, w_eco137975, w_eco137976, w_eco137977, w_eco137978, w_eco137979, w_eco137980, w_eco137981, w_eco137982, w_eco137983, w_eco137984, w_eco137985, w_eco137986, w_eco137987, w_eco137988, w_eco137989, w_eco137990, w_eco137991, w_eco137992, w_eco137993, w_eco137994, w_eco137995, w_eco137996, w_eco137997, w_eco137998, w_eco137999, w_eco138000, w_eco138001, w_eco138002, w_eco138003, w_eco138004, w_eco138005, w_eco138006, w_eco138007, w_eco138008, w_eco138009, w_eco138010, w_eco138011, w_eco138012, w_eco138013, w_eco138014, w_eco138015, w_eco138016, w_eco138017, w_eco138018, w_eco138019, w_eco138020, w_eco138021, w_eco138022, w_eco138023, w_eco138024, w_eco138025, w_eco138026, w_eco138027, w_eco138028, w_eco138029, w_eco138030, w_eco138031, w_eco138032, w_eco138033, w_eco138034, w_eco138035, w_eco138036, w_eco138037, w_eco138038, w_eco138039, w_eco138040, w_eco138041, w_eco138042, w_eco138043, w_eco138044, w_eco138045, w_eco138046, w_eco138047, w_eco138048, w_eco138049, w_eco138050, w_eco138051, w_eco138052, w_eco138053, w_eco138054, w_eco138055, w_eco138056, w_eco138057, w_eco138058, w_eco138059, w_eco138060, w_eco138061, w_eco138062, w_eco138063, w_eco138064, w_eco138065, w_eco138066, w_eco138067, w_eco138068, w_eco138069, w_eco138070, w_eco138071, w_eco138072, w_eco138073, w_eco138074, w_eco138075, w_eco138076, w_eco138077, w_eco138078, w_eco138079, w_eco138080, w_eco138081, w_eco138082, w_eco138083, w_eco138084, w_eco138085, w_eco138086, w_eco138087, w_eco138088, w_eco138089, w_eco138090, w_eco138091, w_eco138092, w_eco138093, w_eco138094, w_eco138095, w_eco138096, w_eco138097, w_eco138098, w_eco138099, w_eco138100, w_eco138101, w_eco138102, w_eco138103, w_eco138104, w_eco138105, w_eco138106, w_eco138107, w_eco138108, w_eco138109, w_eco138110, w_eco138111, w_eco138112, w_eco138113, w_eco138114, w_eco138115, w_eco138116, w_eco138117, w_eco138118, w_eco138119, w_eco138120, w_eco138121, w_eco138122, w_eco138123, w_eco138124, w_eco138125, w_eco138126, w_eco138127, w_eco138128, w_eco138129, w_eco138130, w_eco138131, w_eco138132, w_eco138133, w_eco138134, w_eco138135, w_eco138136, w_eco138137, w_eco138138, w_eco138139, w_eco138140, w_eco138141, w_eco138142, w_eco138143, w_eco138144, w_eco138145, w_eco138146, w_eco138147, w_eco138148, w_eco138149, w_eco138150, w_eco138151, w_eco138152, w_eco138153, w_eco138154, w_eco138155, w_eco138156, w_eco138157, w_eco138158, w_eco138159, w_eco138160, w_eco138161, w_eco138162, w_eco138163, w_eco138164, w_eco138165, w_eco138166, w_eco138167, w_eco138168, w_eco138169, w_eco138170, w_eco138171, w_eco138172, w_eco138173, w_eco138174, w_eco138175, w_eco138176, w_eco138177, w_eco138178, w_eco138179, w_eco138180, w_eco138181, w_eco138182, w_eco138183, w_eco138184, w_eco138185, w_eco138186, w_eco138187, w_eco138188, w_eco138189, w_eco138190, w_eco138191, w_eco138192, w_eco138193, w_eco138194, w_eco138195, w_eco138196, w_eco138197, w_eco138198, w_eco138199, w_eco138200, w_eco138201, w_eco138202, w_eco138203, w_eco138204, w_eco138205, w_eco138206, w_eco138207, w_eco138208, w_eco138209, w_eco138210, w_eco138211, w_eco138212, w_eco138213, w_eco138214, w_eco138215, w_eco138216, w_eco138217, w_eco138218, w_eco138219, w_eco138220, w_eco138221, w_eco138222, w_eco138223, w_eco138224, w_eco138225, w_eco138226, w_eco138227, w_eco138228, w_eco138229, w_eco138230, w_eco138231, w_eco138232, w_eco138233, w_eco138234, w_eco138235, w_eco138236, w_eco138237, w_eco138238, w_eco138239, w_eco138240, w_eco138241, w_eco138242, w_eco138243, w_eco138244, w_eco138245, w_eco138246, w_eco138247, w_eco138248, w_eco138249, w_eco138250, w_eco138251, w_eco138252, w_eco138253, w_eco138254, w_eco138255, w_eco138256, w_eco138257, w_eco138258, w_eco138259, w_eco138260, w_eco138261, w_eco138262, w_eco138263, w_eco138264, w_eco138265, w_eco138266, w_eco138267, w_eco138268, w_eco138269, w_eco138270, w_eco138271, w_eco138272, w_eco138273, w_eco138274, w_eco138275, w_eco138276, w_eco138277, w_eco138278, w_eco138279, w_eco138280, w_eco138281, w_eco138282, w_eco138283, w_eco138284, w_eco138285, w_eco138286, w_eco138287, w_eco138288, w_eco138289, w_eco138290, w_eco138291, w_eco138292, w_eco138293, w_eco138294, w_eco138295, w_eco138296, w_eco138297, w_eco138298, w_eco138299, w_eco138300, w_eco138301, w_eco138302, w_eco138303, w_eco138304, w_eco138305, w_eco138306, w_eco138307, w_eco138308, w_eco138309, w_eco138310, w_eco138311, w_eco138312, w_eco138313, w_eco138314, w_eco138315, w_eco138316, w_eco138317, w_eco138318, w_eco138319, w_eco138320, w_eco138321, w_eco138322, w_eco138323, w_eco138324, w_eco138325, w_eco138326, w_eco138327, w_eco138328, w_eco138329, w_eco138330, w_eco138331, w_eco138332, w_eco138333, w_eco138334, w_eco138335, w_eco138336, w_eco138337, w_eco138338, w_eco138339, w_eco138340, w_eco138341, w_eco138342, w_eco138343, w_eco138344, w_eco138345, w_eco138346, w_eco138347, w_eco138348, w_eco138349, w_eco138350, w_eco138351, w_eco138352, w_eco138353, w_eco138354, w_eco138355, w_eco138356, w_eco138357, w_eco138358, w_eco138359, w_eco138360, w_eco138361, w_eco138362, w_eco138363, w_eco138364, w_eco138365, w_eco138366, w_eco138367, w_eco138368, w_eco138369, w_eco138370, w_eco138371, w_eco138372, w_eco138373, w_eco138374, w_eco138375, w_eco138376, w_eco138377, w_eco138378, w_eco138379, w_eco138380, w_eco138381, w_eco138382, w_eco138383, w_eco138384, w_eco138385, w_eco138386, w_eco138387, w_eco138388, w_eco138389, w_eco138390, w_eco138391, w_eco138392, w_eco138393, w_eco138394, w_eco138395, w_eco138396, w_eco138397, w_eco138398, w_eco138399, w_eco138400, w_eco138401, w_eco138402, w_eco138403, w_eco138404, w_eco138405, w_eco138406, w_eco138407, w_eco138408, w_eco138409, w_eco138410, w_eco138411, w_eco138412, w_eco138413, w_eco138414, w_eco138415, w_eco138416, w_eco138417, w_eco138418, w_eco138419, w_eco138420, w_eco138421, w_eco138422, w_eco138423, w_eco138424, w_eco138425, w_eco138426, w_eco138427, w_eco138428, w_eco138429, w_eco138430, w_eco138431, w_eco138432, w_eco138433, w_eco138434, w_eco138435, w_eco138436, w_eco138437, w_eco138438, w_eco138439, w_eco138440, w_eco138441, w_eco138442, w_eco138443, w_eco138444, w_eco138445, w_eco138446, w_eco138447, w_eco138448, w_eco138449, w_eco138450, w_eco138451, w_eco138452, w_eco138453, w_eco138454, w_eco138455, w_eco138456, w_eco138457, w_eco138458, w_eco138459, w_eco138460, w_eco138461, w_eco138462, w_eco138463, w_eco138464, w_eco138465, w_eco138466, w_eco138467, w_eco138468, w_eco138469, w_eco138470, w_eco138471, w_eco138472, w_eco138473, w_eco138474, w_eco138475, w_eco138476, w_eco138477, w_eco138478, w_eco138479, w_eco138480, w_eco138481, w_eco138482, w_eco138483, w_eco138484, w_eco138485, w_eco138486, w_eco138487, w_eco138488, w_eco138489, w_eco138490, w_eco138491, w_eco138492, w_eco138493, w_eco138494, w_eco138495, w_eco138496, w_eco138497, w_eco138498, w_eco138499, w_eco138500, w_eco138501, w_eco138502, w_eco138503, w_eco138504, w_eco138505, w_eco138506, w_eco138507, w_eco138508, w_eco138509, w_eco138510, w_eco138511, w_eco138512, w_eco138513, w_eco138514, w_eco138515, w_eco138516, w_eco138517, w_eco138518, w_eco138519, w_eco138520, w_eco138521, w_eco138522, w_eco138523, w_eco138524, w_eco138525, w_eco138526, w_eco138527, w_eco138528, w_eco138529, w_eco138530, w_eco138531, w_eco138532, w_eco138533, w_eco138534, w_eco138535, w_eco138536, w_eco138537, w_eco138538, w_eco138539, w_eco138540, w_eco138541, w_eco138542, w_eco138543, w_eco138544, w_eco138545, w_eco138546, w_eco138547, w_eco138548, w_eco138549, w_eco138550, w_eco138551, w_eco138552, w_eco138553, w_eco138554, w_eco138555, w_eco138556, w_eco138557, w_eco138558, w_eco138559, w_eco138560, w_eco138561, w_eco138562, w_eco138563, w_eco138564, w_eco138565, w_eco138566, w_eco138567, w_eco138568, w_eco138569, w_eco138570, w_eco138571, w_eco138572, w_eco138573, w_eco138574, w_eco138575, w_eco138576, w_eco138577, w_eco138578, w_eco138579, w_eco138580, w_eco138581, w_eco138582, w_eco138583, w_eco138584, w_eco138585, w_eco138586, w_eco138587, w_eco138588, w_eco138589, w_eco138590, w_eco138591, w_eco138592, w_eco138593, w_eco138594, w_eco138595, w_eco138596, w_eco138597, w_eco138598, w_eco138599, w_eco138600, w_eco138601, w_eco138602, w_eco138603, w_eco138604, w_eco138605, w_eco138606, w_eco138607, w_eco138608, w_eco138609, w_eco138610, w_eco138611, w_eco138612, w_eco138613, w_eco138614, w_eco138615, w_eco138616, w_eco138617, w_eco138618, w_eco138619, w_eco138620, w_eco138621, w_eco138622, w_eco138623, w_eco138624, w_eco138625, w_eco138626, w_eco138627, w_eco138628, w_eco138629, w_eco138630, w_eco138631, w_eco138632, w_eco138633, w_eco138634, w_eco138635, w_eco138636, w_eco138637, w_eco138638, w_eco138639, w_eco138640, w_eco138641, w_eco138642, w_eco138643, w_eco138644, w_eco138645, w_eco138646, w_eco138647, w_eco138648, w_eco138649, w_eco138650, w_eco138651, w_eco138652, w_eco138653, w_eco138654, w_eco138655, w_eco138656, w_eco138657, w_eco138658, w_eco138659, w_eco138660, w_eco138661, w_eco138662, w_eco138663, w_eco138664, w_eco138665, w_eco138666, w_eco138667, w_eco138668, w_eco138669, w_eco138670, w_eco138671, w_eco138672, w_eco138673, w_eco138674, w_eco138675, w_eco138676, w_eco138677, w_eco138678, w_eco138679, w_eco138680, w_eco138681, w_eco138682, w_eco138683, w_eco138684, w_eco138685, w_eco138686, w_eco138687, w_eco138688, w_eco138689, w_eco138690, w_eco138691, w_eco138692, w_eco138693, w_eco138694, w_eco138695, w_eco138696, w_eco138697, w_eco138698, w_eco138699, w_eco138700, w_eco138701, w_eco138702, w_eco138703, w_eco138704, w_eco138705, w_eco138706, w_eco138707, w_eco138708, w_eco138709, w_eco138710, w_eco138711, w_eco138712, w_eco138713, w_eco138714, w_eco138715, w_eco138716, w_eco138717, w_eco138718, w_eco138719, w_eco138720, w_eco138721, w_eco138722, w_eco138723, w_eco138724, w_eco138725, w_eco138726, w_eco138727, w_eco138728, w_eco138729, w_eco138730, w_eco138731, w_eco138732, w_eco138733, w_eco138734, w_eco138735, w_eco138736, w_eco138737, w_eco138738, w_eco138739, w_eco138740, w_eco138741, w_eco138742, w_eco138743, w_eco138744, w_eco138745, w_eco138746, w_eco138747, w_eco138748, w_eco138749, w_eco138750, w_eco138751, w_eco138752, w_eco138753, w_eco138754, w_eco138755, w_eco138756, w_eco138757, w_eco138758, w_eco138759, w_eco138760, w_eco138761, w_eco138762, w_eco138763, w_eco138764, w_eco138765, w_eco138766, w_eco138767, w_eco138768, w_eco138769, w_eco138770, w_eco138771, w_eco138772, w_eco138773, w_eco138774, w_eco138775, w_eco138776, w_eco138777, w_eco138778, w_eco138779, w_eco138780, w_eco138781, w_eco138782, w_eco138783, w_eco138784, w_eco138785, w_eco138786, w_eco138787, w_eco138788, w_eco138789, w_eco138790, w_eco138791, w_eco138792, w_eco138793, w_eco138794, w_eco138795, w_eco138796, w_eco138797, w_eco138798, w_eco138799, w_eco138800, w_eco138801, w_eco138802, w_eco138803, w_eco138804, w_eco138805, w_eco138806, w_eco138807, w_eco138808, w_eco138809, w_eco138810, w_eco138811, w_eco138812, w_eco138813, w_eco138814, w_eco138815, w_eco138816, w_eco138817, w_eco138818, w_eco138819, w_eco138820, w_eco138821, w_eco138822, w_eco138823, w_eco138824, w_eco138825, w_eco138826, w_eco138827, w_eco138828, w_eco138829, w_eco138830, w_eco138831, w_eco138832, w_eco138833, w_eco138834, w_eco138835, w_eco138836, w_eco138837, w_eco138838, w_eco138839, w_eco138840, w_eco138841, w_eco138842, w_eco138843, w_eco138844, w_eco138845, w_eco138846, w_eco138847, w_eco138848, w_eco138849, w_eco138850, w_eco138851, w_eco138852, w_eco138853, w_eco138854, w_eco138855, w_eco138856, w_eco138857, w_eco138858, w_eco138859, w_eco138860, w_eco138861, w_eco138862, w_eco138863, w_eco138864, w_eco138865, w_eco138866, w_eco138867, w_eco138868, w_eco138869, w_eco138870, w_eco138871, w_eco138872, w_eco138873, w_eco138874, w_eco138875, w_eco138876, w_eco138877, w_eco138878, w_eco138879, w_eco138880, w_eco138881, w_eco138882, w_eco138883, w_eco138884, w_eco138885, w_eco138886, w_eco138887, w_eco138888, w_eco138889, w_eco138890, w_eco138891, w_eco138892, w_eco138893, w_eco138894, w_eco138895, w_eco138896, w_eco138897, w_eco138898, w_eco138899, w_eco138900, w_eco138901, w_eco138902, w_eco138903, w_eco138904, w_eco138905, w_eco138906, w_eco138907, w_eco138908, w_eco138909, w_eco138910, w_eco138911, w_eco138912, w_eco138913, w_eco138914, w_eco138915, w_eco138916, w_eco138917, w_eco138918, w_eco138919, w_eco138920, w_eco138921, w_eco138922, w_eco138923, w_eco138924, w_eco138925, w_eco138926, w_eco138927, w_eco138928, w_eco138929, w_eco138930, w_eco138931, w_eco138932, w_eco138933, w_eco138934, w_eco138935, w_eco138936, w_eco138937, w_eco138938, w_eco138939, w_eco138940, w_eco138941, w_eco138942, w_eco138943, w_eco138944, w_eco138945, w_eco138946, w_eco138947, w_eco138948, w_eco138949, w_eco138950, w_eco138951, w_eco138952, w_eco138953, w_eco138954, w_eco138955, w_eco138956, w_eco138957, w_eco138958, w_eco138959, w_eco138960, w_eco138961, w_eco138962, w_eco138963, w_eco138964, w_eco138965, w_eco138966, w_eco138967, w_eco138968, w_eco138969, w_eco138970, w_eco138971, w_eco138972, w_eco138973, w_eco138974, w_eco138975, w_eco138976, w_eco138977, w_eco138978, w_eco138979, w_eco138980, w_eco138981, w_eco138982, w_eco138983, w_eco138984, w_eco138985, w_eco138986, w_eco138987, w_eco138988, w_eco138989, w_eco138990, w_eco138991, w_eco138992, w_eco138993, w_eco138994, w_eco138995, w_eco138996, w_eco138997, w_eco138998, w_eco138999, w_eco139000, w_eco139001, w_eco139002, w_eco139003, w_eco139004, w_eco139005, w_eco139006, w_eco139007, w_eco139008, w_eco139009, w_eco139010, w_eco139011, w_eco139012, w_eco139013, w_eco139014, w_eco139015, w_eco139016, w_eco139017, w_eco139018, w_eco139019, w_eco139020, w_eco139021, w_eco139022, w_eco139023, w_eco139024, w_eco139025, w_eco139026, w_eco139027, w_eco139028, w_eco139029, w_eco139030, w_eco139031, w_eco139032, w_eco139033, w_eco139034, w_eco139035, w_eco139036, w_eco139037, w_eco139038, w_eco139039, w_eco139040, w_eco139041, w_eco139042, w_eco139043, w_eco139044, w_eco139045, w_eco139046, w_eco139047, w_eco139048, w_eco139049, w_eco139050, w_eco139051, w_eco139052, w_eco139053, w_eco139054, w_eco139055, w_eco139056, w_eco139057, w_eco139058, w_eco139059, w_eco139060, w_eco139061, w_eco139062, w_eco139063, w_eco139064, w_eco139065, w_eco139066, w_eco139067, w_eco139068, w_eco139069, w_eco139070, w_eco139071, w_eco139072, w_eco139073, w_eco139074, w_eco139075, w_eco139076, w_eco139077, w_eco139078, w_eco139079, w_eco139080, w_eco139081, w_eco139082, w_eco139083, w_eco139084, w_eco139085, w_eco139086, w_eco139087, w_eco139088, w_eco139089, w_eco139090, w_eco139091, w_eco139092, w_eco139093, w_eco139094, w_eco139095, w_eco139096, w_eco139097, w_eco139098, w_eco139099, w_eco139100, w_eco139101, w_eco139102, w_eco139103, w_eco139104, w_eco139105, w_eco139106, w_eco139107, w_eco139108, w_eco139109, w_eco139110, w_eco139111, w_eco139112, w_eco139113, w_eco139114, w_eco139115, w_eco139116, w_eco139117, w_eco139118, w_eco139119, w_eco139120, w_eco139121, w_eco139122, w_eco139123, w_eco139124, w_eco139125, w_eco139126, w_eco139127, w_eco139128, w_eco139129, w_eco139130, w_eco139131, w_eco139132, w_eco139133, w_eco139134, w_eco139135, w_eco139136, w_eco139137, w_eco139138, w_eco139139, w_eco139140, w_eco139141, w_eco139142, w_eco139143, w_eco139144, w_eco139145, w_eco139146, w_eco139147, w_eco139148, w_eco139149, w_eco139150, w_eco139151, w_eco139152, w_eco139153, w_eco139154, w_eco139155, w_eco139156, w_eco139157, w_eco139158, w_eco139159, w_eco139160, w_eco139161, w_eco139162, w_eco139163, w_eco139164, w_eco139165, w_eco139166, w_eco139167, w_eco139168, w_eco139169, w_eco139170, w_eco139171, w_eco139172, w_eco139173, w_eco139174, w_eco139175, w_eco139176, w_eco139177, w_eco139178, w_eco139179, w_eco139180, w_eco139181, w_eco139182, w_eco139183, w_eco139184, w_eco139185, w_eco139186, w_eco139187, w_eco139188, w_eco139189, w_eco139190, w_eco139191, w_eco139192, w_eco139193, w_eco139194, w_eco139195, w_eco139196, w_eco139197, w_eco139198, w_eco139199, w_eco139200, w_eco139201, w_eco139202, w_eco139203, w_eco139204, w_eco139205, w_eco139206, w_eco139207, w_eco139208, w_eco139209, w_eco139210, w_eco139211, w_eco139212, w_eco139213, w_eco139214, w_eco139215, w_eco139216, w_eco139217, w_eco139218, w_eco139219, w_eco139220, w_eco139221, w_eco139222, w_eco139223, w_eco139224, w_eco139225, w_eco139226, w_eco139227, w_eco139228, w_eco139229, w_eco139230, w_eco139231, w_eco139232, w_eco139233, w_eco139234, w_eco139235, w_eco139236, w_eco139237, w_eco139238, w_eco139239, w_eco139240, w_eco139241, w_eco139242, w_eco139243, w_eco139244, w_eco139245, w_eco139246, w_eco139247, w_eco139248, w_eco139249, w_eco139250, w_eco139251, w_eco139252, w_eco139253, w_eco139254, w_eco139255, w_eco139256, w_eco139257, w_eco139258, w_eco139259, w_eco139260, w_eco139261, w_eco139262, w_eco139263, w_eco139264, w_eco139265, w_eco139266, w_eco139267, w_eco139268, w_eco139269, w_eco139270, w_eco139271, w_eco139272, w_eco139273, w_eco139274, w_eco139275, w_eco139276, w_eco139277, w_eco139278, w_eco139279, w_eco139280, w_eco139281, w_eco139282, w_eco139283, w_eco139284, w_eco139285, w_eco139286, w_eco139287, w_eco139288, w_eco139289, w_eco139290, w_eco139291, w_eco139292, w_eco139293, w_eco139294, w_eco139295, w_eco139296, w_eco139297, w_eco139298, w_eco139299, w_eco139300, w_eco139301, w_eco139302, w_eco139303, w_eco139304, w_eco139305, w_eco139306, w_eco139307, w_eco139308, w_eco139309, w_eco139310, w_eco139311, w_eco139312, w_eco139313, w_eco139314, w_eco139315, w_eco139316, w_eco139317, w_eco139318, w_eco139319, w_eco139320, w_eco139321, w_eco139322, w_eco139323, w_eco139324, w_eco139325, w_eco139326, w_eco139327, w_eco139328, w_eco139329, w_eco139330, w_eco139331, w_eco139332, w_eco139333, w_eco139334, w_eco139335, w_eco139336, w_eco139337, w_eco139338, w_eco139339, w_eco139340, w_eco139341, w_eco139342, w_eco139343, w_eco139344, w_eco139345, w_eco139346, w_eco139347, w_eco139348, w_eco139349, w_eco139350, w_eco139351, w_eco139352, w_eco139353, w_eco139354, w_eco139355, w_eco139356, w_eco139357, w_eco139358, w_eco139359, w_eco139360, w_eco139361, w_eco139362, w_eco139363, w_eco139364, w_eco139365, w_eco139366, w_eco139367, w_eco139368, w_eco139369, w_eco139370, w_eco139371, w_eco139372, w_eco139373, w_eco139374, w_eco139375, w_eco139376, w_eco139377, w_eco139378, w_eco139379, w_eco139380, w_eco139381, w_eco139382, w_eco139383, w_eco139384, w_eco139385, w_eco139386, w_eco139387, w_eco139388, w_eco139389, w_eco139390, w_eco139391, w_eco139392, w_eco139393, w_eco139394, w_eco139395, w_eco139396, w_eco139397, w_eco139398, w_eco139399, w_eco139400, w_eco139401, w_eco139402, w_eco139403, w_eco139404, w_eco139405, w_eco139406, w_eco139407, w_eco139408, w_eco139409, w_eco139410, w_eco139411, w_eco139412, w_eco139413, w_eco139414, w_eco139415, w_eco139416, w_eco139417, w_eco139418, w_eco139419, w_eco139420, w_eco139421, w_eco139422, w_eco139423, w_eco139424, w_eco139425, w_eco139426, w_eco139427, w_eco139428, w_eco139429, w_eco139430, w_eco139431, w_eco139432, w_eco139433, w_eco139434, w_eco139435, w_eco139436, w_eco139437, w_eco139438, w_eco139439, w_eco139440, w_eco139441, w_eco139442, w_eco139443, w_eco139444, w_eco139445, w_eco139446, w_eco139447, w_eco139448, w_eco139449, w_eco139450, w_eco139451, w_eco139452, w_eco139453, w_eco139454, w_eco139455, w_eco139456, w_eco139457, w_eco139458, w_eco139459, w_eco139460, w_eco139461, w_eco139462, w_eco139463, w_eco139464, w_eco139465, w_eco139466, w_eco139467, w_eco139468, w_eco139469, w_eco139470, w_eco139471, w_eco139472, w_eco139473, w_eco139474, w_eco139475, w_eco139476, w_eco139477, w_eco139478, w_eco139479, w_eco139480, w_eco139481, w_eco139482, w_eco139483, w_eco139484, w_eco139485, w_eco139486, w_eco139487, w_eco139488, w_eco139489, w_eco139490, w_eco139491, w_eco139492, w_eco139493, w_eco139494, w_eco139495, w_eco139496, w_eco139497, w_eco139498, w_eco139499, w_eco139500, w_eco139501, w_eco139502, w_eco139503, w_eco139504, w_eco139505, w_eco139506, w_eco139507, w_eco139508, w_eco139509, w_eco139510, w_eco139511, w_eco139512, w_eco139513, w_eco139514, w_eco139515, w_eco139516, w_eco139517, w_eco139518, w_eco139519, w_eco139520, w_eco139521, w_eco139522, w_eco139523, w_eco139524, w_eco139525, w_eco139526, w_eco139527, w_eco139528, w_eco139529, w_eco139530, w_eco139531, w_eco139532, w_eco139533, w_eco139534, w_eco139535, w_eco139536, w_eco139537, w_eco139538, w_eco139539, w_eco139540, w_eco139541, w_eco139542, w_eco139543, w_eco139544, w_eco139545, w_eco139546, w_eco139547, w_eco139548, w_eco139549, w_eco139550, w_eco139551, w_eco139552, w_eco139553, w_eco139554, w_eco139555, w_eco139556, w_eco139557, w_eco139558, w_eco139559, w_eco139560, w_eco139561, w_eco139562, w_eco139563, w_eco139564, w_eco139565, w_eco139566, w_eco139567, w_eco139568, w_eco139569, w_eco139570, w_eco139571, w_eco139572, w_eco139573, w_eco139574, w_eco139575, w_eco139576, w_eco139577, w_eco139578, w_eco139579, w_eco139580, w_eco139581, w_eco139582, w_eco139583, w_eco139584, w_eco139585, w_eco139586, w_eco139587, w_eco139588, w_eco139589, w_eco139590, w_eco139591, w_eco139592, w_eco139593, w_eco139594, w_eco139595, w_eco139596, w_eco139597, w_eco139598, w_eco139599, w_eco139600, w_eco139601, w_eco139602, w_eco139603, w_eco139604, w_eco139605, w_eco139606, w_eco139607, w_eco139608, w_eco139609, w_eco139610, w_eco139611, w_eco139612, w_eco139613, w_eco139614, w_eco139615, w_eco139616, w_eco139617, w_eco139618, w_eco139619, w_eco139620, w_eco139621, w_eco139622, w_eco139623, w_eco139624, w_eco139625, w_eco139626, w_eco139627, w_eco139628, w_eco139629, w_eco139630, w_eco139631, w_eco139632, w_eco139633, w_eco139634, w_eco139635, w_eco139636, w_eco139637, w_eco139638, w_eco139639, w_eco139640, w_eco139641, w_eco139642, w_eco139643, w_eco139644, w_eco139645, w_eco139646, w_eco139647, w_eco139648, w_eco139649, w_eco139650, w_eco139651, w_eco139652, w_eco139653, w_eco139654, w_eco139655, w_eco139656, w_eco139657, w_eco139658, w_eco139659, w_eco139660, w_eco139661, w_eco139662, w_eco139663, w_eco139664, w_eco139665, w_eco139666, w_eco139667, w_eco139668, w_eco139669, w_eco139670, w_eco139671, w_eco139672, w_eco139673, w_eco139674, w_eco139675, w_eco139676, w_eco139677, w_eco139678, w_eco139679, w_eco139680, w_eco139681, w_eco139682, w_eco139683, w_eco139684, w_eco139685, w_eco139686, w_eco139687, w_eco139688, w_eco139689, w_eco139690, w_eco139691, w_eco139692, w_eco139693, w_eco139694, w_eco139695, w_eco139696, w_eco139697, w_eco139698, w_eco139699, w_eco139700, w_eco139701, w_eco139702, w_eco139703, w_eco139704, w_eco139705, w_eco139706, w_eco139707, w_eco139708, w_eco139709, w_eco139710, w_eco139711, w_eco139712, w_eco139713, w_eco139714, w_eco139715, w_eco139716, w_eco139717, w_eco139718, w_eco139719, w_eco139720, w_eco139721, w_eco139722, w_eco139723, w_eco139724, w_eco139725, w_eco139726, w_eco139727, w_eco139728, w_eco139729, w_eco139730, w_eco139731, w_eco139732, w_eco139733, w_eco139734, w_eco139735, w_eco139736, w_eco139737, w_eco139738, w_eco139739, w_eco139740, w_eco139741, w_eco139742, w_eco139743, w_eco139744, w_eco139745, w_eco139746, w_eco139747, w_eco139748, w_eco139749, w_eco139750, w_eco139751, w_eco139752, w_eco139753, w_eco139754, w_eco139755, w_eco139756, w_eco139757, w_eco139758, w_eco139759, w_eco139760, w_eco139761, w_eco139762, w_eco139763, w_eco139764, w_eco139765, w_eco139766, w_eco139767, w_eco139768, w_eco139769, w_eco139770, w_eco139771, w_eco139772, w_eco139773, w_eco139774, w_eco139775, w_eco139776, w_eco139777, w_eco139778, w_eco139779, w_eco139780, w_eco139781, w_eco139782, w_eco139783, w_eco139784, w_eco139785, w_eco139786, w_eco139787, w_eco139788, w_eco139789, w_eco139790, w_eco139791, w_eco139792, w_eco139793, w_eco139794, w_eco139795, w_eco139796, w_eco139797, w_eco139798, w_eco139799, w_eco139800, w_eco139801, w_eco139802, w_eco139803, w_eco139804, w_eco139805, w_eco139806, w_eco139807, w_eco139808, w_eco139809, w_eco139810, w_eco139811, w_eco139812, w_eco139813, w_eco139814, w_eco139815, w_eco139816, w_eco139817, w_eco139818, w_eco139819, w_eco139820, w_eco139821, w_eco139822, w_eco139823, w_eco139824, w_eco139825, w_eco139826, w_eco139827, w_eco139828, w_eco139829, w_eco139830, w_eco139831, w_eco139832, w_eco139833, w_eco139834, w_eco139835, w_eco139836, w_eco139837, w_eco139838, w_eco139839, w_eco139840, w_eco139841, w_eco139842, w_eco139843, w_eco139844, w_eco139845, w_eco139846, w_eco139847, w_eco139848, w_eco139849, w_eco139850, w_eco139851, w_eco139852, w_eco139853, w_eco139854, w_eco139855, w_eco139856, w_eco139857, w_eco139858, w_eco139859, w_eco139860, w_eco139861, w_eco139862, w_eco139863, w_eco139864, w_eco139865, w_eco139866, w_eco139867, w_eco139868, w_eco139869, w_eco139870, w_eco139871, w_eco139872, w_eco139873, w_eco139874, w_eco139875, w_eco139876, w_eco139877, w_eco139878, w_eco139879, w_eco139880, w_eco139881, w_eco139882, w_eco139883, w_eco139884, w_eco139885, w_eco139886, w_eco139887, w_eco139888, w_eco139889, w_eco139890, w_eco139891, w_eco139892, w_eco139893, w_eco139894, w_eco139895, w_eco139896, w_eco139897, w_eco139898, w_eco139899, w_eco139900, w_eco139901, w_eco139902, w_eco139903, w_eco139904, w_eco139905, w_eco139906, w_eco139907, w_eco139908, w_eco139909, w_eco139910, w_eco139911, w_eco139912, w_eco139913, w_eco139914, w_eco139915, w_eco139916, w_eco139917, w_eco139918, w_eco139919, w_eco139920, w_eco139921, w_eco139922, w_eco139923, w_eco139924, w_eco139925, w_eco139926, w_eco139927, w_eco139928, w_eco139929, w_eco139930, w_eco139931, w_eco139932, w_eco139933, w_eco139934, w_eco139935, w_eco139936, w_eco139937, w_eco139938, w_eco139939, w_eco139940, w_eco139941, w_eco139942, w_eco139943, w_eco139944, w_eco139945, w_eco139946, w_eco139947, w_eco139948, w_eco139949, w_eco139950, w_eco139951, w_eco139952, w_eco139953, w_eco139954, w_eco139955, w_eco139956, w_eco139957, w_eco139958, w_eco139959, w_eco139960, w_eco139961, w_eco139962, w_eco139963, w_eco139964, w_eco139965, w_eco139966, w_eco139967, w_eco139968, w_eco139969, w_eco139970, w_eco139971, w_eco139972, w_eco139973, w_eco139974, w_eco139975, w_eco139976, w_eco139977, w_eco139978, w_eco139979, w_eco139980, w_eco139981, w_eco139982, w_eco139983, w_eco139984, w_eco139985, w_eco139986, w_eco139987, w_eco139988, w_eco139989, w_eco139990, w_eco139991, w_eco139992, w_eco139993, w_eco139994, w_eco139995, w_eco139996, w_eco139997, w_eco139998, w_eco139999, w_eco140000, w_eco140001, w_eco140002, w_eco140003, w_eco140004, w_eco140005, w_eco140006, w_eco140007, w_eco140008, w_eco140009, w_eco140010, w_eco140011, w_eco140012, w_eco140013, w_eco140014, w_eco140015, w_eco140016, w_eco140017, w_eco140018, w_eco140019, w_eco140020, w_eco140021, w_eco140022, w_eco140023, w_eco140024, w_eco140025, w_eco140026, w_eco140027, w_eco140028, w_eco140029, w_eco140030, w_eco140031, w_eco140032, w_eco140033, w_eco140034, w_eco140035, w_eco140036, w_eco140037, w_eco140038, w_eco140039, w_eco140040, w_eco140041, w_eco140042, w_eco140043, w_eco140044, w_eco140045, w_eco140046, w_eco140047, w_eco140048, w_eco140049, w_eco140050, w_eco140051, w_eco140052, w_eco140053, w_eco140054, w_eco140055, w_eco140056, w_eco140057, w_eco140058, w_eco140059, w_eco140060, w_eco140061, w_eco140062, w_eco140063, w_eco140064, w_eco140065, w_eco140066, w_eco140067, w_eco140068, w_eco140069, w_eco140070, w_eco140071, w_eco140072, w_eco140073, w_eco140074, w_eco140075, w_eco140076, w_eco140077, w_eco140078, w_eco140079, w_eco140080, w_eco140081, w_eco140082, w_eco140083, w_eco140084, w_eco140085, w_eco140086, w_eco140087, w_eco140088, w_eco140089, w_eco140090, w_eco140091, w_eco140092, w_eco140093, w_eco140094, w_eco140095, w_eco140096, w_eco140097, w_eco140098, w_eco140099, w_eco140100, w_eco140101, w_eco140102, w_eco140103, w_eco140104, w_eco140105, w_eco140106, w_eco140107, w_eco140108, w_eco140109, w_eco140110, w_eco140111, w_eco140112, w_eco140113, w_eco140114, w_eco140115, w_eco140116, w_eco140117, w_eco140118, w_eco140119, w_eco140120, w_eco140121, w_eco140122, w_eco140123, w_eco140124, w_eco140125, w_eco140126, w_eco140127, w_eco140128, w_eco140129, w_eco140130, w_eco140131, w_eco140132, w_eco140133, w_eco140134, w_eco140135, w_eco140136, w_eco140137, w_eco140138, w_eco140139, w_eco140140, w_eco140141, w_eco140142, w_eco140143, w_eco140144, w_eco140145, w_eco140146, w_eco140147, w_eco140148, w_eco140149, w_eco140150, w_eco140151, w_eco140152, w_eco140153, w_eco140154, w_eco140155, w_eco140156, w_eco140157, w_eco140158, w_eco140159, w_eco140160, w_eco140161, w_eco140162, w_eco140163, w_eco140164, w_eco140165, w_eco140166, w_eco140167, w_eco140168, w_eco140169, w_eco140170, w_eco140171, w_eco140172, w_eco140173, w_eco140174, w_eco140175, w_eco140176, w_eco140177, w_eco140178, w_eco140179, w_eco140180, w_eco140181, w_eco140182, w_eco140183, w_eco140184, w_eco140185, w_eco140186, w_eco140187, w_eco140188, w_eco140189, w_eco140190, w_eco140191, w_eco140192, w_eco140193, w_eco140194, w_eco140195, w_eco140196, w_eco140197, w_eco140198, w_eco140199, w_eco140200, w_eco140201, w_eco140202, w_eco140203, w_eco140204, w_eco140205, w_eco140206, w_eco140207, w_eco140208, w_eco140209, w_eco140210, w_eco140211, w_eco140212, w_eco140213, w_eco140214, w_eco140215, w_eco140216, w_eco140217, w_eco140218, w_eco140219, w_eco140220, w_eco140221, w_eco140222, w_eco140223, w_eco140224, w_eco140225, w_eco140226, w_eco140227, w_eco140228, w_eco140229, w_eco140230, w_eco140231, w_eco140232, w_eco140233, w_eco140234, w_eco140235, w_eco140236, w_eco140237, w_eco140238, w_eco140239, w_eco140240, w_eco140241, w_eco140242, w_eco140243, w_eco140244, w_eco140245, w_eco140246, w_eco140247, w_eco140248, w_eco140249, w_eco140250, w_eco140251, w_eco140252, w_eco140253, w_eco140254, w_eco140255, w_eco140256, w_eco140257, w_eco140258, w_eco140259, w_eco140260, w_eco140261, w_eco140262, w_eco140263, w_eco140264, w_eco140265, w_eco140266, w_eco140267, w_eco140268, w_eco140269, w_eco140270, w_eco140271, w_eco140272, w_eco140273, w_eco140274, w_eco140275, w_eco140276, w_eco140277, w_eco140278, w_eco140279, w_eco140280, w_eco140281, w_eco140282, w_eco140283, w_eco140284, w_eco140285, w_eco140286, w_eco140287, w_eco140288, w_eco140289, w_eco140290, w_eco140291, w_eco140292, w_eco140293, w_eco140294, w_eco140295, w_eco140296, w_eco140297, w_eco140298, w_eco140299, w_eco140300, w_eco140301, w_eco140302, w_eco140303, w_eco140304, w_eco140305, w_eco140306, w_eco140307, w_eco140308, w_eco140309, w_eco140310, w_eco140311, w_eco140312, w_eco140313, w_eco140314, w_eco140315, w_eco140316, w_eco140317, w_eco140318, w_eco140319, w_eco140320, w_eco140321, w_eco140322, w_eco140323, w_eco140324, w_eco140325, w_eco140326, w_eco140327, w_eco140328, w_eco140329, w_eco140330, w_eco140331, w_eco140332, w_eco140333, w_eco140334, w_eco140335, w_eco140336, w_eco140337, w_eco140338, w_eco140339, w_eco140340, w_eco140341, w_eco140342, w_eco140343, w_eco140344, w_eco140345, w_eco140346, w_eco140347, w_eco140348, w_eco140349, w_eco140350, w_eco140351, w_eco140352, w_eco140353, w_eco140354, w_eco140355, w_eco140356, w_eco140357, w_eco140358, w_eco140359, w_eco140360, w_eco140361, w_eco140362, w_eco140363, w_eco140364, w_eco140365, w_eco140366, w_eco140367, w_eco140368, w_eco140369, w_eco140370, w_eco140371, w_eco140372, w_eco140373, w_eco140374, w_eco140375, w_eco140376, w_eco140377, w_eco140378, w_eco140379, w_eco140380, w_eco140381, w_eco140382, w_eco140383, w_eco140384, w_eco140385, w_eco140386, w_eco140387, w_eco140388, w_eco140389, w_eco140390, w_eco140391, w_eco140392, w_eco140393, w_eco140394, w_eco140395, w_eco140396, w_eco140397, w_eco140398, w_eco140399, w_eco140400, w_eco140401, w_eco140402, w_eco140403, w_eco140404, w_eco140405, w_eco140406, w_eco140407, w_eco140408, w_eco140409, w_eco140410, w_eco140411, w_eco140412, w_eco140413, w_eco140414, w_eco140415, w_eco140416, w_eco140417, w_eco140418, w_eco140419, w_eco140420, w_eco140421, w_eco140422, w_eco140423, w_eco140424, w_eco140425, w_eco140426, w_eco140427, w_eco140428, w_eco140429, w_eco140430, w_eco140431, w_eco140432, w_eco140433, w_eco140434, w_eco140435, w_eco140436, w_eco140437, w_eco140438, w_eco140439, w_eco140440, w_eco140441, w_eco140442, w_eco140443, w_eco140444, w_eco140445, w_eco140446, w_eco140447, w_eco140448, w_eco140449, w_eco140450, w_eco140451, w_eco140452, w_eco140453, w_eco140454, w_eco140455, w_eco140456, w_eco140457, w_eco140458, w_eco140459, w_eco140460, w_eco140461, w_eco140462, w_eco140463, w_eco140464, w_eco140465, w_eco140466, w_eco140467, w_eco140468, w_eco140469, w_eco140470, w_eco140471, w_eco140472, w_eco140473, w_eco140474, w_eco140475, w_eco140476, w_eco140477, w_eco140478, w_eco140479, w_eco140480, w_eco140481, w_eco140482, w_eco140483, w_eco140484, w_eco140485, w_eco140486, w_eco140487, w_eco140488, w_eco140489, w_eco140490, w_eco140491, w_eco140492, w_eco140493, w_eco140494, w_eco140495, w_eco140496, w_eco140497, w_eco140498, w_eco140499, w_eco140500, w_eco140501, w_eco140502, w_eco140503, w_eco140504, w_eco140505, w_eco140506, w_eco140507, w_eco140508, w_eco140509, w_eco140510, w_eco140511, w_eco140512, w_eco140513, w_eco140514, w_eco140515, w_eco140516, w_eco140517, w_eco140518, w_eco140519, w_eco140520, w_eco140521, w_eco140522, w_eco140523, w_eco140524, w_eco140525, w_eco140526, w_eco140527, w_eco140528, w_eco140529, w_eco140530, w_eco140531, w_eco140532, w_eco140533, w_eco140534, w_eco140535, w_eco140536, w_eco140537, w_eco140538, w_eco140539, w_eco140540, w_eco140541, w_eco140542, w_eco140543, w_eco140544, w_eco140545, w_eco140546, w_eco140547, w_eco140548, w_eco140549, w_eco140550, w_eco140551, w_eco140552, w_eco140553, w_eco140554, w_eco140555, w_eco140556, w_eco140557, w_eco140558, w_eco140559, w_eco140560, w_eco140561, w_eco140562, w_eco140563, w_eco140564, w_eco140565, w_eco140566, w_eco140567, w_eco140568, w_eco140569, w_eco140570, w_eco140571, w_eco140572, w_eco140573, w_eco140574, w_eco140575, w_eco140576, w_eco140577, w_eco140578, w_eco140579, w_eco140580, w_eco140581, w_eco140582, w_eco140583, w_eco140584, w_eco140585, w_eco140586, w_eco140587, w_eco140588, w_eco140589, w_eco140590, w_eco140591, w_eco140592, w_eco140593, w_eco140594, w_eco140595, w_eco140596, w_eco140597, w_eco140598, w_eco140599, w_eco140600, w_eco140601, w_eco140602, w_eco140603, w_eco140604, w_eco140605, w_eco140606, w_eco140607, w_eco140608, w_eco140609, w_eco140610, w_eco140611, w_eco140612, w_eco140613, w_eco140614, w_eco140615, w_eco140616, w_eco140617, w_eco140618, w_eco140619, w_eco140620, w_eco140621, w_eco140622, w_eco140623, w_eco140624, w_eco140625, w_eco140626, w_eco140627, w_eco140628, w_eco140629, w_eco140630, w_eco140631, w_eco140632, w_eco140633, w_eco140634, w_eco140635, w_eco140636, w_eco140637, w_eco140638, w_eco140639, w_eco140640, w_eco140641, w_eco140642, w_eco140643, w_eco140644, w_eco140645, w_eco140646, w_eco140647, w_eco140648, w_eco140649, w_eco140650, w_eco140651, w_eco140652, w_eco140653, w_eco140654, w_eco140655, w_eco140656, w_eco140657, w_eco140658, w_eco140659, w_eco140660, w_eco140661, w_eco140662, w_eco140663, w_eco140664, w_eco140665, w_eco140666, w_eco140667, w_eco140668, w_eco140669, w_eco140670, w_eco140671, w_eco140672, w_eco140673, w_eco140674, w_eco140675, w_eco140676, w_eco140677, w_eco140678, w_eco140679, w_eco140680, w_eco140681, w_eco140682, w_eco140683, w_eco140684, w_eco140685, w_eco140686, w_eco140687, w_eco140688, w_eco140689, w_eco140690, w_eco140691, w_eco140692, w_eco140693, w_eco140694, w_eco140695, w_eco140696, w_eco140697, w_eco140698, w_eco140699, w_eco140700, w_eco140701, w_eco140702, w_eco140703, w_eco140704, w_eco140705, w_eco140706, w_eco140707, w_eco140708, w_eco140709, w_eco140710, w_eco140711, w_eco140712, w_eco140713, w_eco140714, w_eco140715, w_eco140716, w_eco140717, w_eco140718, w_eco140719, w_eco140720, w_eco140721, w_eco140722, w_eco140723, w_eco140724, w_eco140725, w_eco140726, w_eco140727, w_eco140728, w_eco140729, w_eco140730, w_eco140731, w_eco140732, w_eco140733, w_eco140734, w_eco140735, w_eco140736, w_eco140737, w_eco140738, w_eco140739, w_eco140740, w_eco140741, w_eco140742, w_eco140743, w_eco140744, w_eco140745, w_eco140746, w_eco140747, w_eco140748, w_eco140749, w_eco140750, w_eco140751, w_eco140752, w_eco140753, w_eco140754, w_eco140755, w_eco140756, w_eco140757, w_eco140758, w_eco140759, w_eco140760, w_eco140761, w_eco140762, w_eco140763, w_eco140764, w_eco140765, w_eco140766, w_eco140767, w_eco140768, w_eco140769, w_eco140770, w_eco140771, w_eco140772, w_eco140773, w_eco140774, w_eco140775, w_eco140776, w_eco140777, w_eco140778, w_eco140779, w_eco140780, w_eco140781, w_eco140782, w_eco140783, w_eco140784, w_eco140785, w_eco140786, w_eco140787, w_eco140788, w_eco140789, w_eco140790, w_eco140791, w_eco140792, w_eco140793, w_eco140794, w_eco140795, w_eco140796, w_eco140797, w_eco140798, w_eco140799, w_eco140800, w_eco140801, w_eco140802, w_eco140803, w_eco140804, w_eco140805, w_eco140806, w_eco140807, w_eco140808, w_eco140809, w_eco140810, w_eco140811, w_eco140812, w_eco140813, w_eco140814, w_eco140815, w_eco140816, w_eco140817, w_eco140818, w_eco140819, w_eco140820, w_eco140821, w_eco140822, w_eco140823, w_eco140824, w_eco140825, w_eco140826, w_eco140827, w_eco140828, w_eco140829, w_eco140830, w_eco140831, w_eco140832, w_eco140833, w_eco140834, w_eco140835, w_eco140836, w_eco140837, w_eco140838, w_eco140839, w_eco140840, w_eco140841, w_eco140842, w_eco140843, w_eco140844, w_eco140845, w_eco140846, w_eco140847, w_eco140848, w_eco140849, w_eco140850, w_eco140851, w_eco140852, w_eco140853, w_eco140854, w_eco140855, w_eco140856, w_eco140857, w_eco140858, w_eco140859, w_eco140860, w_eco140861, w_eco140862, w_eco140863, w_eco140864, w_eco140865, w_eco140866, w_eco140867, w_eco140868, w_eco140869, w_eco140870, w_eco140871, w_eco140872, w_eco140873, w_eco140874, w_eco140875, w_eco140876, w_eco140877, w_eco140878, w_eco140879, w_eco140880, w_eco140881, w_eco140882, w_eco140883, w_eco140884, w_eco140885, w_eco140886, w_eco140887, w_eco140888, w_eco140889, w_eco140890, w_eco140891, w_eco140892, w_eco140893, w_eco140894, w_eco140895, w_eco140896, w_eco140897, w_eco140898, w_eco140899, w_eco140900, w_eco140901, w_eco140902, w_eco140903, w_eco140904, w_eco140905, w_eco140906, w_eco140907, w_eco140908, w_eco140909, w_eco140910, w_eco140911, w_eco140912, w_eco140913, w_eco140914, w_eco140915, w_eco140916, w_eco140917, w_eco140918, w_eco140919, w_eco140920, w_eco140921, w_eco140922, w_eco140923, w_eco140924, w_eco140925, w_eco140926, w_eco140927, w_eco140928, w_eco140929, w_eco140930, w_eco140931, w_eco140932, w_eco140933, w_eco140934, w_eco140935, w_eco140936, w_eco140937, w_eco140938, w_eco140939, w_eco140940, w_eco140941, w_eco140942, w_eco140943, w_eco140944, w_eco140945, w_eco140946, w_eco140947, w_eco140948, w_eco140949, w_eco140950, w_eco140951, w_eco140952, w_eco140953, w_eco140954, w_eco140955, w_eco140956, w_eco140957, w_eco140958, w_eco140959, w_eco140960, w_eco140961, w_eco140962, w_eco140963, w_eco140964, w_eco140965, w_eco140966, w_eco140967, w_eco140968, w_eco140969, w_eco140970, w_eco140971, w_eco140972, w_eco140973, w_eco140974, w_eco140975, w_eco140976, w_eco140977, w_eco140978, w_eco140979, w_eco140980, w_eco140981, w_eco140982, w_eco140983, w_eco140984, w_eco140985, w_eco140986, w_eco140987, w_eco140988, w_eco140989, w_eco140990, w_eco140991, w_eco140992, w_eco140993, w_eco140994, w_eco140995, w_eco140996, w_eco140997, w_eco140998, w_eco140999, w_eco141000, w_eco141001, w_eco141002, w_eco141003, w_eco141004, w_eco141005, w_eco141006, w_eco141007, w_eco141008, w_eco141009, w_eco141010, w_eco141011, w_eco141012, w_eco141013, w_eco141014, w_eco141015, w_eco141016, w_eco141017, w_eco141018, w_eco141019, w_eco141020, w_eco141021, w_eco141022, w_eco141023, w_eco141024, w_eco141025, w_eco141026, w_eco141027, w_eco141028, w_eco141029, w_eco141030, w_eco141031, w_eco141032, w_eco141033, w_eco141034, w_eco141035, w_eco141036, w_eco141037, w_eco141038, w_eco141039, w_eco141040, w_eco141041, w_eco141042, w_eco141043, w_eco141044, w_eco141045, w_eco141046, w_eco141047, w_eco141048, w_eco141049, w_eco141050, w_eco141051, w_eco141052, w_eco141053, w_eco141054, w_eco141055, w_eco141056, w_eco141057, w_eco141058, w_eco141059, w_eco141060, w_eco141061, w_eco141062, w_eco141063, w_eco141064, w_eco141065, w_eco141066, w_eco141067, w_eco141068, w_eco141069, w_eco141070, w_eco141071, w_eco141072, w_eco141073, w_eco141074, w_eco141075, w_eco141076, w_eco141077, w_eco141078, w_eco141079, w_eco141080, w_eco141081, w_eco141082, w_eco141083, w_eco141084, w_eco141085, w_eco141086, w_eco141087, w_eco141088, w_eco141089, w_eco141090, w_eco141091, w_eco141092, w_eco141093, w_eco141094, w_eco141095, w_eco141096, w_eco141097, w_eco141098, w_eco141099, w_eco141100, w_eco141101, w_eco141102, w_eco141103, w_eco141104, w_eco141105, w_eco141106, w_eco141107, w_eco141108, w_eco141109, w_eco141110, w_eco141111, w_eco141112, w_eco141113, w_eco141114, w_eco141115, w_eco141116, w_eco141117, w_eco141118, w_eco141119, w_eco141120, w_eco141121, w_eco141122, w_eco141123, w_eco141124, w_eco141125, w_eco141126, w_eco141127, w_eco141128, w_eco141129, w_eco141130, w_eco141131, w_eco141132, w_eco141133, w_eco141134, w_eco141135, w_eco141136, w_eco141137, w_eco141138, w_eco141139, w_eco141140, w_eco141141, w_eco141142, w_eco141143, w_eco141144, w_eco141145, w_eco141146, w_eco141147, w_eco141148, w_eco141149, w_eco141150, w_eco141151, w_eco141152, w_eco141153, w_eco141154, w_eco141155, w_eco141156, w_eco141157, w_eco141158, w_eco141159, w_eco141160, w_eco141161, w_eco141162, w_eco141163, w_eco141164, w_eco141165, w_eco141166, w_eco141167, w_eco141168, w_eco141169, w_eco141170, w_eco141171, w_eco141172, w_eco141173, w_eco141174, w_eco141175, w_eco141176, w_eco141177, w_eco141178, w_eco141179, w_eco141180, w_eco141181, w_eco141182, w_eco141183, w_eco141184, w_eco141185, w_eco141186, w_eco141187, w_eco141188, w_eco141189, w_eco141190, w_eco141191, w_eco141192, w_eco141193, w_eco141194, w_eco141195, w_eco141196, w_eco141197, w_eco141198, w_eco141199, w_eco141200, w_eco141201, w_eco141202, w_eco141203, w_eco141204, w_eco141205, w_eco141206, w_eco141207, w_eco141208, w_eco141209, w_eco141210, w_eco141211, w_eco141212, w_eco141213, w_eco141214, w_eco141215, w_eco141216, w_eco141217, w_eco141218, w_eco141219, w_eco141220, w_eco141221, w_eco141222, w_eco141223, w_eco141224, w_eco141225, w_eco141226, w_eco141227, w_eco141228, w_eco141229, w_eco141230, w_eco141231, w_eco141232, w_eco141233, w_eco141234, w_eco141235, w_eco141236, w_eco141237, w_eco141238, w_eco141239, w_eco141240, w_eco141241, w_eco141242, w_eco141243, w_eco141244, w_eco141245, w_eco141246, w_eco141247, w_eco141248, w_eco141249, w_eco141250, w_eco141251, w_eco141252, w_eco141253, w_eco141254, w_eco141255, w_eco141256, w_eco141257, w_eco141258, w_eco141259, w_eco141260, w_eco141261, w_eco141262, w_eco141263, w_eco141264, w_eco141265, w_eco141266, w_eco141267, w_eco141268, w_eco141269, w_eco141270, w_eco141271, w_eco141272, w_eco141273, w_eco141274, w_eco141275, w_eco141276, w_eco141277, w_eco141278, w_eco141279, w_eco141280, w_eco141281, w_eco141282, w_eco141283, w_eco141284, w_eco141285, w_eco141286, w_eco141287, w_eco141288, w_eco141289, w_eco141290, w_eco141291, w_eco141292, w_eco141293, w_eco141294, w_eco141295, w_eco141296, w_eco141297, w_eco141298, w_eco141299, w_eco141300, w_eco141301, w_eco141302, w_eco141303, w_eco141304, w_eco141305, w_eco141306, w_eco141307, w_eco141308, w_eco141309, w_eco141310, w_eco141311, w_eco141312, w_eco141313, w_eco141314, w_eco141315, w_eco141316, w_eco141317, w_eco141318, w_eco141319, w_eco141320, w_eco141321, w_eco141322, w_eco141323, w_eco141324, w_eco141325, w_eco141326, w_eco141327, w_eco141328, w_eco141329, w_eco141330, w_eco141331, w_eco141332, w_eco141333, w_eco141334, w_eco141335, w_eco141336, w_eco141337, w_eco141338, w_eco141339, w_eco141340, w_eco141341, w_eco141342, w_eco141343, w_eco141344, w_eco141345, w_eco141346, w_eco141347, w_eco141348, w_eco141349, w_eco141350, w_eco141351, w_eco141352, w_eco141353, w_eco141354, w_eco141355, w_eco141356, w_eco141357, w_eco141358, w_eco141359, w_eco141360, w_eco141361, w_eco141362, w_eco141363, w_eco141364, w_eco141365, w_eco141366, w_eco141367, w_eco141368, w_eco141369, w_eco141370, w_eco141371, w_eco141372, w_eco141373, w_eco141374, w_eco141375, w_eco141376, w_eco141377, w_eco141378, w_eco141379, w_eco141380, w_eco141381, w_eco141382, w_eco141383, w_eco141384, w_eco141385, w_eco141386, w_eco141387, w_eco141388, w_eco141389, w_eco141390, w_eco141391, w_eco141392, w_eco141393, w_eco141394, w_eco141395, w_eco141396, w_eco141397, w_eco141398, w_eco141399, w_eco141400, w_eco141401, w_eco141402, w_eco141403, w_eco141404, w_eco141405, w_eco141406, w_eco141407, w_eco141408, w_eco141409, w_eco141410, w_eco141411, w_eco141412, w_eco141413, w_eco141414, w_eco141415, w_eco141416, w_eco141417, w_eco141418, w_eco141419, w_eco141420, w_eco141421, w_eco141422, w_eco141423, w_eco141424, w_eco141425, w_eco141426, w_eco141427, w_eco141428, w_eco141429, w_eco141430, w_eco141431, w_eco141432, w_eco141433, w_eco141434, w_eco141435, w_eco141436, w_eco141437, w_eco141438, w_eco141439, w_eco141440, w_eco141441, w_eco141442, w_eco141443, w_eco141444, w_eco141445, w_eco141446, w_eco141447, w_eco141448, w_eco141449, w_eco141450, w_eco141451, w_eco141452, w_eco141453, w_eco141454, w_eco141455, w_eco141456, w_eco141457, w_eco141458, w_eco141459, w_eco141460, w_eco141461, w_eco141462, w_eco141463, w_eco141464, w_eco141465, w_eco141466, w_eco141467, w_eco141468, w_eco141469, w_eco141470, w_eco141471, w_eco141472, w_eco141473, w_eco141474, w_eco141475, w_eco141476, w_eco141477, w_eco141478, w_eco141479, w_eco141480, w_eco141481, w_eco141482, w_eco141483, w_eco141484, w_eco141485, w_eco141486, w_eco141487, w_eco141488, w_eco141489, w_eco141490, w_eco141491, w_eco141492, w_eco141493, w_eco141494, w_eco141495, w_eco141496, w_eco141497, w_eco141498, w_eco141499, w_eco141500, w_eco141501, w_eco141502, w_eco141503, w_eco141504, w_eco141505, w_eco141506, w_eco141507, w_eco141508, w_eco141509, w_eco141510, w_eco141511, w_eco141512, w_eco141513, w_eco141514, w_eco141515, w_eco141516, w_eco141517, w_eco141518, w_eco141519, w_eco141520, w_eco141521, w_eco141522, w_eco141523, w_eco141524, w_eco141525, w_eco141526, w_eco141527, w_eco141528, w_eco141529, w_eco141530, w_eco141531, w_eco141532, w_eco141533, w_eco141534, w_eco141535, w_eco141536, w_eco141537, w_eco141538, w_eco141539, w_eco141540, w_eco141541, w_eco141542, w_eco141543, w_eco141544, w_eco141545, w_eco141546, w_eco141547, w_eco141548, w_eco141549, w_eco141550, w_eco141551, w_eco141552, w_eco141553, w_eco141554, w_eco141555, w_eco141556, w_eco141557, w_eco141558, w_eco141559, w_eco141560, w_eco141561, w_eco141562, w_eco141563, w_eco141564, w_eco141565, w_eco141566, w_eco141567, w_eco141568, w_eco141569, w_eco141570, w_eco141571, w_eco141572, w_eco141573, w_eco141574, w_eco141575, w_eco141576, w_eco141577, w_eco141578, w_eco141579, w_eco141580, w_eco141581, w_eco141582, w_eco141583, w_eco141584, w_eco141585, w_eco141586, w_eco141587, w_eco141588, w_eco141589, w_eco141590, w_eco141591, w_eco141592, w_eco141593, w_eco141594, w_eco141595, w_eco141596, w_eco141597, w_eco141598, w_eco141599, w_eco141600, w_eco141601, w_eco141602, w_eco141603, w_eco141604, w_eco141605, w_eco141606, w_eco141607, w_eco141608, w_eco141609, w_eco141610, w_eco141611, w_eco141612, w_eco141613, w_eco141614, w_eco141615, w_eco141616, w_eco141617, w_eco141618, w_eco141619, w_eco141620, w_eco141621, w_eco141622, w_eco141623, w_eco141624, w_eco141625, w_eco141626, w_eco141627, w_eco141628, w_eco141629, w_eco141630, w_eco141631, w_eco141632, w_eco141633, w_eco141634, w_eco141635, w_eco141636, w_eco141637, w_eco141638, w_eco141639, w_eco141640, w_eco141641, w_eco141642, w_eco141643, w_eco141644, w_eco141645, w_eco141646, w_eco141647, w_eco141648, w_eco141649, w_eco141650, w_eco141651, w_eco141652, w_eco141653, w_eco141654, w_eco141655, w_eco141656, w_eco141657, w_eco141658, w_eco141659, w_eco141660, w_eco141661, w_eco141662, w_eco141663, w_eco141664, w_eco141665, w_eco141666, w_eco141667, w_eco141668, w_eco141669, w_eco141670, w_eco141671, w_eco141672, w_eco141673, w_eco141674, w_eco141675, w_eco141676, w_eco141677, w_eco141678, w_eco141679, w_eco141680, w_eco141681, w_eco141682, w_eco141683, w_eco141684, w_eco141685, w_eco141686, w_eco141687, w_eco141688, w_eco141689, w_eco141690, w_eco141691, w_eco141692, w_eco141693, w_eco141694, w_eco141695, w_eco141696, w_eco141697, w_eco141698, w_eco141699, w_eco141700, w_eco141701, w_eco141702, w_eco141703, w_eco141704, w_eco141705, w_eco141706, w_eco141707, w_eco141708, w_eco141709, w_eco141710, w_eco141711, w_eco141712, w_eco141713, w_eco141714, w_eco141715, w_eco141716, w_eco141717, w_eco141718, w_eco141719, w_eco141720, w_eco141721, w_eco141722, w_eco141723, w_eco141724, w_eco141725, w_eco141726, w_eco141727, w_eco141728, w_eco141729, w_eco141730, w_eco141731, w_eco141732, w_eco141733, w_eco141734, w_eco141735, w_eco141736, w_eco141737, w_eco141738, w_eco141739, w_eco141740, w_eco141741, w_eco141742, w_eco141743, w_eco141744, w_eco141745, w_eco141746, w_eco141747, w_eco141748, w_eco141749, w_eco141750, w_eco141751, w_eco141752, w_eco141753, w_eco141754, w_eco141755, w_eco141756, w_eco141757, w_eco141758, w_eco141759, w_eco141760, w_eco141761, w_eco141762, w_eco141763, w_eco141764, w_eco141765, w_eco141766, w_eco141767, w_eco141768, w_eco141769, w_eco141770, w_eco141771, w_eco141772, w_eco141773, w_eco141774, w_eco141775, w_eco141776, w_eco141777, w_eco141778, w_eco141779, w_eco141780, w_eco141781, w_eco141782, w_eco141783, w_eco141784, w_eco141785, w_eco141786, w_eco141787, w_eco141788, w_eco141789, w_eco141790, w_eco141791, w_eco141792, w_eco141793, w_eco141794, w_eco141795, w_eco141796, w_eco141797, w_eco141798, w_eco141799, w_eco141800, w_eco141801, w_eco141802, w_eco141803, w_eco141804, w_eco141805, w_eco141806, w_eco141807, w_eco141808, w_eco141809, w_eco141810, w_eco141811, w_eco141812, w_eco141813, w_eco141814, w_eco141815, w_eco141816, w_eco141817, w_eco141818, w_eco141819, w_eco141820, w_eco141821, w_eco141822, w_eco141823, w_eco141824, w_eco141825, w_eco141826, w_eco141827, w_eco141828, w_eco141829, w_eco141830, w_eco141831, w_eco141832, w_eco141833, w_eco141834, w_eco141835, w_eco141836, w_eco141837, w_eco141838, w_eco141839, w_eco141840, w_eco141841, w_eco141842, w_eco141843, w_eco141844, w_eco141845, w_eco141846, w_eco141847, w_eco141848, w_eco141849, w_eco141850, w_eco141851, w_eco141852, w_eco141853, w_eco141854, w_eco141855, w_eco141856, w_eco141857, w_eco141858, w_eco141859, w_eco141860, w_eco141861, w_eco141862, w_eco141863, w_eco141864, w_eco141865, w_eco141866, w_eco141867, w_eco141868, w_eco141869, w_eco141870, w_eco141871, w_eco141872, w_eco141873, w_eco141874, w_eco141875, w_eco141876, w_eco141877, w_eco141878, w_eco141879, w_eco141880, w_eco141881, w_eco141882, w_eco141883, w_eco141884, w_eco141885, w_eco141886, w_eco141887, w_eco141888, w_eco141889, w_eco141890, w_eco141891, w_eco141892, w_eco141893, w_eco141894, w_eco141895, w_eco141896, w_eco141897, w_eco141898, w_eco141899, w_eco141900, w_eco141901, w_eco141902, w_eco141903, w_eco141904, w_eco141905, w_eco141906, w_eco141907, w_eco141908, w_eco141909, w_eco141910, w_eco141911, w_eco141912, w_eco141913, w_eco141914, w_eco141915, w_eco141916, w_eco141917, w_eco141918, w_eco141919, w_eco141920, w_eco141921, w_eco141922, w_eco141923, w_eco141924, w_eco141925, w_eco141926, w_eco141927, w_eco141928, w_eco141929, w_eco141930, w_eco141931, w_eco141932, w_eco141933, w_eco141934, w_eco141935, w_eco141936, w_eco141937, w_eco141938, w_eco141939, w_eco141940, w_eco141941, w_eco141942, w_eco141943, w_eco141944, w_eco141945, w_eco141946, w_eco141947, w_eco141948, w_eco141949, w_eco141950, w_eco141951, w_eco141952, w_eco141953, w_eco141954, w_eco141955, w_eco141956, w_eco141957, w_eco141958, w_eco141959, w_eco141960, w_eco141961, w_eco141962, w_eco141963, w_eco141964, w_eco141965, w_eco141966, w_eco141967, w_eco141968, w_eco141969, w_eco141970, w_eco141971, w_eco141972, w_eco141973, w_eco141974, w_eco141975, w_eco141976, w_eco141977, w_eco141978, w_eco141979, w_eco141980, w_eco141981, w_eco141982, w_eco141983, w_eco141984, w_eco141985, w_eco141986, w_eco141987, w_eco141988, w_eco141989, w_eco141990, w_eco141991, w_eco141992, w_eco141993, w_eco141994, w_eco141995, w_eco141996, w_eco141997, w_eco141998, w_eco141999, w_eco142000, w_eco142001, w_eco142002, w_eco142003, w_eco142004, w_eco142005, w_eco142006, w_eco142007, w_eco142008, w_eco142009, w_eco142010, w_eco142011, w_eco142012, w_eco142013, w_eco142014, w_eco142015, w_eco142016, w_eco142017, w_eco142018, w_eco142019, w_eco142020, w_eco142021, w_eco142022, w_eco142023, w_eco142024, w_eco142025, w_eco142026, w_eco142027, w_eco142028, w_eco142029, w_eco142030, w_eco142031, w_eco142032, w_eco142033, w_eco142034, w_eco142035, w_eco142036, w_eco142037, w_eco142038, w_eco142039, w_eco142040, w_eco142041, w_eco142042, w_eco142043, w_eco142044, w_eco142045, w_eco142046, w_eco142047, w_eco142048, w_eco142049, w_eco142050, w_eco142051, w_eco142052, w_eco142053, w_eco142054, w_eco142055, w_eco142056, w_eco142057, w_eco142058, w_eco142059, w_eco142060, w_eco142061, w_eco142062, w_eco142063, w_eco142064, w_eco142065, w_eco142066, w_eco142067, w_eco142068, w_eco142069, w_eco142070, w_eco142071, w_eco142072, w_eco142073, w_eco142074, w_eco142075, w_eco142076, w_eco142077, w_eco142078, w_eco142079, w_eco142080, w_eco142081, w_eco142082, w_eco142083, w_eco142084, w_eco142085, w_eco142086, w_eco142087, w_eco142088, w_eco142089, w_eco142090, w_eco142091, w_eco142092, w_eco142093, w_eco142094, w_eco142095, w_eco142096, w_eco142097, w_eco142098, w_eco142099, w_eco142100, w_eco142101, w_eco142102, w_eco142103, w_eco142104, w_eco142105, w_eco142106, w_eco142107, w_eco142108, w_eco142109, w_eco142110, w_eco142111, w_eco142112, w_eco142113, w_eco142114, w_eco142115, w_eco142116, w_eco142117, w_eco142118, w_eco142119, w_eco142120, w_eco142121, w_eco142122, w_eco142123, w_eco142124, w_eco142125, w_eco142126, w_eco142127, w_eco142128, w_eco142129, w_eco142130, w_eco142131, w_eco142132, w_eco142133, w_eco142134, w_eco142135, w_eco142136, w_eco142137, w_eco142138, w_eco142139, w_eco142140, w_eco142141, w_eco142142, w_eco142143, w_eco142144, w_eco142145, w_eco142146, w_eco142147, w_eco142148, w_eco142149, w_eco142150, w_eco142151, w_eco142152, w_eco142153, w_eco142154, w_eco142155, w_eco142156, w_eco142157, w_eco142158, w_eco142159, w_eco142160, w_eco142161, w_eco142162, w_eco142163, w_eco142164, w_eco142165, w_eco142166, w_eco142167, w_eco142168, w_eco142169, w_eco142170, w_eco142171, w_eco142172, w_eco142173, w_eco142174, w_eco142175, w_eco142176, w_eco142177, w_eco142178, w_eco142179, w_eco142180, w_eco142181, w_eco142182, w_eco142183, w_eco142184, w_eco142185, w_eco142186, w_eco142187, w_eco142188, w_eco142189, w_eco142190, w_eco142191, w_eco142192, w_eco142193, w_eco142194, w_eco142195, w_eco142196, w_eco142197, w_eco142198, w_eco142199, w_eco142200, w_eco142201, w_eco142202, w_eco142203, w_eco142204, w_eco142205, w_eco142206, w_eco142207, w_eco142208, w_eco142209, w_eco142210, w_eco142211, w_eco142212, w_eco142213, w_eco142214, w_eco142215, w_eco142216, w_eco142217, w_eco142218, w_eco142219, w_eco142220, w_eco142221, w_eco142222, w_eco142223, w_eco142224, w_eco142225, w_eco142226, w_eco142227, w_eco142228, w_eco142229, w_eco142230, w_eco142231, w_eco142232, w_eco142233, w_eco142234, w_eco142235, w_eco142236, w_eco142237, w_eco142238, w_eco142239, w_eco142240, w_eco142241, w_eco142242, w_eco142243, w_eco142244, w_eco142245, w_eco142246, w_eco142247, w_eco142248, w_eco142249, w_eco142250, w_eco142251, w_eco142252, w_eco142253, w_eco142254, w_eco142255, w_eco142256, w_eco142257, w_eco142258, w_eco142259, w_eco142260, w_eco142261, w_eco142262, w_eco142263, w_eco142264, w_eco142265, w_eco142266, w_eco142267, w_eco142268, w_eco142269, w_eco142270, w_eco142271, w_eco142272, w_eco142273, w_eco142274, w_eco142275, w_eco142276, w_eco142277, w_eco142278, w_eco142279, w_eco142280, w_eco142281, w_eco142282, w_eco142283, w_eco142284, w_eco142285, w_eco142286, w_eco142287, w_eco142288, w_eco142289, w_eco142290, w_eco142291, w_eco142292, w_eco142293, w_eco142294, w_eco142295, w_eco142296, w_eco142297, w_eco142298, w_eco142299, w_eco142300, w_eco142301, w_eco142302, w_eco142303, w_eco142304, w_eco142305, w_eco142306, w_eco142307, w_eco142308, w_eco142309, w_eco142310, w_eco142311, w_eco142312, w_eco142313, w_eco142314, w_eco142315, w_eco142316, w_eco142317, w_eco142318, w_eco142319, w_eco142320, w_eco142321, w_eco142322, w_eco142323, w_eco142324, w_eco142325, w_eco142326, w_eco142327, w_eco142328, w_eco142329, w_eco142330, w_eco142331, w_eco142332, w_eco142333, w_eco142334, w_eco142335, w_eco142336, w_eco142337, w_eco142338, w_eco142339, w_eco142340, w_eco142341, w_eco142342, w_eco142343, w_eco142344, w_eco142345, w_eco142346, w_eco142347, w_eco142348, w_eco142349, w_eco142350, w_eco142351, w_eco142352, w_eco142353, w_eco142354, w_eco142355, w_eco142356, w_eco142357, w_eco142358, w_eco142359, w_eco142360, w_eco142361, w_eco142362, w_eco142363, w_eco142364, w_eco142365, w_eco142366, w_eco142367, w_eco142368, w_eco142369, w_eco142370, w_eco142371, w_eco142372, w_eco142373, w_eco142374, w_eco142375, w_eco142376, w_eco142377, w_eco142378, w_eco142379, w_eco142380, w_eco142381, w_eco142382, w_eco142383, w_eco142384, w_eco142385, w_eco142386, w_eco142387, w_eco142388, w_eco142389, w_eco142390, w_eco142391, w_eco142392, w_eco142393, w_eco142394, w_eco142395, w_eco142396, w_eco142397, w_eco142398, w_eco142399, w_eco142400, w_eco142401, w_eco142402, w_eco142403, w_eco142404, w_eco142405, w_eco142406, w_eco142407, w_eco142408, w_eco142409, w_eco142410, w_eco142411, w_eco142412, w_eco142413, w_eco142414, w_eco142415, w_eco142416, w_eco142417, w_eco142418, w_eco142419, w_eco142420, w_eco142421, w_eco142422, w_eco142423, w_eco142424, w_eco142425, w_eco142426, w_eco142427, w_eco142428, w_eco142429, w_eco142430, w_eco142431, w_eco142432, w_eco142433, w_eco142434, w_eco142435, w_eco142436, w_eco142437, w_eco142438, w_eco142439, w_eco142440, w_eco142441, w_eco142442, w_eco142443, w_eco142444, w_eco142445, w_eco142446, w_eco142447, w_eco142448, w_eco142449, w_eco142450, w_eco142451, w_eco142452, w_eco142453, w_eco142454, w_eco142455, w_eco142456, w_eco142457, w_eco142458, w_eco142459, w_eco142460, w_eco142461, w_eco142462, w_eco142463, w_eco142464, w_eco142465, w_eco142466, w_eco142467, w_eco142468, w_eco142469, w_eco142470, w_eco142471, w_eco142472, w_eco142473, w_eco142474, w_eco142475, w_eco142476, w_eco142477, w_eco142478, w_eco142479, w_eco142480, w_eco142481, w_eco142482, w_eco142483, w_eco142484, w_eco142485, w_eco142486, w_eco142487, w_eco142488, w_eco142489, w_eco142490, w_eco142491, w_eco142492, w_eco142493, w_eco142494, w_eco142495, w_eco142496, w_eco142497, w_eco142498, w_eco142499, w_eco142500, w_eco142501, w_eco142502, w_eco142503, w_eco142504, w_eco142505, w_eco142506, w_eco142507, w_eco142508, w_eco142509, w_eco142510, w_eco142511, w_eco142512, w_eco142513, w_eco142514, w_eco142515, w_eco142516, w_eco142517, w_eco142518, w_eco142519, w_eco142520, w_eco142521, w_eco142522, w_eco142523, w_eco142524, w_eco142525, w_eco142526, w_eco142527, w_eco142528, w_eco142529, w_eco142530, w_eco142531, w_eco142532, w_eco142533, w_eco142534, w_eco142535, w_eco142536, w_eco142537, w_eco142538, w_eco142539, w_eco142540, w_eco142541, w_eco142542, w_eco142543, w_eco142544, w_eco142545, w_eco142546, w_eco142547, w_eco142548, w_eco142549, w_eco142550, w_eco142551, w_eco142552, w_eco142553, w_eco142554, w_eco142555, w_eco142556, w_eco142557, w_eco142558, w_eco142559, w_eco142560, w_eco142561, w_eco142562, w_eco142563, w_eco142564, w_eco142565, w_eco142566, w_eco142567, w_eco142568, w_eco142569, w_eco142570, w_eco142571, w_eco142572, w_eco142573, w_eco142574, w_eco142575, w_eco142576, w_eco142577, w_eco142578, w_eco142579, w_eco142580, w_eco142581, w_eco142582, w_eco142583, w_eco142584, w_eco142585, w_eco142586, w_eco142587, w_eco142588, w_eco142589, w_eco142590, w_eco142591, w_eco142592, w_eco142593, w_eco142594, w_eco142595, w_eco142596, w_eco142597, w_eco142598, w_eco142599, w_eco142600, w_eco142601, w_eco142602, w_eco142603, w_eco142604, w_eco142605, w_eco142606, w_eco142607, w_eco142608, w_eco142609, w_eco142610, w_eco142611, w_eco142612, w_eco142613, w_eco142614, w_eco142615, w_eco142616, w_eco142617, w_eco142618, w_eco142619, w_eco142620, w_eco142621, w_eco142622, w_eco142623, w_eco142624, w_eco142625, w_eco142626, w_eco142627, w_eco142628, w_eco142629, w_eco142630, w_eco142631, w_eco142632, w_eco142633, w_eco142634, w_eco142635, w_eco142636, w_eco142637, w_eco142638, w_eco142639, w_eco142640, w_eco142641, w_eco142642, w_eco142643, w_eco142644, w_eco142645, w_eco142646, w_eco142647, w_eco142648, w_eco142649, w_eco142650, w_eco142651, w_eco142652, w_eco142653, w_eco142654, w_eco142655, w_eco142656, w_eco142657, w_eco142658, w_eco142659, w_eco142660, w_eco142661, w_eco142662, w_eco142663, w_eco142664, w_eco142665, w_eco142666, w_eco142667, w_eco142668, w_eco142669, w_eco142670, w_eco142671, w_eco142672, w_eco142673, w_eco142674, w_eco142675, w_eco142676, w_eco142677, w_eco142678, w_eco142679, w_eco142680, w_eco142681, w_eco142682, w_eco142683, w_eco142684, w_eco142685, w_eco142686, w_eco142687, w_eco142688, w_eco142689, w_eco142690, w_eco142691, w_eco142692, w_eco142693, w_eco142694, w_eco142695, w_eco142696, w_eco142697, w_eco142698, w_eco142699, w_eco142700, w_eco142701, w_eco142702, w_eco142703, w_eco142704, w_eco142705, w_eco142706, w_eco142707, w_eco142708, w_eco142709, w_eco142710, w_eco142711, w_eco142712, w_eco142713, w_eco142714, w_eco142715, w_eco142716, w_eco142717, w_eco142718, w_eco142719, w_eco142720, w_eco142721, w_eco142722, w_eco142723, w_eco142724, w_eco142725, w_eco142726, w_eco142727, w_eco142728, w_eco142729, w_eco142730, w_eco142731, w_eco142732, w_eco142733, w_eco142734, w_eco142735, w_eco142736, w_eco142737, w_eco142738, w_eco142739, w_eco142740, w_eco142741, w_eco142742, w_eco142743, w_eco142744, w_eco142745, w_eco142746, w_eco142747, w_eco142748, w_eco142749, w_eco142750, w_eco142751, w_eco142752, w_eco142753, w_eco142754, w_eco142755, w_eco142756, w_eco142757, w_eco142758, w_eco142759, w_eco142760, w_eco142761, w_eco142762, w_eco142763, w_eco142764, w_eco142765, w_eco142766, w_eco142767, w_eco142768, w_eco142769, w_eco142770, w_eco142771, w_eco142772, w_eco142773, w_eco142774, w_eco142775, w_eco142776, w_eco142777, w_eco142778, w_eco142779, w_eco142780, w_eco142781, w_eco142782, w_eco142783, w_eco142784, w_eco142785, w_eco142786, w_eco142787, w_eco142788, w_eco142789, w_eco142790, w_eco142791, w_eco142792, w_eco142793, w_eco142794, w_eco142795, w_eco142796, w_eco142797, w_eco142798, w_eco142799, w_eco142800, w_eco142801, w_eco142802, w_eco142803, w_eco142804, w_eco142805, w_eco142806, w_eco142807, w_eco142808, w_eco142809, w_eco142810, w_eco142811, w_eco142812, w_eco142813, w_eco142814, w_eco142815, w_eco142816, w_eco142817, w_eco142818, w_eco142819, w_eco142820, w_eco142821, w_eco142822, w_eco142823, w_eco142824, w_eco142825, w_eco142826, w_eco142827, w_eco142828, w_eco142829, w_eco142830, w_eco142831, w_eco142832, w_eco142833, w_eco142834, w_eco142835, w_eco142836, w_eco142837, w_eco142838, w_eco142839, w_eco142840, w_eco142841, w_eco142842, w_eco142843, w_eco142844, w_eco142845, w_eco142846, w_eco142847, w_eco142848, w_eco142849, w_eco142850, w_eco142851, w_eco142852, w_eco142853, w_eco142854, w_eco142855, w_eco142856, w_eco142857, w_eco142858, w_eco142859, w_eco142860, w_eco142861, w_eco142862, w_eco142863, w_eco142864, w_eco142865, w_eco142866, w_eco142867, w_eco142868, w_eco142869, w_eco142870, w_eco142871, w_eco142872, w_eco142873, w_eco142874, w_eco142875, w_eco142876, w_eco142877, w_eco142878, w_eco142879, w_eco142880, w_eco142881, w_eco142882, w_eco142883, w_eco142884, w_eco142885, w_eco142886, w_eco142887, w_eco142888, w_eco142889, w_eco142890, w_eco142891, w_eco142892, w_eco142893, w_eco142894, w_eco142895, w_eco142896, w_eco142897, w_eco142898, w_eco142899, w_eco142900, w_eco142901, w_eco142902, w_eco142903, w_eco142904, w_eco142905, w_eco142906, w_eco142907, w_eco142908, w_eco142909, w_eco142910, w_eco142911, w_eco142912, w_eco142913, w_eco142914, w_eco142915, w_eco142916, w_eco142917, w_eco142918, w_eco142919, w_eco142920, w_eco142921, w_eco142922, w_eco142923, w_eco142924, w_eco142925, w_eco142926, w_eco142927, w_eco142928, w_eco142929, w_eco142930, w_eco142931, w_eco142932, w_eco142933, w_eco142934, w_eco142935, w_eco142936, w_eco142937, w_eco142938, w_eco142939, w_eco142940, w_eco142941, w_eco142942, w_eco142943, w_eco142944, w_eco142945, w_eco142946, w_eco142947, w_eco142948, w_eco142949, w_eco142950, w_eco142951, w_eco142952, w_eco142953, w_eco142954, w_eco142955, w_eco142956, w_eco142957, w_eco142958, w_eco142959, w_eco142960, w_eco142961, w_eco142962, w_eco142963, w_eco142964, w_eco142965, w_eco142966, w_eco142967, w_eco142968, w_eco142969, w_eco142970, w_eco142971, w_eco142972, w_eco142973, w_eco142974, w_eco142975, w_eco142976, w_eco142977, w_eco142978, w_eco142979, w_eco142980, w_eco142981, w_eco142982, w_eco142983, w_eco142984, w_eco142985, w_eco142986, w_eco142987, w_eco142988, w_eco142989, w_eco142990, w_eco142991, w_eco142992, w_eco142993, w_eco142994, w_eco142995, w_eco142996, w_eco142997, w_eco142998, w_eco142999, w_eco143000, w_eco143001, w_eco143002, w_eco143003, w_eco143004, w_eco143005, w_eco143006, w_eco143007, w_eco143008, w_eco143009, w_eco143010, w_eco143011, w_eco143012, w_eco143013, w_eco143014, w_eco143015, w_eco143016, w_eco143017, w_eco143018, w_eco143019, w_eco143020, w_eco143021, w_eco143022, w_eco143023, w_eco143024, w_eco143025, w_eco143026, w_eco143027, w_eco143028, w_eco143029, w_eco143030, w_eco143031, w_eco143032, w_eco143033, w_eco143034, w_eco143035, w_eco143036, w_eco143037, w_eco143038, w_eco143039, w_eco143040, w_eco143041, w_eco143042, w_eco143043, w_eco143044, w_eco143045, w_eco143046, w_eco143047, w_eco143048, w_eco143049, w_eco143050, w_eco143051, w_eco143052, w_eco143053, w_eco143054, w_eco143055, w_eco143056, w_eco143057, w_eco143058, w_eco143059, w_eco143060, w_eco143061, w_eco143062, w_eco143063, w_eco143064, w_eco143065, w_eco143066, w_eco143067, w_eco143068, w_eco143069, w_eco143070, w_eco143071, w_eco143072, w_eco143073, w_eco143074, w_eco143075, w_eco143076, w_eco143077, w_eco143078, w_eco143079, w_eco143080, w_eco143081, w_eco143082, w_eco143083, w_eco143084, w_eco143085, w_eco143086, w_eco143087, w_eco143088, w_eco143089, w_eco143090, w_eco143091, w_eco143092, w_eco143093, w_eco143094, w_eco143095, w_eco143096, w_eco143097, w_eco143098, w_eco143099, w_eco143100, w_eco143101, w_eco143102, w_eco143103, w_eco143104, w_eco143105, w_eco143106, w_eco143107, w_eco143108, w_eco143109, w_eco143110, w_eco143111, w_eco143112, w_eco143113, w_eco143114, w_eco143115, w_eco143116, w_eco143117, w_eco143118, w_eco143119, w_eco143120, w_eco143121, w_eco143122, w_eco143123, w_eco143124, w_eco143125, w_eco143126, w_eco143127, w_eco143128, w_eco143129, w_eco143130, w_eco143131, w_eco143132, w_eco143133, w_eco143134, w_eco143135, w_eco143136, w_eco143137, w_eco143138, w_eco143139, w_eco143140, w_eco143141, w_eco143142, w_eco143143, w_eco143144, w_eco143145, w_eco143146, w_eco143147, w_eco143148, w_eco143149, w_eco143150, w_eco143151, w_eco143152, w_eco143153, w_eco143154, w_eco143155, w_eco143156, w_eco143157, w_eco143158, w_eco143159, w_eco143160, w_eco143161, w_eco143162, w_eco143163, w_eco143164, w_eco143165, w_eco143166, w_eco143167, w_eco143168, w_eco143169, w_eco143170, w_eco143171, w_eco143172, w_eco143173, w_eco143174, w_eco143175, w_eco143176, w_eco143177, w_eco143178, w_eco143179, w_eco143180, w_eco143181, w_eco143182, w_eco143183, w_eco143184, w_eco143185, w_eco143186, w_eco143187, w_eco143188, w_eco143189, w_eco143190, w_eco143191, w_eco143192, w_eco143193, w_eco143194, w_eco143195, w_eco143196, w_eco143197, w_eco143198, w_eco143199, w_eco143200, w_eco143201, w_eco143202, w_eco143203, w_eco143204, w_eco143205, w_eco143206, w_eco143207, w_eco143208, w_eco143209, w_eco143210, w_eco143211, w_eco143212, w_eco143213, w_eco143214, w_eco143215, w_eco143216, w_eco143217, w_eco143218, w_eco143219, w_eco143220, w_eco143221, w_eco143222, w_eco143223, w_eco143224, w_eco143225, w_eco143226, w_eco143227, w_eco143228, w_eco143229, w_eco143230, w_eco143231, w_eco143232, w_eco143233, w_eco143234, w_eco143235, w_eco143236, w_eco143237, w_eco143238, w_eco143239, w_eco143240, w_eco143241, w_eco143242, w_eco143243, w_eco143244, w_eco143245, w_eco143246, w_eco143247, w_eco143248, w_eco143249, w_eco143250, w_eco143251, w_eco143252, w_eco143253, w_eco143254, w_eco143255, w_eco143256, w_eco143257, w_eco143258, w_eco143259, w_eco143260, w_eco143261, w_eco143262, w_eco143263, w_eco143264, w_eco143265, w_eco143266, w_eco143267, w_eco143268, w_eco143269, w_eco143270, w_eco143271, w_eco143272, w_eco143273, w_eco143274, w_eco143275, w_eco143276, w_eco143277, w_eco143278, w_eco143279, w_eco143280, w_eco143281, w_eco143282, w_eco143283, w_eco143284, w_eco143285, w_eco143286, w_eco143287, w_eco143288, w_eco143289, w_eco143290, w_eco143291, w_eco143292, w_eco143293, w_eco143294, w_eco143295, w_eco143296, w_eco143297, w_eco143298, w_eco143299, w_eco143300, w_eco143301, w_eco143302, w_eco143303, w_eco143304, w_eco143305, w_eco143306, w_eco143307, w_eco143308, w_eco143309, w_eco143310, w_eco143311, w_eco143312, w_eco143313, w_eco143314, w_eco143315, w_eco143316, w_eco143317, w_eco143318, w_eco143319, w_eco143320, w_eco143321, w_eco143322, w_eco143323, w_eco143324, w_eco143325, w_eco143326, w_eco143327, w_eco143328, w_eco143329, w_eco143330, w_eco143331, w_eco143332, w_eco143333, w_eco143334, w_eco143335, w_eco143336, w_eco143337, w_eco143338, w_eco143339, w_eco143340, w_eco143341, w_eco143342, w_eco143343, w_eco143344, w_eco143345, w_eco143346, w_eco143347, w_eco143348, w_eco143349, w_eco143350, w_eco143351, w_eco143352, w_eco143353, w_eco143354, w_eco143355, w_eco143356, w_eco143357, w_eco143358, w_eco143359, w_eco143360, w_eco143361, w_eco143362, w_eco143363, w_eco143364, w_eco143365, w_eco143366, w_eco143367, w_eco143368, w_eco143369, w_eco143370, w_eco143371, w_eco143372, w_eco143373, w_eco143374, w_eco143375, w_eco143376, w_eco143377, w_eco143378, w_eco143379, w_eco143380, w_eco143381, w_eco143382, w_eco143383, w_eco143384, w_eco143385, w_eco143386, w_eco143387, w_eco143388, w_eco143389, w_eco143390, w_eco143391, w_eco143392, w_eco143393, w_eco143394, w_eco143395, w_eco143396, w_eco143397, w_eco143398, w_eco143399, w_eco143400, w_eco143401, w_eco143402, w_eco143403, w_eco143404, w_eco143405, w_eco143406, w_eco143407, w_eco143408, w_eco143409, w_eco143410, w_eco143411, w_eco143412, w_eco143413, w_eco143414, w_eco143415, w_eco143416, w_eco143417, w_eco143418, w_eco143419, w_eco143420, w_eco143421, w_eco143422, w_eco143423, w_eco143424, w_eco143425, w_eco143426, w_eco143427, w_eco143428, w_eco143429, w_eco143430, w_eco143431, w_eco143432, w_eco143433, w_eco143434, w_eco143435, w_eco143436, w_eco143437, w_eco143438, w_eco143439, w_eco143440, w_eco143441, w_eco143442, w_eco143443, w_eco143444, w_eco143445, w_eco143446, w_eco143447, w_eco143448, w_eco143449, w_eco143450, w_eco143451, w_eco143452, w_eco143453, w_eco143454, w_eco143455, w_eco143456, w_eco143457, w_eco143458, w_eco143459, w_eco143460, w_eco143461, w_eco143462, w_eco143463, w_eco143464, w_eco143465, w_eco143466, w_eco143467, w_eco143468, w_eco143469, w_eco143470, w_eco143471, w_eco143472, w_eco143473, w_eco143474, w_eco143475, w_eco143476, w_eco143477, w_eco143478, w_eco143479, w_eco143480, w_eco143481, w_eco143482, w_eco143483, w_eco143484, w_eco143485, w_eco143486, w_eco143487, w_eco143488, w_eco143489, w_eco143490, w_eco143491, w_eco143492, w_eco143493, w_eco143494, w_eco143495, w_eco143496, w_eco143497, w_eco143498, w_eco143499, w_eco143500, w_eco143501, w_eco143502, w_eco143503, w_eco143504, w_eco143505, w_eco143506, w_eco143507, w_eco143508, w_eco143509, w_eco143510, w_eco143511, w_eco143512, w_eco143513, w_eco143514, w_eco143515, w_eco143516, w_eco143517, w_eco143518, w_eco143519, w_eco143520, w_eco143521, w_eco143522, w_eco143523, w_eco143524, w_eco143525, w_eco143526, w_eco143527, w_eco143528, w_eco143529, w_eco143530, w_eco143531, w_eco143532, w_eco143533, w_eco143534, w_eco143535, w_eco143536, w_eco143537, w_eco143538, w_eco143539, w_eco143540, w_eco143541, w_eco143542, w_eco143543, w_eco143544, w_eco143545, w_eco143546, w_eco143547, w_eco143548, w_eco143549, w_eco143550, w_eco143551, w_eco143552, w_eco143553, w_eco143554, w_eco143555, w_eco143556, w_eco143557, w_eco143558, w_eco143559, w_eco143560, w_eco143561, w_eco143562, w_eco143563, w_eco143564, w_eco143565, w_eco143566, w_eco143567, w_eco143568, w_eco143569, w_eco143570, w_eco143571, w_eco143572, w_eco143573, w_eco143574, w_eco143575, w_eco143576, w_eco143577, w_eco143578, w_eco143579, w_eco143580, w_eco143581, w_eco143582, w_eco143583, w_eco143584, w_eco143585, w_eco143586, w_eco143587, w_eco143588, w_eco143589, w_eco143590, w_eco143591, w_eco143592, w_eco143593, w_eco143594, w_eco143595, w_eco143596, w_eco143597, w_eco143598, w_eco143599, w_eco143600, w_eco143601, w_eco143602, w_eco143603, w_eco143604, w_eco143605, w_eco143606, w_eco143607, w_eco143608, w_eco143609, w_eco143610, w_eco143611, w_eco143612, w_eco143613, w_eco143614, w_eco143615, w_eco143616, w_eco143617, w_eco143618, w_eco143619, w_eco143620, w_eco143621, w_eco143622, w_eco143623, w_eco143624, w_eco143625, w_eco143626, w_eco143627, w_eco143628, w_eco143629, w_eco143630, w_eco143631, w_eco143632, w_eco143633, w_eco143634, w_eco143635, w_eco143636, w_eco143637, w_eco143638, w_eco143639, w_eco143640, w_eco143641, w_eco143642, w_eco143643, w_eco143644, w_eco143645, w_eco143646, w_eco143647, w_eco143648, w_eco143649, w_eco143650, w_eco143651, w_eco143652, w_eco143653, w_eco143654, w_eco143655, w_eco143656, w_eco143657, w_eco143658, w_eco143659, w_eco143660, w_eco143661, w_eco143662, w_eco143663, w_eco143664, w_eco143665, w_eco143666, w_eco143667, w_eco143668, w_eco143669, w_eco143670, w_eco143671, w_eco143672, w_eco143673, w_eco143674, w_eco143675, w_eco143676, w_eco143677, w_eco143678, w_eco143679, w_eco143680, w_eco143681, w_eco143682, w_eco143683, w_eco143684, w_eco143685, w_eco143686, w_eco143687, w_eco143688, w_eco143689, w_eco143690, w_eco143691, w_eco143692, w_eco143693, w_eco143694, w_eco143695, w_eco143696, w_eco143697, w_eco143698, w_eco143699, w_eco143700, w_eco143701, w_eco143702, w_eco143703, w_eco143704, w_eco143705, w_eco143706, w_eco143707, w_eco143708, w_eco143709, w_eco143710, w_eco143711, w_eco143712, w_eco143713, w_eco143714, w_eco143715, w_eco143716, w_eco143717, w_eco143718, w_eco143719, w_eco143720, w_eco143721, w_eco143722, w_eco143723, w_eco143724, w_eco143725, w_eco143726, w_eco143727, w_eco143728, w_eco143729, w_eco143730, w_eco143731, w_eco143732, w_eco143733, w_eco143734, w_eco143735, w_eco143736, w_eco143737, w_eco143738, w_eco143739, w_eco143740, w_eco143741, w_eco143742, w_eco143743, w_eco143744, w_eco143745, w_eco143746, w_eco143747, w_eco143748, w_eco143749, w_eco143750, w_eco143751, w_eco143752, w_eco143753, w_eco143754, w_eco143755, w_eco143756, w_eco143757, w_eco143758, w_eco143759, w_eco143760, w_eco143761, w_eco143762, w_eco143763, w_eco143764, w_eco143765, w_eco143766, w_eco143767, w_eco143768, w_eco143769, w_eco143770, w_eco143771, w_eco143772, w_eco143773, w_eco143774, w_eco143775, w_eco143776, w_eco143777, w_eco143778, w_eco143779, w_eco143780, w_eco143781, w_eco143782, w_eco143783, w_eco143784, w_eco143785, w_eco143786, w_eco143787, w_eco143788, w_eco143789, w_eco143790, w_eco143791, w_eco143792, w_eco143793, w_eco143794, w_eco143795, w_eco143796, w_eco143797, w_eco143798, w_eco143799, w_eco143800, w_eco143801, w_eco143802, w_eco143803, w_eco143804, w_eco143805, w_eco143806, w_eco143807, w_eco143808, w_eco143809, w_eco143810, w_eco143811, w_eco143812, w_eco143813, w_eco143814, w_eco143815, w_eco143816, w_eco143817, w_eco143818, w_eco143819, w_eco143820, w_eco143821, w_eco143822, w_eco143823, w_eco143824, w_eco143825, w_eco143826, w_eco143827, w_eco143828, w_eco143829, w_eco143830, w_eco143831, w_eco143832, w_eco143833, w_eco143834, w_eco143835, w_eco143836, w_eco143837, w_eco143838, w_eco143839, w_eco143840, w_eco143841, w_eco143842, w_eco143843, w_eco143844, w_eco143845, w_eco143846, w_eco143847, w_eco143848, w_eco143849, w_eco143850, w_eco143851, w_eco143852, w_eco143853, w_eco143854, w_eco143855, w_eco143856, w_eco143857, w_eco143858, w_eco143859, w_eco143860, w_eco143861, w_eco143862, w_eco143863, w_eco143864, w_eco143865, w_eco143866, w_eco143867, w_eco143868, w_eco143869, w_eco143870, w_eco143871, w_eco143872, w_eco143873, w_eco143874, w_eco143875, w_eco143876, w_eco143877, w_eco143878, w_eco143879, w_eco143880, w_eco143881, w_eco143882, w_eco143883, w_eco143884, w_eco143885, w_eco143886, w_eco143887, w_eco143888, w_eco143889, w_eco143890, w_eco143891, w_eco143892, w_eco143893, w_eco143894, w_eco143895, w_eco143896, w_eco143897, w_eco143898, w_eco143899, w_eco143900, w_eco143901, w_eco143902, w_eco143903, w_eco143904, w_eco143905, w_eco143906, w_eco143907, w_eco143908, w_eco143909, w_eco143910, w_eco143911, w_eco143912, w_eco143913, w_eco143914, w_eco143915, w_eco143916, w_eco143917, w_eco143918, w_eco143919, w_eco143920, w_eco143921, w_eco143922, w_eco143923, w_eco143924, w_eco143925, w_eco143926, w_eco143927, w_eco143928, w_eco143929, w_eco143930, w_eco143931, w_eco143932, w_eco143933, w_eco143934, w_eco143935, w_eco143936, w_eco143937, w_eco143938, w_eco143939, w_eco143940, w_eco143941, w_eco143942, w_eco143943, w_eco143944, w_eco143945, w_eco143946, w_eco143947, w_eco143948, w_eco143949, w_eco143950, w_eco143951, w_eco143952, w_eco143953, w_eco143954, w_eco143955, w_eco143956, w_eco143957, w_eco143958, w_eco143959, w_eco143960, w_eco143961, w_eco143962, w_eco143963, w_eco143964, w_eco143965, w_eco143966, w_eco143967, w_eco143968, w_eco143969, w_eco143970, w_eco143971, w_eco143972, w_eco143973, w_eco143974, w_eco143975, w_eco143976, w_eco143977, w_eco143978, w_eco143979, w_eco143980, w_eco143981, w_eco143982, w_eco143983, w_eco143984, w_eco143985, w_eco143986, w_eco143987, w_eco143988, w_eco143989, w_eco143990, w_eco143991, w_eco143992, w_eco143993, w_eco143994, w_eco143995, w_eco143996, w_eco143997, w_eco143998, w_eco143999, w_eco144000, w_eco144001, w_eco144002, w_eco144003, w_eco144004, w_eco144005, w_eco144006, w_eco144007, w_eco144008, w_eco144009, w_eco144010, w_eco144011, w_eco144012, w_eco144013, w_eco144014, w_eco144015, w_eco144016, w_eco144017, w_eco144018, w_eco144019, w_eco144020, w_eco144021, w_eco144022, w_eco144023, w_eco144024, w_eco144025, w_eco144026, w_eco144027, w_eco144028, w_eco144029, w_eco144030, w_eco144031, w_eco144032, w_eco144033, w_eco144034, w_eco144035, w_eco144036, w_eco144037, w_eco144038, w_eco144039, w_eco144040, w_eco144041, w_eco144042, w_eco144043, w_eco144044, w_eco144045, w_eco144046, w_eco144047, w_eco144048, w_eco144049, w_eco144050, w_eco144051, w_eco144052, w_eco144053, w_eco144054, w_eco144055, w_eco144056, w_eco144057, w_eco144058, w_eco144059, w_eco144060, w_eco144061, w_eco144062, w_eco144063, w_eco144064, w_eco144065, w_eco144066, w_eco144067, w_eco144068, w_eco144069, w_eco144070, w_eco144071, w_eco144072, w_eco144073, w_eco144074, w_eco144075, w_eco144076, w_eco144077, w_eco144078, w_eco144079, w_eco144080, w_eco144081, w_eco144082, w_eco144083, w_eco144084, w_eco144085, w_eco144086, w_eco144087, w_eco144088, w_eco144089, w_eco144090, w_eco144091, w_eco144092, w_eco144093, w_eco144094, w_eco144095, w_eco144096, w_eco144097, w_eco144098, w_eco144099, w_eco144100, w_eco144101, w_eco144102, w_eco144103, w_eco144104, w_eco144105, w_eco144106, w_eco144107, w_eco144108, w_eco144109, w_eco144110, w_eco144111, w_eco144112, w_eco144113, w_eco144114, w_eco144115, w_eco144116, w_eco144117, w_eco144118, w_eco144119, w_eco144120, w_eco144121, w_eco144122, w_eco144123, w_eco144124, w_eco144125, w_eco144126, w_eco144127, w_eco144128, w_eco144129, w_eco144130, w_eco144131, w_eco144132, w_eco144133, w_eco144134, w_eco144135, w_eco144136, w_eco144137, w_eco144138, w_eco144139, w_eco144140, w_eco144141, w_eco144142, w_eco144143, w_eco144144, w_eco144145, w_eco144146, w_eco144147, w_eco144148, w_eco144149, w_eco144150, w_eco144151, w_eco144152, w_eco144153, w_eco144154, w_eco144155, w_eco144156, w_eco144157, w_eco144158, w_eco144159, w_eco144160, w_eco144161, w_eco144162, w_eco144163, w_eco144164, w_eco144165, w_eco144166, w_eco144167, w_eco144168, w_eco144169, w_eco144170, w_eco144171, w_eco144172, w_eco144173, w_eco144174, w_eco144175, w_eco144176, w_eco144177, w_eco144178, w_eco144179, w_eco144180, w_eco144181, w_eco144182, w_eco144183, w_eco144184, w_eco144185, w_eco144186, w_eco144187, w_eco144188, w_eco144189, w_eco144190, w_eco144191, w_eco144192, w_eco144193, w_eco144194, w_eco144195, w_eco144196, w_eco144197, w_eco144198, w_eco144199, w_eco144200, w_eco144201, w_eco144202, w_eco144203, w_eco144204, w_eco144205, w_eco144206, w_eco144207, w_eco144208, w_eco144209, w_eco144210, w_eco144211, w_eco144212, w_eco144213, w_eco144214, w_eco144215, w_eco144216, w_eco144217, w_eco144218, w_eco144219, w_eco144220, w_eco144221, w_eco144222, w_eco144223, w_eco144224, w_eco144225, w_eco144226, w_eco144227, w_eco144228, w_eco144229, w_eco144230, w_eco144231, w_eco144232, w_eco144233, w_eco144234, w_eco144235, w_eco144236, w_eco144237, w_eco144238, w_eco144239, w_eco144240, w_eco144241, w_eco144242, w_eco144243, w_eco144244, w_eco144245, w_eco144246, w_eco144247, w_eco144248, w_eco144249, w_eco144250, w_eco144251, w_eco144252, w_eco144253, w_eco144254, w_eco144255, w_eco144256, w_eco144257, w_eco144258, w_eco144259, w_eco144260, w_eco144261, w_eco144262, w_eco144263, w_eco144264, w_eco144265, w_eco144266, w_eco144267, w_eco144268, w_eco144269, w_eco144270, w_eco144271, w_eco144272, w_eco144273, w_eco144274, w_eco144275, w_eco144276, w_eco144277, w_eco144278, w_eco144279, w_eco144280, w_eco144281, w_eco144282, w_eco144283, w_eco144284, w_eco144285, w_eco144286, w_eco144287, w_eco144288, w_eco144289, w_eco144290, w_eco144291, w_eco144292, w_eco144293, w_eco144294, w_eco144295, w_eco144296, w_eco144297, w_eco144298, w_eco144299, w_eco144300, w_eco144301, w_eco144302, w_eco144303, w_eco144304, w_eco144305, w_eco144306, w_eco144307, w_eco144308, w_eco144309, w_eco144310, w_eco144311, w_eco144312, w_eco144313, w_eco144314, w_eco144315, w_eco144316, w_eco144317, w_eco144318, w_eco144319, w_eco144320, w_eco144321, w_eco144322, w_eco144323, w_eco144324, w_eco144325, w_eco144326, w_eco144327, w_eco144328, w_eco144329, w_eco144330, w_eco144331, w_eco144332, w_eco144333, w_eco144334, w_eco144335, w_eco144336, w_eco144337, w_eco144338, w_eco144339, w_eco144340, w_eco144341, w_eco144342, w_eco144343, w_eco144344, w_eco144345, w_eco144346, w_eco144347, w_eco144348, w_eco144349, w_eco144350, w_eco144351, w_eco144352, w_eco144353, w_eco144354, w_eco144355, w_eco144356, w_eco144357, w_eco144358, w_eco144359, w_eco144360, w_eco144361, w_eco144362, w_eco144363, w_eco144364, w_eco144365, w_eco144366, w_eco144367, w_eco144368, w_eco144369, w_eco144370, w_eco144371, w_eco144372, w_eco144373, w_eco144374, w_eco144375, w_eco144376, w_eco144377, w_eco144378, w_eco144379, w_eco144380, w_eco144381, w_eco144382, w_eco144383, w_eco144384, w_eco144385, w_eco144386, w_eco144387, w_eco144388, w_eco144389, w_eco144390, w_eco144391, w_eco144392, w_eco144393, w_eco144394, w_eco144395, w_eco144396, w_eco144397, w_eco144398, w_eco144399, w_eco144400, w_eco144401, w_eco144402, w_eco144403, w_eco144404, w_eco144405, w_eco144406, w_eco144407, w_eco144408, w_eco144409, w_eco144410, w_eco144411, w_eco144412, w_eco144413, w_eco144414, w_eco144415, w_eco144416, w_eco144417, w_eco144418, w_eco144419, w_eco144420, w_eco144421, w_eco144422, w_eco144423, w_eco144424, w_eco144425, w_eco144426, w_eco144427, w_eco144428, w_eco144429, w_eco144430, w_eco144431, w_eco144432, w_eco144433, w_eco144434, w_eco144435, w_eco144436, w_eco144437, w_eco144438, w_eco144439, w_eco144440, w_eco144441, w_eco144442, w_eco144443, w_eco144444, w_eco144445, w_eco144446, w_eco144447, w_eco144448, w_eco144449, w_eco144450, w_eco144451, w_eco144452, w_eco144453, w_eco144454, w_eco144455, w_eco144456, w_eco144457, w_eco144458, w_eco144459, w_eco144460, w_eco144461, w_eco144462, w_eco144463, w_eco144464, w_eco144465, w_eco144466, w_eco144467, w_eco144468, w_eco144469, w_eco144470, w_eco144471, w_eco144472, w_eco144473, w_eco144474, w_eco144475, w_eco144476, w_eco144477, w_eco144478, w_eco144479, w_eco144480, w_eco144481, w_eco144482, w_eco144483, w_eco144484, w_eco144485, w_eco144486, w_eco144487, w_eco144488, w_eco144489, w_eco144490, w_eco144491, w_eco144492, w_eco144493, w_eco144494, w_eco144495, w_eco144496, w_eco144497, w_eco144498, w_eco144499, w_eco144500, w_eco144501, w_eco144502, w_eco144503, w_eco144504, w_eco144505, w_eco144506, w_eco144507, w_eco144508, w_eco144509, w_eco144510, w_eco144511, w_eco144512, w_eco144513, w_eco144514, w_eco144515, w_eco144516, w_eco144517, w_eco144518, w_eco144519, w_eco144520, w_eco144521, w_eco144522, w_eco144523, w_eco144524, w_eco144525, w_eco144526, w_eco144527, w_eco144528, w_eco144529, w_eco144530, w_eco144531, w_eco144532, w_eco144533, w_eco144534, w_eco144535, w_eco144536, w_eco144537, w_eco144538, w_eco144539, w_eco144540, w_eco144541, w_eco144542, w_eco144543, w_eco144544, w_eco144545, w_eco144546, w_eco144547, w_eco144548, w_eco144549, w_eco144550, w_eco144551, w_eco144552, w_eco144553, w_eco144554, w_eco144555, w_eco144556, w_eco144557, w_eco144558, w_eco144559, w_eco144560, w_eco144561, w_eco144562, w_eco144563, w_eco144564, w_eco144565, w_eco144566, w_eco144567, w_eco144568, w_eco144569, w_eco144570, w_eco144571, w_eco144572, w_eco144573, w_eco144574, w_eco144575, w_eco144576, w_eco144577, w_eco144578, w_eco144579, w_eco144580, w_eco144581, w_eco144582, w_eco144583, w_eco144584, w_eco144585, w_eco144586, w_eco144587, w_eco144588, w_eco144589, w_eco144590, w_eco144591, w_eco144592, w_eco144593, w_eco144594, w_eco144595, w_eco144596, w_eco144597, w_eco144598, w_eco144599, w_eco144600, w_eco144601, w_eco144602, w_eco144603, w_eco144604, w_eco144605, w_eco144606, w_eco144607, w_eco144608, w_eco144609, w_eco144610, w_eco144611, w_eco144612, w_eco144613, w_eco144614, w_eco144615, w_eco144616, w_eco144617, w_eco144618, w_eco144619, w_eco144620, w_eco144621, w_eco144622, w_eco144623, w_eco144624, w_eco144625, w_eco144626, w_eco144627, w_eco144628, w_eco144629, w_eco144630, w_eco144631, w_eco144632, w_eco144633, w_eco144634, w_eco144635, w_eco144636, w_eco144637, w_eco144638, w_eco144639, w_eco144640, w_eco144641, w_eco144642, w_eco144643, w_eco144644, w_eco144645, w_eco144646, w_eco144647, w_eco144648, w_eco144649, w_eco144650, w_eco144651, w_eco144652, w_eco144653, w_eco144654, w_eco144655, w_eco144656, w_eco144657, w_eco144658, w_eco144659, w_eco144660, w_eco144661, w_eco144662, w_eco144663, w_eco144664, w_eco144665, w_eco144666, w_eco144667, w_eco144668, w_eco144669, w_eco144670, w_eco144671, w_eco144672, w_eco144673, w_eco144674, w_eco144675, w_eco144676, w_eco144677, w_eco144678, w_eco144679, w_eco144680, w_eco144681, w_eco144682, w_eco144683, w_eco144684, w_eco144685, w_eco144686, w_eco144687, w_eco144688, w_eco144689, w_eco144690, w_eco144691, w_eco144692, w_eco144693, w_eco144694, w_eco144695, w_eco144696, w_eco144697, w_eco144698, w_eco144699, w_eco144700, w_eco144701, w_eco144702, w_eco144703, w_eco144704, w_eco144705, w_eco144706, w_eco144707, w_eco144708, w_eco144709, w_eco144710, w_eco144711, w_eco144712, w_eco144713, w_eco144714, w_eco144715, w_eco144716, w_eco144717, w_eco144718, w_eco144719, w_eco144720, w_eco144721, w_eco144722, w_eco144723, w_eco144724, w_eco144725, w_eco144726, w_eco144727, w_eco144728, w_eco144729, w_eco144730, w_eco144731, w_eco144732, w_eco144733, w_eco144734, w_eco144735, w_eco144736, w_eco144737, w_eco144738, w_eco144739, w_eco144740, w_eco144741, w_eco144742, w_eco144743, w_eco144744, w_eco144745, w_eco144746, w_eco144747, w_eco144748, w_eco144749, w_eco144750, w_eco144751, w_eco144752, w_eco144753, w_eco144754, w_eco144755, w_eco144756, w_eco144757, w_eco144758, w_eco144759, w_eco144760, w_eco144761, w_eco144762, w_eco144763, w_eco144764, w_eco144765, w_eco144766, w_eco144767, w_eco144768, w_eco144769, w_eco144770, w_eco144771, w_eco144772, w_eco144773, w_eco144774, w_eco144775, w_eco144776, w_eco144777, w_eco144778, w_eco144779, w_eco144780, w_eco144781, w_eco144782, w_eco144783, w_eco144784, w_eco144785, w_eco144786, w_eco144787, w_eco144788, w_eco144789, w_eco144790, w_eco144791, w_eco144792, w_eco144793, w_eco144794, w_eco144795, w_eco144796, w_eco144797, w_eco144798, w_eco144799, w_eco144800, w_eco144801, w_eco144802, w_eco144803, w_eco144804, w_eco144805, w_eco144806, w_eco144807, w_eco144808, w_eco144809, w_eco144810, w_eco144811, w_eco144812, w_eco144813, w_eco144814, w_eco144815, w_eco144816, w_eco144817, w_eco144818, w_eco144819, w_eco144820, w_eco144821, w_eco144822, w_eco144823, w_eco144824, w_eco144825, w_eco144826, w_eco144827, w_eco144828, w_eco144829, w_eco144830, w_eco144831, w_eco144832, w_eco144833, w_eco144834, w_eco144835, w_eco144836, w_eco144837, w_eco144838, w_eco144839, w_eco144840, w_eco144841, w_eco144842, w_eco144843, w_eco144844, w_eco144845, w_eco144846, w_eco144847, w_eco144848, w_eco144849, w_eco144850, w_eco144851, w_eco144852, w_eco144853, w_eco144854, w_eco144855, w_eco144856, w_eco144857, w_eco144858, w_eco144859, w_eco144860, w_eco144861, w_eco144862, w_eco144863, w_eco144864, w_eco144865, w_eco144866, w_eco144867, w_eco144868, w_eco144869, w_eco144870, w_eco144871, w_eco144872, w_eco144873, w_eco144874, w_eco144875, w_eco144876, w_eco144877, w_eco144878, w_eco144879, w_eco144880, w_eco144881, w_eco144882, w_eco144883, w_eco144884, w_eco144885, w_eco144886, w_eco144887, w_eco144888, w_eco144889, w_eco144890, w_eco144891, w_eco144892, w_eco144893, w_eco144894, w_eco144895, w_eco144896, w_eco144897, w_eco144898, w_eco144899, w_eco144900, w_eco144901, w_eco144902, w_eco144903, w_eco144904, w_eco144905, w_eco144906, w_eco144907, w_eco144908, w_eco144909, w_eco144910, w_eco144911, w_eco144912, w_eco144913, w_eco144914, w_eco144915, w_eco144916, w_eco144917, w_eco144918, w_eco144919, w_eco144920, w_eco144921, w_eco144922, w_eco144923, w_eco144924, w_eco144925, w_eco144926, w_eco144927, w_eco144928, w_eco144929, w_eco144930, w_eco144931, w_eco144932, w_eco144933, w_eco144934, w_eco144935, w_eco144936, w_eco144937, w_eco144938, w_eco144939, w_eco144940, w_eco144941, w_eco144942, w_eco144943, w_eco144944, w_eco144945, w_eco144946, w_eco144947, w_eco144948, w_eco144949, w_eco144950, w_eco144951, w_eco144952, w_eco144953, w_eco144954, w_eco144955, w_eco144956, w_eco144957, w_eco144958, w_eco144959, w_eco144960, w_eco144961, w_eco144962, w_eco144963, w_eco144964, w_eco144965, w_eco144966, w_eco144967, w_eco144968, w_eco144969, w_eco144970, w_eco144971, w_eco144972, w_eco144973, w_eco144974, w_eco144975, w_eco144976, w_eco144977, w_eco144978, w_eco144979, w_eco144980, w_eco144981, w_eco144982, w_eco144983, w_eco144984, w_eco144985, w_eco144986, w_eco144987, w_eco144988, w_eco144989, w_eco144990, w_eco144991, w_eco144992, w_eco144993, w_eco144994, w_eco144995, w_eco144996, w_eco144997, w_eco144998, w_eco144999, w_eco145000, w_eco145001, w_eco145002, w_eco145003, w_eco145004, w_eco145005, w_eco145006, w_eco145007, w_eco145008, w_eco145009, w_eco145010, w_eco145011, w_eco145012, w_eco145013, w_eco145014, w_eco145015, w_eco145016, w_eco145017, w_eco145018, w_eco145019, w_eco145020, w_eco145021, w_eco145022, w_eco145023, w_eco145024, w_eco145025, w_eco145026, w_eco145027, w_eco145028, w_eco145029, w_eco145030, w_eco145031, w_eco145032, w_eco145033, w_eco145034, w_eco145035, w_eco145036, w_eco145037, w_eco145038, w_eco145039, w_eco145040, w_eco145041, w_eco145042, w_eco145043, w_eco145044, w_eco145045, w_eco145046, w_eco145047, w_eco145048, w_eco145049, w_eco145050, w_eco145051, w_eco145052, w_eco145053, w_eco145054, w_eco145055, w_eco145056, w_eco145057, w_eco145058, w_eco145059, w_eco145060, w_eco145061, w_eco145062, w_eco145063, w_eco145064, w_eco145065, w_eco145066, w_eco145067, w_eco145068, w_eco145069, w_eco145070, w_eco145071, w_eco145072, w_eco145073, w_eco145074, w_eco145075, w_eco145076, w_eco145077, w_eco145078, w_eco145079, w_eco145080, w_eco145081, w_eco145082, w_eco145083, w_eco145084, w_eco145085, w_eco145086, w_eco145087, w_eco145088, w_eco145089, w_eco145090, w_eco145091, w_eco145092, w_eco145093, w_eco145094, w_eco145095, w_eco145096, w_eco145097, w_eco145098, w_eco145099, w_eco145100, w_eco145101, w_eco145102, w_eco145103, w_eco145104, w_eco145105, w_eco145106, w_eco145107, w_eco145108, w_eco145109, w_eco145110, w_eco145111, w_eco145112, w_eco145113, w_eco145114, w_eco145115, w_eco145116, w_eco145117, w_eco145118, w_eco145119, w_eco145120, w_eco145121, w_eco145122, w_eco145123, w_eco145124, w_eco145125, w_eco145126, w_eco145127, w_eco145128, w_eco145129, w_eco145130, w_eco145131, w_eco145132, w_eco145133, w_eco145134, w_eco145135, w_eco145136, w_eco145137, w_eco145138, w_eco145139, w_eco145140, w_eco145141, w_eco145142, w_eco145143, w_eco145144, w_eco145145, w_eco145146, w_eco145147, w_eco145148, w_eco145149, w_eco145150, w_eco145151, w_eco145152, w_eco145153, w_eco145154, w_eco145155, w_eco145156, w_eco145157, w_eco145158, w_eco145159, w_eco145160, w_eco145161, w_eco145162, w_eco145163, w_eco145164, w_eco145165, w_eco145166, w_eco145167, w_eco145168, w_eco145169, w_eco145170, w_eco145171, w_eco145172, w_eco145173, w_eco145174, w_eco145175, w_eco145176, w_eco145177, w_eco145178, w_eco145179, w_eco145180, w_eco145181, w_eco145182, w_eco145183, w_eco145184, w_eco145185, w_eco145186, w_eco145187, w_eco145188, w_eco145189, w_eco145190, w_eco145191, w_eco145192, w_eco145193, w_eco145194, w_eco145195, w_eco145196, w_eco145197, w_eco145198, w_eco145199, w_eco145200, w_eco145201, w_eco145202, w_eco145203, w_eco145204, w_eco145205, w_eco145206, w_eco145207, w_eco145208, w_eco145209, w_eco145210, w_eco145211, w_eco145212, w_eco145213, w_eco145214, w_eco145215, w_eco145216, w_eco145217, w_eco145218, w_eco145219, w_eco145220, w_eco145221, w_eco145222, w_eco145223, w_eco145224, w_eco145225, w_eco145226, w_eco145227, w_eco145228, w_eco145229, w_eco145230, w_eco145231, w_eco145232, w_eco145233, w_eco145234, w_eco145235, w_eco145236, w_eco145237, w_eco145238, w_eco145239, w_eco145240, w_eco145241, w_eco145242, w_eco145243, w_eco145244, w_eco145245, w_eco145246, w_eco145247, w_eco145248, w_eco145249, w_eco145250, w_eco145251, w_eco145252, w_eco145253, w_eco145254, w_eco145255, w_eco145256, w_eco145257, w_eco145258, w_eco145259, w_eco145260, w_eco145261, w_eco145262, w_eco145263, w_eco145264, w_eco145265, w_eco145266, w_eco145267, w_eco145268, w_eco145269, w_eco145270, w_eco145271, w_eco145272, w_eco145273, w_eco145274, w_eco145275, w_eco145276, w_eco145277, w_eco145278, w_eco145279, w_eco145280, w_eco145281, w_eco145282, w_eco145283, w_eco145284, w_eco145285, w_eco145286, w_eco145287, w_eco145288, w_eco145289, w_eco145290, w_eco145291, w_eco145292, w_eco145293, w_eco145294, w_eco145295, w_eco145296, w_eco145297, w_eco145298, w_eco145299, w_eco145300, w_eco145301, w_eco145302, w_eco145303, w_eco145304, w_eco145305, w_eco145306, w_eco145307, w_eco145308, w_eco145309, w_eco145310, w_eco145311, w_eco145312, w_eco145313, w_eco145314, w_eco145315, w_eco145316, w_eco145317, w_eco145318, w_eco145319, w_eco145320, w_eco145321, w_eco145322, w_eco145323, w_eco145324, w_eco145325, w_eco145326, w_eco145327, w_eco145328, w_eco145329, w_eco145330, w_eco145331, w_eco145332, w_eco145333, w_eco145334, w_eco145335, w_eco145336, w_eco145337, w_eco145338, w_eco145339, w_eco145340, w_eco145341, w_eco145342, w_eco145343, w_eco145344, w_eco145345, w_eco145346, w_eco145347, w_eco145348, w_eco145349, w_eco145350, w_eco145351, w_eco145352, w_eco145353, w_eco145354, w_eco145355, w_eco145356, w_eco145357, w_eco145358, w_eco145359, w_eco145360, w_eco145361, w_eco145362, w_eco145363, w_eco145364, w_eco145365, w_eco145366, w_eco145367, w_eco145368, w_eco145369, w_eco145370, w_eco145371, w_eco145372, w_eco145373, w_eco145374, w_eco145375, w_eco145376, w_eco145377, w_eco145378, w_eco145379, w_eco145380, w_eco145381, w_eco145382, w_eco145383, w_eco145384, w_eco145385, w_eco145386, w_eco145387, w_eco145388, w_eco145389, w_eco145390, w_eco145391, w_eco145392, w_eco145393, w_eco145394, w_eco145395, w_eco145396, w_eco145397, w_eco145398, w_eco145399, w_eco145400, w_eco145401, w_eco145402, w_eco145403, w_eco145404, w_eco145405, w_eco145406, w_eco145407, w_eco145408, w_eco145409, w_eco145410, w_eco145411, w_eco145412, w_eco145413, w_eco145414, w_eco145415, w_eco145416, w_eco145417, w_eco145418, w_eco145419, w_eco145420, w_eco145421, w_eco145422, w_eco145423, w_eco145424, w_eco145425, w_eco145426, w_eco145427, w_eco145428, w_eco145429, w_eco145430, w_eco145431, w_eco145432, w_eco145433, w_eco145434, w_eco145435, w_eco145436, w_eco145437, w_eco145438, w_eco145439, w_eco145440, w_eco145441, w_eco145442, w_eco145443, w_eco145444, w_eco145445, w_eco145446, w_eco145447, w_eco145448, w_eco145449, w_eco145450, w_eco145451, w_eco145452, w_eco145453, w_eco145454, w_eco145455, w_eco145456, w_eco145457, w_eco145458, w_eco145459, w_eco145460, w_eco145461, w_eco145462, w_eco145463, w_eco145464, w_eco145465, w_eco145466, w_eco145467, w_eco145468, w_eco145469, w_eco145470, w_eco145471, w_eco145472, w_eco145473, w_eco145474, w_eco145475, w_eco145476, w_eco145477, w_eco145478, w_eco145479, w_eco145480, w_eco145481, w_eco145482, w_eco145483, w_eco145484, w_eco145485, w_eco145486, w_eco145487, w_eco145488, w_eco145489, w_eco145490, w_eco145491, w_eco145492, w_eco145493, w_eco145494, w_eco145495, w_eco145496, w_eco145497, w_eco145498, w_eco145499, w_eco145500, w_eco145501, w_eco145502, w_eco145503, w_eco145504, w_eco145505, w_eco145506, w_eco145507, w_eco145508, w_eco145509, w_eco145510, w_eco145511, w_eco145512, w_eco145513, w_eco145514, w_eco145515, w_eco145516, w_eco145517, w_eco145518, w_eco145519, w_eco145520, w_eco145521, w_eco145522, w_eco145523, w_eco145524, w_eco145525, w_eco145526, w_eco145527, w_eco145528, w_eco145529, w_eco145530, w_eco145531, w_eco145532, w_eco145533, w_eco145534, w_eco145535, w_eco145536, w_eco145537, w_eco145538, w_eco145539, w_eco145540, w_eco145541, w_eco145542, w_eco145543, w_eco145544, w_eco145545, w_eco145546, w_eco145547, w_eco145548, w_eco145549, w_eco145550, w_eco145551, w_eco145552, w_eco145553, w_eco145554, w_eco145555, w_eco145556, w_eco145557, w_eco145558, w_eco145559, w_eco145560, w_eco145561, w_eco145562, w_eco145563, w_eco145564, w_eco145565, w_eco145566, w_eco145567, w_eco145568, w_eco145569, w_eco145570, w_eco145571, w_eco145572, w_eco145573, w_eco145574, w_eco145575, w_eco145576, w_eco145577, w_eco145578, w_eco145579, w_eco145580, w_eco145581, w_eco145582, w_eco145583, w_eco145584, w_eco145585, w_eco145586, w_eco145587, w_eco145588, w_eco145589, w_eco145590, w_eco145591, w_eco145592, w_eco145593, w_eco145594, w_eco145595, w_eco145596, w_eco145597, w_eco145598, w_eco145599, w_eco145600, w_eco145601, w_eco145602, w_eco145603, w_eco145604, w_eco145605, w_eco145606, w_eco145607, w_eco145608, w_eco145609, w_eco145610, w_eco145611, w_eco145612, w_eco145613, w_eco145614, w_eco145615, w_eco145616, w_eco145617, w_eco145618, w_eco145619, w_eco145620, w_eco145621, w_eco145622, w_eco145623, w_eco145624, w_eco145625, w_eco145626, w_eco145627, w_eco145628, w_eco145629, w_eco145630, w_eco145631, w_eco145632, w_eco145633, w_eco145634, w_eco145635, w_eco145636, w_eco145637, w_eco145638, w_eco145639, w_eco145640, w_eco145641, w_eco145642, w_eco145643, w_eco145644, w_eco145645, w_eco145646, w_eco145647, w_eco145648, w_eco145649, w_eco145650, w_eco145651, w_eco145652, w_eco145653, w_eco145654, w_eco145655, w_eco145656, w_eco145657, w_eco145658, w_eco145659, w_eco145660, w_eco145661, w_eco145662, w_eco145663, w_eco145664, w_eco145665, w_eco145666, w_eco145667, w_eco145668, w_eco145669, w_eco145670, w_eco145671, w_eco145672, w_eco145673, w_eco145674, w_eco145675, w_eco145676, w_eco145677, w_eco145678, w_eco145679, w_eco145680, w_eco145681, w_eco145682, w_eco145683, w_eco145684, w_eco145685, w_eco145686, w_eco145687, w_eco145688, w_eco145689, w_eco145690, w_eco145691, w_eco145692, w_eco145693, w_eco145694, w_eco145695, w_eco145696, w_eco145697, w_eco145698, w_eco145699, w_eco145700, w_eco145701, w_eco145702, w_eco145703, w_eco145704, w_eco145705, w_eco145706, w_eco145707, w_eco145708, w_eco145709, w_eco145710, w_eco145711, w_eco145712, w_eco145713, w_eco145714, w_eco145715, w_eco145716, w_eco145717, w_eco145718, w_eco145719, w_eco145720, w_eco145721, w_eco145722, w_eco145723, w_eco145724, w_eco145725, w_eco145726, w_eco145727, w_eco145728, w_eco145729, w_eco145730, w_eco145731, w_eco145732, w_eco145733, w_eco145734, w_eco145735, w_eco145736, w_eco145737, w_eco145738, w_eco145739, w_eco145740, w_eco145741, w_eco145742, w_eco145743, w_eco145744, w_eco145745, w_eco145746, w_eco145747, w_eco145748, w_eco145749, w_eco145750, w_eco145751, w_eco145752, w_eco145753, w_eco145754, w_eco145755, w_eco145756, w_eco145757, w_eco145758, w_eco145759, w_eco145760, w_eco145761, w_eco145762, w_eco145763, w_eco145764, w_eco145765, w_eco145766, w_eco145767, w_eco145768, w_eco145769, w_eco145770, w_eco145771, w_eco145772, w_eco145773, w_eco145774, w_eco145775, w_eco145776, w_eco145777, w_eco145778, w_eco145779, w_eco145780, w_eco145781, w_eco145782, w_eco145783, w_eco145784, w_eco145785, w_eco145786, w_eco145787, w_eco145788, w_eco145789, w_eco145790, w_eco145791, w_eco145792, w_eco145793, w_eco145794, w_eco145795, w_eco145796, w_eco145797, w_eco145798, w_eco145799, w_eco145800, w_eco145801, w_eco145802, w_eco145803, w_eco145804, w_eco145805, w_eco145806, w_eco145807, w_eco145808, w_eco145809, w_eco145810, w_eco145811, w_eco145812, w_eco145813, w_eco145814, w_eco145815, w_eco145816, w_eco145817, w_eco145818, w_eco145819, w_eco145820, w_eco145821, w_eco145822, w_eco145823, w_eco145824, w_eco145825, w_eco145826, w_eco145827, w_eco145828, w_eco145829, w_eco145830, w_eco145831, w_eco145832, w_eco145833, w_eco145834, w_eco145835, w_eco145836, w_eco145837, w_eco145838, w_eco145839, w_eco145840, w_eco145841, w_eco145842, w_eco145843, w_eco145844, w_eco145845, w_eco145846, w_eco145847, w_eco145848, w_eco145849, w_eco145850, w_eco145851, w_eco145852, w_eco145853, w_eco145854, w_eco145855, w_eco145856, w_eco145857, w_eco145858, w_eco145859, w_eco145860, w_eco145861, w_eco145862, w_eco145863, w_eco145864, w_eco145865, w_eco145866, w_eco145867, w_eco145868, w_eco145869, w_eco145870, w_eco145871, w_eco145872, w_eco145873, w_eco145874, w_eco145875, w_eco145876, w_eco145877, w_eco145878, w_eco145879, w_eco145880, w_eco145881, w_eco145882, w_eco145883, w_eco145884, w_eco145885, w_eco145886, w_eco145887, w_eco145888, w_eco145889, w_eco145890, w_eco145891, w_eco145892, w_eco145893, w_eco145894, w_eco145895, w_eco145896, w_eco145897, w_eco145898, w_eco145899, w_eco145900, w_eco145901, w_eco145902, w_eco145903, w_eco145904, w_eco145905, w_eco145906, w_eco145907, w_eco145908, w_eco145909, w_eco145910, w_eco145911, w_eco145912, w_eco145913, w_eco145914, w_eco145915, w_eco145916, w_eco145917, w_eco145918, w_eco145919, w_eco145920, w_eco145921, w_eco145922, w_eco145923, w_eco145924, w_eco145925, w_eco145926, w_eco145927, w_eco145928, w_eco145929, w_eco145930, w_eco145931, w_eco145932, w_eco145933, w_eco145934, w_eco145935, w_eco145936, w_eco145937, w_eco145938, w_eco145939, w_eco145940, w_eco145941, w_eco145942, w_eco145943, w_eco145944, w_eco145945, w_eco145946, w_eco145947, w_eco145948, w_eco145949, w_eco145950, w_eco145951, w_eco145952, w_eco145953, w_eco145954, w_eco145955, w_eco145956, w_eco145957, w_eco145958, w_eco145959, w_eco145960, w_eco145961, w_eco145962, w_eco145963, w_eco145964, w_eco145965, w_eco145966, w_eco145967, w_eco145968, w_eco145969, w_eco145970, w_eco145971, w_eco145972, w_eco145973, w_eco145974, w_eco145975, w_eco145976, w_eco145977, w_eco145978, w_eco145979, w_eco145980, w_eco145981, w_eco145982, w_eco145983, w_eco145984, w_eco145985, w_eco145986, w_eco145987, w_eco145988, w_eco145989, w_eco145990, w_eco145991, w_eco145992, w_eco145993, w_eco145994, w_eco145995, w_eco145996, w_eco145997, w_eco145998, w_eco145999, w_eco146000, w_eco146001, w_eco146002, w_eco146003, w_eco146004, w_eco146005, w_eco146006, w_eco146007, w_eco146008, w_eco146009, w_eco146010, w_eco146011, w_eco146012, w_eco146013, w_eco146014, w_eco146015, w_eco146016, w_eco146017, w_eco146018, w_eco146019, w_eco146020, w_eco146021, w_eco146022, w_eco146023, w_eco146024, w_eco146025, w_eco146026, w_eco146027, w_eco146028, w_eco146029, w_eco146030, w_eco146031, w_eco146032, w_eco146033, w_eco146034, w_eco146035, w_eco146036, w_eco146037, w_eco146038, w_eco146039, w_eco146040, w_eco146041, w_eco146042, w_eco146043, w_eco146044, w_eco146045, w_eco146046, w_eco146047, w_eco146048, w_eco146049, w_eco146050, w_eco146051, w_eco146052, w_eco146053, w_eco146054, w_eco146055, w_eco146056, w_eco146057, w_eco146058, w_eco146059, w_eco146060, w_eco146061, w_eco146062, w_eco146063, w_eco146064, w_eco146065, w_eco146066, w_eco146067, w_eco146068, w_eco146069, w_eco146070, w_eco146071, w_eco146072, w_eco146073, w_eco146074, w_eco146075, w_eco146076, w_eco146077, w_eco146078, w_eco146079, w_eco146080, w_eco146081, w_eco146082, w_eco146083, w_eco146084, w_eco146085, w_eco146086, w_eco146087, w_eco146088, w_eco146089, w_eco146090, w_eco146091, w_eco146092, w_eco146093, w_eco146094, w_eco146095, w_eco146096, w_eco146097, w_eco146098, w_eco146099, w_eco146100, w_eco146101, w_eco146102, w_eco146103, w_eco146104, w_eco146105, w_eco146106, w_eco146107, w_eco146108, w_eco146109, w_eco146110, w_eco146111, w_eco146112, w_eco146113, w_eco146114, w_eco146115, w_eco146116, w_eco146117, w_eco146118, w_eco146119, w_eco146120, w_eco146121, w_eco146122, w_eco146123, w_eco146124, w_eco146125, w_eco146126, w_eco146127, w_eco146128, w_eco146129, w_eco146130, w_eco146131, w_eco146132, w_eco146133, w_eco146134, w_eco146135, w_eco146136, w_eco146137, w_eco146138, w_eco146139, w_eco146140, w_eco146141, w_eco146142, w_eco146143, w_eco146144, w_eco146145, w_eco146146, w_eco146147, w_eco146148, w_eco146149, w_eco146150, w_eco146151, w_eco146152, w_eco146153, w_eco146154, w_eco146155, w_eco146156, w_eco146157, w_eco146158, w_eco146159, w_eco146160, w_eco146161, w_eco146162, w_eco146163, w_eco146164, w_eco146165, w_eco146166, w_eco146167, w_eco146168, w_eco146169, w_eco146170, w_eco146171, w_eco146172, w_eco146173, w_eco146174, w_eco146175, w_eco146176, w_eco146177, w_eco146178, w_eco146179, w_eco146180, w_eco146181, w_eco146182, w_eco146183, w_eco146184, w_eco146185, w_eco146186, w_eco146187, w_eco146188, w_eco146189, w_eco146190, w_eco146191, w_eco146192, w_eco146193, w_eco146194, w_eco146195, w_eco146196, w_eco146197, w_eco146198, w_eco146199, w_eco146200, w_eco146201, w_eco146202, w_eco146203, w_eco146204, w_eco146205, w_eco146206, w_eco146207, w_eco146208, w_eco146209, w_eco146210, w_eco146211, w_eco146212, w_eco146213, w_eco146214, w_eco146215, w_eco146216, w_eco146217, w_eco146218, w_eco146219, w_eco146220, w_eco146221, w_eco146222, w_eco146223, w_eco146224, w_eco146225, w_eco146226, w_eco146227, w_eco146228, w_eco146229, w_eco146230, w_eco146231, w_eco146232, w_eco146233, w_eco146234, w_eco146235, w_eco146236, w_eco146237, w_eco146238, w_eco146239, w_eco146240, w_eco146241, w_eco146242, w_eco146243, w_eco146244, w_eco146245, w_eco146246, w_eco146247, w_eco146248, w_eco146249, w_eco146250, w_eco146251, w_eco146252, w_eco146253, w_eco146254, w_eco146255, w_eco146256, w_eco146257, w_eco146258, w_eco146259, w_eco146260, w_eco146261, w_eco146262, w_eco146263, w_eco146264, w_eco146265, w_eco146266, w_eco146267, w_eco146268, w_eco146269, w_eco146270, w_eco146271, w_eco146272, w_eco146273, w_eco146274, w_eco146275, w_eco146276, w_eco146277, w_eco146278, w_eco146279, w_eco146280, w_eco146281, w_eco146282, w_eco146283, w_eco146284, w_eco146285, w_eco146286, w_eco146287, w_eco146288, w_eco146289, w_eco146290, w_eco146291, w_eco146292, w_eco146293, w_eco146294, w_eco146295, w_eco146296, w_eco146297, w_eco146298, w_eco146299, w_eco146300, w_eco146301, w_eco146302, w_eco146303, w_eco146304, w_eco146305, w_eco146306, w_eco146307, w_eco146308, w_eco146309, w_eco146310, w_eco146311, w_eco146312, w_eco146313, w_eco146314, w_eco146315, w_eco146316, w_eco146317, w_eco146318, w_eco146319, w_eco146320, w_eco146321, w_eco146322, w_eco146323, w_eco146324, w_eco146325, w_eco146326, w_eco146327, w_eco146328, w_eco146329, w_eco146330, w_eco146331, w_eco146332, w_eco146333, w_eco146334, w_eco146335, w_eco146336, w_eco146337, w_eco146338, w_eco146339, w_eco146340, w_eco146341, w_eco146342, w_eco146343, w_eco146344, w_eco146345, w_eco146346, w_eco146347, w_eco146348, w_eco146349, w_eco146350, w_eco146351, w_eco146352, w_eco146353, w_eco146354, w_eco146355, w_eco146356, w_eco146357, w_eco146358, w_eco146359, w_eco146360, w_eco146361, w_eco146362, w_eco146363, w_eco146364, w_eco146365, w_eco146366, w_eco146367, w_eco146368, w_eco146369, w_eco146370, w_eco146371, w_eco146372, w_eco146373, w_eco146374, w_eco146375, w_eco146376, w_eco146377, w_eco146378, w_eco146379, w_eco146380, w_eco146381, w_eco146382, w_eco146383, w_eco146384, w_eco146385, w_eco146386, w_eco146387, w_eco146388, w_eco146389, w_eco146390, w_eco146391, w_eco146392, w_eco146393, w_eco146394, w_eco146395, w_eco146396, w_eco146397, w_eco146398, w_eco146399, w_eco146400, w_eco146401, w_eco146402, w_eco146403, w_eco146404, w_eco146405, w_eco146406, w_eco146407, w_eco146408, w_eco146409, w_eco146410, w_eco146411, w_eco146412, w_eco146413, w_eco146414, w_eco146415, w_eco146416, w_eco146417, w_eco146418, w_eco146419, w_eco146420, w_eco146421, w_eco146422, w_eco146423, w_eco146424, w_eco146425, w_eco146426, w_eco146427, w_eco146428, w_eco146429, w_eco146430, w_eco146431, w_eco146432, w_eco146433, w_eco146434, w_eco146435, w_eco146436, w_eco146437, w_eco146438, w_eco146439, w_eco146440, w_eco146441, w_eco146442, w_eco146443, w_eco146444, w_eco146445, w_eco146446, w_eco146447, w_eco146448, w_eco146449, w_eco146450, w_eco146451, w_eco146452, w_eco146453, w_eco146454, w_eco146455, w_eco146456, w_eco146457, w_eco146458, w_eco146459, w_eco146460, w_eco146461, w_eco146462, w_eco146463, w_eco146464, w_eco146465, w_eco146466, w_eco146467, w_eco146468, w_eco146469, w_eco146470, w_eco146471, w_eco146472, w_eco146473, w_eco146474, w_eco146475, w_eco146476, w_eco146477, w_eco146478, w_eco146479, w_eco146480, w_eco146481, w_eco146482, w_eco146483, w_eco146484, w_eco146485, w_eco146486, w_eco146487, w_eco146488, w_eco146489, w_eco146490, w_eco146491, w_eco146492, w_eco146493, w_eco146494, w_eco146495, w_eco146496, w_eco146497, w_eco146498, w_eco146499, w_eco146500, w_eco146501, w_eco146502, w_eco146503, w_eco146504, w_eco146505, w_eco146506, w_eco146507, w_eco146508, w_eco146509, w_eco146510, w_eco146511, w_eco146512, w_eco146513, w_eco146514, w_eco146515, w_eco146516, w_eco146517, w_eco146518, w_eco146519, w_eco146520, w_eco146521, w_eco146522, w_eco146523, w_eco146524, w_eco146525, w_eco146526, w_eco146527, w_eco146528, w_eco146529, w_eco146530, w_eco146531, w_eco146532, w_eco146533, w_eco146534, w_eco146535, w_eco146536, w_eco146537, w_eco146538, w_eco146539, w_eco146540, w_eco146541, w_eco146542, w_eco146543, w_eco146544, w_eco146545, w_eco146546, w_eco146547, w_eco146548, w_eco146549, w_eco146550, w_eco146551, w_eco146552, w_eco146553, w_eco146554, w_eco146555, w_eco146556, w_eco146557, w_eco146558, w_eco146559, w_eco146560, w_eco146561, w_eco146562, w_eco146563, w_eco146564, w_eco146565, w_eco146566, w_eco146567, w_eco146568, w_eco146569, w_eco146570, w_eco146571, w_eco146572, w_eco146573, w_eco146574, w_eco146575, w_eco146576, w_eco146577, w_eco146578, w_eco146579, w_eco146580, w_eco146581, w_eco146582, w_eco146583, w_eco146584, w_eco146585, w_eco146586, w_eco146587, w_eco146588, w_eco146589, w_eco146590, w_eco146591, w_eco146592, w_eco146593, w_eco146594, w_eco146595, w_eco146596, w_eco146597, w_eco146598, w_eco146599, w_eco146600, w_eco146601, w_eco146602, w_eco146603, w_eco146604, w_eco146605, w_eco146606, w_eco146607, w_eco146608, w_eco146609, w_eco146610, w_eco146611, w_eco146612, w_eco146613, w_eco146614, w_eco146615, w_eco146616, w_eco146617, w_eco146618, w_eco146619, w_eco146620, w_eco146621, w_eco146622, w_eco146623, w_eco146624, w_eco146625, w_eco146626, w_eco146627, w_eco146628, w_eco146629, w_eco146630, w_eco146631, w_eco146632, w_eco146633, w_eco146634, w_eco146635, w_eco146636, w_eco146637, w_eco146638, w_eco146639, w_eco146640, w_eco146641, w_eco146642, w_eco146643, w_eco146644, w_eco146645, w_eco146646, w_eco146647, w_eco146648, w_eco146649, w_eco146650, w_eco146651, w_eco146652, w_eco146653, w_eco146654, w_eco146655, w_eco146656, w_eco146657, w_eco146658, w_eco146659, w_eco146660, w_eco146661, w_eco146662, w_eco146663, w_eco146664, w_eco146665, w_eco146666, w_eco146667, w_eco146668, w_eco146669, w_eco146670, w_eco146671, w_eco146672, w_eco146673, w_eco146674, w_eco146675, w_eco146676, w_eco146677, w_eco146678, w_eco146679, w_eco146680, w_eco146681, w_eco146682, w_eco146683, w_eco146684, w_eco146685, w_eco146686, w_eco146687, w_eco146688, w_eco146689, w_eco146690, w_eco146691, w_eco146692, w_eco146693, w_eco146694, w_eco146695, w_eco146696, w_eco146697, w_eco146698, w_eco146699, w_eco146700, w_eco146701, w_eco146702, w_eco146703, w_eco146704, w_eco146705, w_eco146706, w_eco146707, w_eco146708, w_eco146709, w_eco146710, w_eco146711, w_eco146712, w_eco146713, w_eco146714, w_eco146715, w_eco146716, w_eco146717, w_eco146718, w_eco146719, w_eco146720, w_eco146721, w_eco146722, w_eco146723, w_eco146724, w_eco146725, w_eco146726, w_eco146727, w_eco146728, w_eco146729, w_eco146730, w_eco146731, w_eco146732, w_eco146733, w_eco146734, w_eco146735, w_eco146736, w_eco146737, w_eco146738, w_eco146739, w_eco146740, w_eco146741, w_eco146742, w_eco146743, w_eco146744, w_eco146745, w_eco146746, w_eco146747, w_eco146748, w_eco146749, w_eco146750, w_eco146751, w_eco146752, w_eco146753, w_eco146754, w_eco146755, w_eco146756, w_eco146757, w_eco146758, w_eco146759, w_eco146760, w_eco146761, w_eco146762, w_eco146763, w_eco146764, w_eco146765, w_eco146766, w_eco146767, w_eco146768, w_eco146769, w_eco146770, w_eco146771, w_eco146772, w_eco146773, w_eco146774, w_eco146775, w_eco146776, w_eco146777, w_eco146778, w_eco146779, w_eco146780, w_eco146781, w_eco146782, w_eco146783, w_eco146784, w_eco146785, w_eco146786, w_eco146787, w_eco146788, w_eco146789, w_eco146790, w_eco146791, w_eco146792, w_eco146793, w_eco146794, w_eco146795, w_eco146796, w_eco146797, w_eco146798, w_eco146799, w_eco146800, w_eco146801, w_eco146802, w_eco146803, w_eco146804, w_eco146805, w_eco146806, w_eco146807, w_eco146808, w_eco146809, w_eco146810, w_eco146811, w_eco146812, w_eco146813, w_eco146814, w_eco146815, w_eco146816, w_eco146817, w_eco146818, w_eco146819, w_eco146820, w_eco146821, w_eco146822, w_eco146823, w_eco146824, w_eco146825, w_eco146826, w_eco146827, w_eco146828, w_eco146829, w_eco146830, w_eco146831, w_eco146832, w_eco146833, w_eco146834, w_eco146835, w_eco146836, w_eco146837, w_eco146838, w_eco146839, w_eco146840, w_eco146841, w_eco146842, w_eco146843, w_eco146844, w_eco146845, w_eco146846, w_eco146847, w_eco146848, w_eco146849, w_eco146850, w_eco146851, w_eco146852, w_eco146853, w_eco146854, w_eco146855, w_eco146856, w_eco146857, w_eco146858, w_eco146859, w_eco146860, w_eco146861, w_eco146862, w_eco146863, w_eco146864, w_eco146865, w_eco146866, w_eco146867, w_eco146868, w_eco146869, w_eco146870, w_eco146871, w_eco146872, w_eco146873, w_eco146874, w_eco146875, w_eco146876, w_eco146877, w_eco146878, w_eco146879, w_eco146880, w_eco146881, w_eco146882, w_eco146883, w_eco146884, w_eco146885, w_eco146886, w_eco146887, w_eco146888, w_eco146889, w_eco146890, w_eco146891, w_eco146892, w_eco146893, w_eco146894, w_eco146895, w_eco146896, w_eco146897, w_eco146898, w_eco146899, w_eco146900, w_eco146901, w_eco146902, w_eco146903, w_eco146904, w_eco146905, w_eco146906, w_eco146907, w_eco146908, w_eco146909, w_eco146910, w_eco146911, w_eco146912, w_eco146913, w_eco146914, w_eco146915, w_eco146916, w_eco146917, w_eco146918, w_eco146919, w_eco146920, w_eco146921, w_eco146922, w_eco146923, w_eco146924, w_eco146925, w_eco146926, w_eco146927, w_eco146928, w_eco146929, w_eco146930, w_eco146931, w_eco146932, w_eco146933, w_eco146934, w_eco146935, w_eco146936, w_eco146937, w_eco146938, w_eco146939, w_eco146940, w_eco146941, w_eco146942, w_eco146943, w_eco146944, w_eco146945, w_eco146946, w_eco146947, w_eco146948, w_eco146949, w_eco146950, w_eco146951, w_eco146952, w_eco146953, w_eco146954, w_eco146955, w_eco146956, w_eco146957, w_eco146958, w_eco146959, w_eco146960, w_eco146961, w_eco146962, w_eco146963, w_eco146964, w_eco146965, w_eco146966, w_eco146967, w_eco146968, w_eco146969, w_eco146970, w_eco146971, w_eco146972, w_eco146973, w_eco146974, w_eco146975, w_eco146976, w_eco146977, w_eco146978, w_eco146979, w_eco146980, w_eco146981, w_eco146982, w_eco146983, w_eco146984, w_eco146985, w_eco146986, w_eco146987, w_eco146988, w_eco146989, w_eco146990, w_eco146991, w_eco146992, w_eco146993, w_eco146994, w_eco146995, w_eco146996, w_eco146997, w_eco146998, w_eco146999, w_eco147000, w_eco147001, w_eco147002, w_eco147003, w_eco147004, w_eco147005, w_eco147006, w_eco147007, w_eco147008, w_eco147009, w_eco147010, w_eco147011, w_eco147012, w_eco147013, w_eco147014, w_eco147015, w_eco147016, w_eco147017, w_eco147018, w_eco147019, w_eco147020, w_eco147021, w_eco147022, w_eco147023, w_eco147024, w_eco147025, w_eco147026, w_eco147027, w_eco147028, w_eco147029, w_eco147030, w_eco147031, w_eco147032, w_eco147033, w_eco147034, w_eco147035, w_eco147036, w_eco147037, w_eco147038, w_eco147039, w_eco147040, w_eco147041, w_eco147042, w_eco147043, w_eco147044, w_eco147045, w_eco147046, w_eco147047, w_eco147048, w_eco147049, w_eco147050, w_eco147051, w_eco147052, w_eco147053, w_eco147054, w_eco147055, w_eco147056, w_eco147057, w_eco147058, w_eco147059, w_eco147060, w_eco147061, w_eco147062, w_eco147063, w_eco147064, w_eco147065, w_eco147066, w_eco147067, w_eco147068, w_eco147069, w_eco147070, w_eco147071, w_eco147072, w_eco147073, w_eco147074, w_eco147075, w_eco147076, w_eco147077, w_eco147078, w_eco147079, w_eco147080, w_eco147081, w_eco147082, w_eco147083, w_eco147084, w_eco147085, w_eco147086, w_eco147087, w_eco147088, w_eco147089, w_eco147090, w_eco147091, w_eco147092, w_eco147093, w_eco147094, w_eco147095, w_eco147096, w_eco147097, w_eco147098, w_eco147099, w_eco147100, w_eco147101, w_eco147102, w_eco147103, w_eco147104, w_eco147105, w_eco147106, w_eco147107, w_eco147108, w_eco147109, w_eco147110, w_eco147111, w_eco147112, w_eco147113, w_eco147114, w_eco147115, w_eco147116, w_eco147117, w_eco147118, w_eco147119, w_eco147120, w_eco147121, w_eco147122, w_eco147123, w_eco147124, w_eco147125, w_eco147126, w_eco147127, w_eco147128, w_eco147129, w_eco147130, w_eco147131, w_eco147132, w_eco147133, w_eco147134, w_eco147135, w_eco147136, w_eco147137, w_eco147138, w_eco147139, w_eco147140, w_eco147141, w_eco147142, w_eco147143, w_eco147144, w_eco147145, w_eco147146, w_eco147147, w_eco147148, w_eco147149, w_eco147150, w_eco147151, w_eco147152, w_eco147153, w_eco147154, w_eco147155, w_eco147156, w_eco147157, w_eco147158, w_eco147159, w_eco147160, w_eco147161, w_eco147162, w_eco147163, w_eco147164, w_eco147165, w_eco147166, w_eco147167, w_eco147168, w_eco147169, w_eco147170, w_eco147171, w_eco147172, w_eco147173, w_eco147174, w_eco147175, w_eco147176, w_eco147177, w_eco147178, w_eco147179, w_eco147180, w_eco147181, w_eco147182, w_eco147183, w_eco147184, w_eco147185, w_eco147186, w_eco147187, w_eco147188, w_eco147189, w_eco147190, w_eco147191, w_eco147192, w_eco147193, w_eco147194, w_eco147195, w_eco147196, w_eco147197, w_eco147198, w_eco147199, w_eco147200, w_eco147201, w_eco147202, w_eco147203, w_eco147204, w_eco147205, w_eco147206, w_eco147207, w_eco147208, w_eco147209, w_eco147210, w_eco147211, w_eco147212, w_eco147213, w_eco147214, w_eco147215, w_eco147216, w_eco147217, w_eco147218, w_eco147219, w_eco147220, w_eco147221, w_eco147222, w_eco147223, w_eco147224, w_eco147225, w_eco147226, w_eco147227, w_eco147228, w_eco147229, w_eco147230, w_eco147231, w_eco147232, w_eco147233, w_eco147234, w_eco147235, w_eco147236, w_eco147237, w_eco147238, w_eco147239, w_eco147240, w_eco147241, w_eco147242, w_eco147243, w_eco147244, w_eco147245, w_eco147246, w_eco147247, w_eco147248, w_eco147249, w_eco147250, w_eco147251, w_eco147252, w_eco147253, w_eco147254, w_eco147255, w_eco147256, w_eco147257, w_eco147258, w_eco147259, w_eco147260, w_eco147261, w_eco147262, w_eco147263, w_eco147264, w_eco147265, w_eco147266, w_eco147267, w_eco147268, w_eco147269, w_eco147270, w_eco147271, w_eco147272, w_eco147273, w_eco147274, w_eco147275, w_eco147276, w_eco147277, w_eco147278, w_eco147279, w_eco147280, w_eco147281, w_eco147282, w_eco147283, w_eco147284, w_eco147285, w_eco147286, w_eco147287, w_eco147288, w_eco147289, w_eco147290, w_eco147291, w_eco147292, w_eco147293, w_eco147294, w_eco147295, w_eco147296, w_eco147297, w_eco147298, w_eco147299, w_eco147300, w_eco147301, w_eco147302, w_eco147303, w_eco147304, w_eco147305, w_eco147306, w_eco147307, w_eco147308, w_eco147309, w_eco147310, w_eco147311, w_eco147312, w_eco147313, w_eco147314, w_eco147315, w_eco147316, w_eco147317, w_eco147318, w_eco147319, w_eco147320, w_eco147321, w_eco147322, w_eco147323, w_eco147324, w_eco147325, w_eco147326, w_eco147327, w_eco147328, w_eco147329, w_eco147330, w_eco147331, w_eco147332, w_eco147333, w_eco147334, w_eco147335, w_eco147336, w_eco147337, w_eco147338, w_eco147339, w_eco147340, w_eco147341, w_eco147342, w_eco147343, w_eco147344, w_eco147345, w_eco147346, w_eco147347, w_eco147348, w_eco147349, w_eco147350, w_eco147351, w_eco147352, w_eco147353, w_eco147354, w_eco147355, w_eco147356, w_eco147357, w_eco147358, w_eco147359, w_eco147360, w_eco147361, w_eco147362, w_eco147363, w_eco147364, w_eco147365, w_eco147366, w_eco147367, w_eco147368, w_eco147369, w_eco147370, w_eco147371, w_eco147372, w_eco147373, w_eco147374, w_eco147375, w_eco147376, w_eco147377, w_eco147378, w_eco147379, w_eco147380, w_eco147381, w_eco147382, w_eco147383, w_eco147384, w_eco147385, w_eco147386, w_eco147387, w_eco147388, w_eco147389, w_eco147390, w_eco147391, w_eco147392, w_eco147393, w_eco147394, w_eco147395, w_eco147396, w_eco147397, w_eco147398, w_eco147399, w_eco147400, w_eco147401, w_eco147402, w_eco147403, w_eco147404, w_eco147405, w_eco147406, w_eco147407, w_eco147408, w_eco147409, w_eco147410, w_eco147411, w_eco147412, w_eco147413, w_eco147414, w_eco147415, w_eco147416, w_eco147417, w_eco147418, w_eco147419, w_eco147420, w_eco147421, w_eco147422, w_eco147423, w_eco147424, w_eco147425, w_eco147426, w_eco147427, w_eco147428, w_eco147429, w_eco147430, w_eco147431, w_eco147432, w_eco147433, w_eco147434, w_eco147435, w_eco147436, w_eco147437, w_eco147438, w_eco147439, w_eco147440, w_eco147441, w_eco147442, w_eco147443, w_eco147444, w_eco147445, w_eco147446, w_eco147447, w_eco147448, w_eco147449, w_eco147450, w_eco147451, w_eco147452, w_eco147453, w_eco147454, w_eco147455, w_eco147456, w_eco147457, w_eco147458, w_eco147459, w_eco147460, w_eco147461, w_eco147462, w_eco147463, w_eco147464, w_eco147465, w_eco147466, w_eco147467, w_eco147468, w_eco147469, w_eco147470, w_eco147471, w_eco147472, w_eco147473, w_eco147474, w_eco147475, w_eco147476, w_eco147477, w_eco147478, w_eco147479, w_eco147480, w_eco147481, w_eco147482, w_eco147483, w_eco147484, w_eco147485, w_eco147486, w_eco147487, w_eco147488, w_eco147489, w_eco147490, w_eco147491, w_eco147492, w_eco147493, w_eco147494, w_eco147495, w_eco147496, w_eco147497, w_eco147498, w_eco147499, w_eco147500, w_eco147501, w_eco147502, w_eco147503, w_eco147504, w_eco147505, w_eco147506, w_eco147507, w_eco147508, w_eco147509, w_eco147510, w_eco147511, w_eco147512, w_eco147513, w_eco147514, w_eco147515, w_eco147516, w_eco147517, w_eco147518, w_eco147519, w_eco147520, w_eco147521, w_eco147522, w_eco147523, w_eco147524, w_eco147525, w_eco147526, w_eco147527, w_eco147528, w_eco147529, w_eco147530, w_eco147531, w_eco147532, w_eco147533, w_eco147534, w_eco147535, w_eco147536, w_eco147537, w_eco147538, w_eco147539, w_eco147540, w_eco147541, w_eco147542, w_eco147543, w_eco147544, w_eco147545, w_eco147546, w_eco147547, w_eco147548, w_eco147549, w_eco147550, w_eco147551, w_eco147552, w_eco147553, w_eco147554, w_eco147555, w_eco147556, w_eco147557, w_eco147558, w_eco147559, w_eco147560, w_eco147561, w_eco147562, w_eco147563, w_eco147564, w_eco147565, w_eco147566, w_eco147567, w_eco147568, w_eco147569, w_eco147570, w_eco147571, w_eco147572, w_eco147573, w_eco147574, w_eco147575, w_eco147576, w_eco147577, w_eco147578, w_eco147579, w_eco147580, w_eco147581, w_eco147582, w_eco147583, w_eco147584, w_eco147585, w_eco147586, w_eco147587, w_eco147588, w_eco147589, w_eco147590, w_eco147591, w_eco147592, w_eco147593, w_eco147594, w_eco147595, w_eco147596, w_eco147597, w_eco147598, w_eco147599, w_eco147600, w_eco147601, w_eco147602, w_eco147603, w_eco147604, w_eco147605, w_eco147606, w_eco147607, w_eco147608, w_eco147609, w_eco147610, w_eco147611, w_eco147612, w_eco147613, w_eco147614, w_eco147615, w_eco147616, w_eco147617, w_eco147618, w_eco147619, w_eco147620, w_eco147621, w_eco147622, w_eco147623, w_eco147624, w_eco147625, w_eco147626, w_eco147627, w_eco147628, w_eco147629, w_eco147630, w_eco147631, w_eco147632, w_eco147633, w_eco147634, w_eco147635, w_eco147636, w_eco147637, w_eco147638, w_eco147639, w_eco147640, w_eco147641, w_eco147642, w_eco147643, w_eco147644, w_eco147645, w_eco147646, w_eco147647, w_eco147648, w_eco147649, w_eco147650, w_eco147651, w_eco147652, w_eco147653, w_eco147654, w_eco147655, w_eco147656, w_eco147657, w_eco147658, w_eco147659, w_eco147660, w_eco147661, w_eco147662, w_eco147663, w_eco147664, w_eco147665, w_eco147666, w_eco147667, w_eco147668, w_eco147669, w_eco147670, w_eco147671, w_eco147672, w_eco147673, w_eco147674, w_eco147675, w_eco147676, w_eco147677, w_eco147678, w_eco147679, w_eco147680, w_eco147681, w_eco147682, w_eco147683, w_eco147684, w_eco147685, w_eco147686, w_eco147687, w_eco147688, w_eco147689, w_eco147690, w_eco147691, w_eco147692, w_eco147693, w_eco147694, w_eco147695, w_eco147696, w_eco147697, w_eco147698, w_eco147699, w_eco147700, w_eco147701, w_eco147702, w_eco147703, w_eco147704, w_eco147705, w_eco147706, w_eco147707, w_eco147708, w_eco147709, w_eco147710, w_eco147711, w_eco147712, w_eco147713, w_eco147714, w_eco147715, w_eco147716, w_eco147717, w_eco147718, w_eco147719, w_eco147720, w_eco147721, w_eco147722, w_eco147723, w_eco147724, w_eco147725, w_eco147726, w_eco147727, w_eco147728, w_eco147729, w_eco147730, w_eco147731, w_eco147732, w_eco147733, w_eco147734, w_eco147735, w_eco147736, w_eco147737, w_eco147738, w_eco147739, w_eco147740, w_eco147741, w_eco147742, w_eco147743, w_eco147744, w_eco147745, w_eco147746, w_eco147747, w_eco147748, w_eco147749, w_eco147750, w_eco147751, w_eco147752, w_eco147753, w_eco147754, w_eco147755, w_eco147756, w_eco147757, w_eco147758, w_eco147759, w_eco147760, w_eco147761, w_eco147762, w_eco147763, w_eco147764, w_eco147765, w_eco147766, w_eco147767, w_eco147768, w_eco147769, w_eco147770, w_eco147771, w_eco147772, w_eco147773, w_eco147774, w_eco147775, w_eco147776, w_eco147777, w_eco147778, w_eco147779, w_eco147780, w_eco147781, w_eco147782, w_eco147783, w_eco147784, w_eco147785, w_eco147786, w_eco147787, w_eco147788, w_eco147789, w_eco147790, w_eco147791, w_eco147792, w_eco147793, w_eco147794, w_eco147795, w_eco147796, w_eco147797, w_eco147798, w_eco147799, w_eco147800, w_eco147801, w_eco147802, w_eco147803, w_eco147804, w_eco147805, w_eco147806, w_eco147807, w_eco147808, w_eco147809, w_eco147810, w_eco147811, w_eco147812, w_eco147813, w_eco147814, w_eco147815, w_eco147816, w_eco147817, w_eco147818, w_eco147819, w_eco147820, w_eco147821, w_eco147822, w_eco147823, w_eco147824, w_eco147825, w_eco147826, w_eco147827, w_eco147828, w_eco147829, w_eco147830, w_eco147831, w_eco147832, w_eco147833, w_eco147834, w_eco147835, w_eco147836, w_eco147837, w_eco147838, w_eco147839, w_eco147840, w_eco147841, w_eco147842, w_eco147843, w_eco147844, w_eco147845, w_eco147846, w_eco147847, w_eco147848, w_eco147849, w_eco147850, w_eco147851, w_eco147852, w_eco147853, w_eco147854, w_eco147855, w_eco147856, w_eco147857, w_eco147858, w_eco147859, w_eco147860, w_eco147861, w_eco147862, w_eco147863, w_eco147864, w_eco147865, w_eco147866, w_eco147867, w_eco147868, w_eco147869, w_eco147870, w_eco147871, w_eco147872, w_eco147873, w_eco147874, w_eco147875, w_eco147876, w_eco147877, w_eco147878, w_eco147879, w_eco147880, w_eco147881, w_eco147882, w_eco147883, w_eco147884, w_eco147885, w_eco147886, w_eco147887, w_eco147888, w_eco147889, w_eco147890, w_eco147891, w_eco147892, w_eco147893, w_eco147894, w_eco147895, w_eco147896, w_eco147897, w_eco147898, w_eco147899, w_eco147900, w_eco147901, w_eco147902, w_eco147903, w_eco147904, w_eco147905, w_eco147906, w_eco147907, w_eco147908, w_eco147909, w_eco147910, w_eco147911, w_eco147912, w_eco147913, w_eco147914, w_eco147915, w_eco147916, w_eco147917, w_eco147918, w_eco147919, w_eco147920, w_eco147921, w_eco147922, w_eco147923, w_eco147924, w_eco147925, w_eco147926, w_eco147927, w_eco147928, w_eco147929, w_eco147930, w_eco147931, w_eco147932, w_eco147933, w_eco147934, w_eco147935, w_eco147936, w_eco147937, w_eco147938, w_eco147939, w_eco147940, w_eco147941, w_eco147942, w_eco147943, w_eco147944, w_eco147945, w_eco147946, w_eco147947, w_eco147948, w_eco147949, w_eco147950, w_eco147951, w_eco147952, w_eco147953, w_eco147954, w_eco147955, w_eco147956, w_eco147957, w_eco147958, w_eco147959, w_eco147960, w_eco147961, w_eco147962, w_eco147963, w_eco147964, w_eco147965, w_eco147966, w_eco147967, w_eco147968, w_eco147969, w_eco147970, w_eco147971, w_eco147972, w_eco147973, w_eco147974, w_eco147975, w_eco147976, w_eco147977, w_eco147978, w_eco147979, w_eco147980, w_eco147981, w_eco147982, w_eco147983, w_eco147984, w_eco147985, w_eco147986, w_eco147987, w_eco147988, w_eco147989, w_eco147990, w_eco147991, w_eco147992, w_eco147993, w_eco147994, w_eco147995, w_eco147996, w_eco147997, w_eco147998, w_eco147999, w_eco148000, w_eco148001, w_eco148002, w_eco148003, w_eco148004, w_eco148005, w_eco148006, w_eco148007, w_eco148008, w_eco148009, w_eco148010, w_eco148011, w_eco148012, w_eco148013, w_eco148014, w_eco148015, w_eco148016, w_eco148017, w_eco148018, w_eco148019, w_eco148020, w_eco148021, w_eco148022, w_eco148023, w_eco148024, w_eco148025, w_eco148026, w_eco148027, w_eco148028, w_eco148029, w_eco148030, w_eco148031, w_eco148032, w_eco148033, w_eco148034, w_eco148035, w_eco148036, w_eco148037, w_eco148038, w_eco148039, w_eco148040, w_eco148041, w_eco148042, w_eco148043, w_eco148044, w_eco148045, w_eco148046, w_eco148047, w_eco148048, w_eco148049, w_eco148050, w_eco148051, w_eco148052, w_eco148053, w_eco148054, w_eco148055, w_eco148056, w_eco148057, w_eco148058, w_eco148059, w_eco148060, w_eco148061, w_eco148062, w_eco148063, w_eco148064, w_eco148065, w_eco148066, w_eco148067, w_eco148068, w_eco148069, w_eco148070, w_eco148071, w_eco148072, w_eco148073, w_eco148074, w_eco148075, w_eco148076, w_eco148077, w_eco148078, w_eco148079, w_eco148080, w_eco148081, w_eco148082, w_eco148083, w_eco148084, w_eco148085, w_eco148086, w_eco148087, w_eco148088, w_eco148089, w_eco148090, w_eco148091, w_eco148092, w_eco148093, w_eco148094, w_eco148095, w_eco148096, w_eco148097, w_eco148098, w_eco148099, w_eco148100, w_eco148101, w_eco148102, w_eco148103, w_eco148104, w_eco148105, w_eco148106, w_eco148107, w_eco148108, w_eco148109, w_eco148110, w_eco148111, w_eco148112, w_eco148113, w_eco148114, w_eco148115, w_eco148116, w_eco148117, w_eco148118, w_eco148119, w_eco148120, w_eco148121, w_eco148122, w_eco148123, w_eco148124, w_eco148125, w_eco148126, w_eco148127, w_eco148128, w_eco148129, w_eco148130, w_eco148131, w_eco148132, w_eco148133, w_eco148134, w_eco148135, w_eco148136, w_eco148137, w_eco148138, w_eco148139, w_eco148140, w_eco148141, w_eco148142, w_eco148143, w_eco148144, w_eco148145, w_eco148146, w_eco148147, w_eco148148, w_eco148149, w_eco148150, w_eco148151, w_eco148152, w_eco148153, w_eco148154, w_eco148155, w_eco148156, w_eco148157, w_eco148158, w_eco148159, w_eco148160, w_eco148161, w_eco148162, w_eco148163, w_eco148164, w_eco148165, w_eco148166, w_eco148167, w_eco148168, w_eco148169, w_eco148170, w_eco148171, w_eco148172, w_eco148173, w_eco148174, w_eco148175, w_eco148176, w_eco148177, w_eco148178, w_eco148179, w_eco148180, w_eco148181, w_eco148182, w_eco148183, w_eco148184, w_eco148185, w_eco148186, w_eco148187, w_eco148188, w_eco148189, w_eco148190, w_eco148191, w_eco148192, w_eco148193, w_eco148194, w_eco148195, w_eco148196, w_eco148197, w_eco148198, w_eco148199, w_eco148200, w_eco148201, w_eco148202, w_eco148203, w_eco148204, w_eco148205, w_eco148206, w_eco148207, w_eco148208, w_eco148209, w_eco148210, w_eco148211, w_eco148212, w_eco148213, w_eco148214, w_eco148215, w_eco148216, w_eco148217, w_eco148218, w_eco148219, w_eco148220, w_eco148221, w_eco148222, w_eco148223, w_eco148224, w_eco148225, w_eco148226, w_eco148227, w_eco148228, w_eco148229, w_eco148230, w_eco148231, w_eco148232, w_eco148233, w_eco148234, w_eco148235, w_eco148236, w_eco148237, w_eco148238, w_eco148239, w_eco148240, w_eco148241, w_eco148242, w_eco148243, w_eco148244, w_eco148245, w_eco148246, w_eco148247, w_eco148248, w_eco148249, w_eco148250, w_eco148251, w_eco148252, w_eco148253, w_eco148254, w_eco148255, w_eco148256, w_eco148257, w_eco148258, w_eco148259, w_eco148260, w_eco148261, w_eco148262, w_eco148263, w_eco148264, w_eco148265, w_eco148266, w_eco148267, w_eco148268, w_eco148269, w_eco148270, w_eco148271, w_eco148272, w_eco148273, w_eco148274, w_eco148275, w_eco148276, w_eco148277, w_eco148278, w_eco148279, w_eco148280, w_eco148281, w_eco148282, w_eco148283, w_eco148284, w_eco148285, w_eco148286, w_eco148287, w_eco148288, w_eco148289, w_eco148290, w_eco148291, w_eco148292, w_eco148293, w_eco148294, w_eco148295, w_eco148296, w_eco148297, w_eco148298, w_eco148299, w_eco148300, w_eco148301, w_eco148302, w_eco148303, w_eco148304, w_eco148305, w_eco148306, w_eco148307, w_eco148308, w_eco148309, w_eco148310, w_eco148311, w_eco148312, w_eco148313, w_eco148314, w_eco148315, w_eco148316, w_eco148317, w_eco148318, w_eco148319, w_eco148320, w_eco148321, w_eco148322, w_eco148323, w_eco148324, w_eco148325, w_eco148326, w_eco148327, w_eco148328, w_eco148329, w_eco148330, w_eco148331, w_eco148332, w_eco148333, w_eco148334, w_eco148335, w_eco148336, w_eco148337, w_eco148338, w_eco148339, w_eco148340, w_eco148341, w_eco148342, w_eco148343, w_eco148344, w_eco148345, w_eco148346, w_eco148347, w_eco148348, w_eco148349, w_eco148350, w_eco148351, w_eco148352, w_eco148353, w_eco148354, w_eco148355, w_eco148356, w_eco148357, w_eco148358, w_eco148359, w_eco148360, w_eco148361, w_eco148362, w_eco148363, w_eco148364, w_eco148365, w_eco148366, w_eco148367, w_eco148368, w_eco148369, w_eco148370, w_eco148371, w_eco148372, w_eco148373, w_eco148374, w_eco148375, w_eco148376, w_eco148377, w_eco148378, w_eco148379, w_eco148380, w_eco148381, w_eco148382, w_eco148383, w_eco148384, w_eco148385, w_eco148386, w_eco148387, w_eco148388, w_eco148389, w_eco148390, w_eco148391, w_eco148392, w_eco148393, w_eco148394, w_eco148395, w_eco148396, w_eco148397, w_eco148398, w_eco148399, w_eco148400, w_eco148401, w_eco148402, w_eco148403, w_eco148404, w_eco148405, w_eco148406, w_eco148407, w_eco148408, w_eco148409, w_eco148410, w_eco148411, w_eco148412, w_eco148413, w_eco148414, w_eco148415, w_eco148416, w_eco148417, w_eco148418, w_eco148419, w_eco148420, w_eco148421, w_eco148422, w_eco148423, w_eco148424, w_eco148425, w_eco148426, w_eco148427, w_eco148428, w_eco148429, w_eco148430, w_eco148431, w_eco148432, w_eco148433, w_eco148434, w_eco148435, w_eco148436, w_eco148437, w_eco148438, w_eco148439, w_eco148440, w_eco148441, w_eco148442, w_eco148443, w_eco148444, w_eco148445, w_eco148446, w_eco148447, w_eco148448, w_eco148449, w_eco148450, w_eco148451, w_eco148452, w_eco148453, w_eco148454, w_eco148455, w_eco148456, w_eco148457, w_eco148458, w_eco148459, w_eco148460, w_eco148461, w_eco148462, w_eco148463, w_eco148464, w_eco148465, w_eco148466, w_eco148467, w_eco148468, w_eco148469, w_eco148470, w_eco148471, w_eco148472, w_eco148473, w_eco148474, w_eco148475, w_eco148476, w_eco148477, w_eco148478, w_eco148479, w_eco148480, w_eco148481, w_eco148482, w_eco148483, w_eco148484, w_eco148485, w_eco148486, w_eco148487, w_eco148488, w_eco148489, w_eco148490, w_eco148491, w_eco148492, w_eco148493, w_eco148494, w_eco148495, w_eco148496, w_eco148497, w_eco148498, w_eco148499, w_eco148500, w_eco148501, w_eco148502, w_eco148503, w_eco148504, w_eco148505, w_eco148506, w_eco148507, w_eco148508, w_eco148509, w_eco148510, w_eco148511, w_eco148512, w_eco148513, w_eco148514, w_eco148515, w_eco148516, w_eco148517, w_eco148518, w_eco148519, w_eco148520, w_eco148521, w_eco148522, w_eco148523, w_eco148524, w_eco148525, w_eco148526, w_eco148527, w_eco148528, w_eco148529, w_eco148530, w_eco148531, w_eco148532, w_eco148533, w_eco148534, w_eco148535, w_eco148536, w_eco148537, w_eco148538, w_eco148539, w_eco148540, w_eco148541, w_eco148542, w_eco148543, w_eco148544, w_eco148545, w_eco148546, w_eco148547, w_eco148548, w_eco148549, w_eco148550, w_eco148551, w_eco148552, w_eco148553, w_eco148554, w_eco148555, w_eco148556, w_eco148557, w_eco148558, w_eco148559, w_eco148560, w_eco148561, w_eco148562, w_eco148563, w_eco148564, w_eco148565, w_eco148566, w_eco148567, w_eco148568, w_eco148569, w_eco148570, w_eco148571, w_eco148572, w_eco148573, w_eco148574, w_eco148575, w_eco148576, w_eco148577, w_eco148578, w_eco148579, w_eco148580, w_eco148581, w_eco148582, w_eco148583, w_eco148584, w_eco148585, w_eco148586, w_eco148587, w_eco148588, w_eco148589, w_eco148590, w_eco148591, w_eco148592, w_eco148593, w_eco148594, w_eco148595, w_eco148596, w_eco148597, w_eco148598, w_eco148599, w_eco148600, w_eco148601, w_eco148602, w_eco148603, w_eco148604, w_eco148605, w_eco148606, w_eco148607, w_eco148608, w_eco148609, w_eco148610, w_eco148611, w_eco148612, w_eco148613, w_eco148614, w_eco148615, w_eco148616, w_eco148617, w_eco148618, w_eco148619, w_eco148620, w_eco148621, w_eco148622, w_eco148623, w_eco148624, w_eco148625, w_eco148626, w_eco148627, w_eco148628, w_eco148629, w_eco148630, w_eco148631, w_eco148632, w_eco148633, w_eco148634, w_eco148635, w_eco148636, w_eco148637, w_eco148638, w_eco148639, w_eco148640, w_eco148641, w_eco148642, w_eco148643, w_eco148644, w_eco148645, w_eco148646, w_eco148647, w_eco148648, w_eco148649, w_eco148650, w_eco148651, w_eco148652, w_eco148653, w_eco148654, w_eco148655, w_eco148656, w_eco148657, w_eco148658, w_eco148659, w_eco148660, w_eco148661, w_eco148662, w_eco148663, w_eco148664, w_eco148665, w_eco148666, w_eco148667, w_eco148668, w_eco148669, w_eco148670, w_eco148671, w_eco148672, w_eco148673, w_eco148674, w_eco148675, w_eco148676, w_eco148677, w_eco148678, w_eco148679, w_eco148680, w_eco148681, w_eco148682, w_eco148683, w_eco148684, w_eco148685, w_eco148686, w_eco148687, w_eco148688, w_eco148689, w_eco148690, w_eco148691, w_eco148692, w_eco148693, w_eco148694, w_eco148695, w_eco148696, w_eco148697, w_eco148698, w_eco148699, w_eco148700, w_eco148701, w_eco148702, w_eco148703, w_eco148704, w_eco148705, w_eco148706, w_eco148707, w_eco148708, w_eco148709, w_eco148710, w_eco148711, w_eco148712, w_eco148713, w_eco148714, w_eco148715, w_eco148716, w_eco148717, w_eco148718, w_eco148719, w_eco148720, w_eco148721, w_eco148722, w_eco148723, w_eco148724, w_eco148725, w_eco148726, w_eco148727, w_eco148728, w_eco148729, w_eco148730, w_eco148731, w_eco148732, w_eco148733, w_eco148734, w_eco148735, w_eco148736, w_eco148737, w_eco148738, w_eco148739, w_eco148740, w_eco148741, w_eco148742, w_eco148743, w_eco148744, w_eco148745, w_eco148746, w_eco148747, w_eco148748, w_eco148749, w_eco148750, w_eco148751, w_eco148752, w_eco148753, w_eco148754, w_eco148755, w_eco148756, w_eco148757, w_eco148758, w_eco148759, w_eco148760, w_eco148761, w_eco148762, w_eco148763, w_eco148764, w_eco148765, w_eco148766, w_eco148767, w_eco148768, w_eco148769, w_eco148770, w_eco148771, w_eco148772, w_eco148773, w_eco148774, w_eco148775, w_eco148776, w_eco148777, w_eco148778, w_eco148779, w_eco148780, w_eco148781, w_eco148782, w_eco148783, w_eco148784, w_eco148785, w_eco148786, w_eco148787, w_eco148788, w_eco148789, w_eco148790, w_eco148791, w_eco148792, w_eco148793, w_eco148794, w_eco148795, w_eco148796, w_eco148797, w_eco148798, w_eco148799, w_eco148800, w_eco148801, w_eco148802, w_eco148803, w_eco148804, w_eco148805, w_eco148806, w_eco148807, w_eco148808, w_eco148809, w_eco148810, w_eco148811, w_eco148812, w_eco148813, w_eco148814, w_eco148815, w_eco148816, w_eco148817, w_eco148818, w_eco148819, w_eco148820, w_eco148821, w_eco148822, w_eco148823, w_eco148824, w_eco148825, w_eco148826, w_eco148827, w_eco148828, w_eco148829, w_eco148830, w_eco148831, w_eco148832, w_eco148833, w_eco148834, w_eco148835, w_eco148836, w_eco148837, w_eco148838, w_eco148839, w_eco148840, w_eco148841, w_eco148842, w_eco148843, w_eco148844, w_eco148845, w_eco148846, w_eco148847, w_eco148848, w_eco148849, w_eco148850, w_eco148851, w_eco148852, w_eco148853, w_eco148854, w_eco148855, w_eco148856, w_eco148857, w_eco148858, w_eco148859, w_eco148860, w_eco148861, w_eco148862, w_eco148863, w_eco148864, w_eco148865, w_eco148866, w_eco148867, w_eco148868, w_eco148869, w_eco148870, w_eco148871, w_eco148872, w_eco148873, w_eco148874, w_eco148875, w_eco148876, w_eco148877, w_eco148878, w_eco148879, w_eco148880, w_eco148881, w_eco148882, w_eco148883, w_eco148884, w_eco148885, w_eco148886, w_eco148887, w_eco148888, w_eco148889, w_eco148890, w_eco148891, w_eco148892, w_eco148893, w_eco148894, w_eco148895, w_eco148896, w_eco148897, w_eco148898, w_eco148899, w_eco148900, w_eco148901, w_eco148902, w_eco148903, w_eco148904, w_eco148905, w_eco148906, w_eco148907, w_eco148908, w_eco148909, w_eco148910, w_eco148911, w_eco148912, w_eco148913, w_eco148914, w_eco148915, w_eco148916, w_eco148917, w_eco148918, w_eco148919, w_eco148920, w_eco148921, w_eco148922, w_eco148923, w_eco148924, w_eco148925, w_eco148926, w_eco148927, w_eco148928, w_eco148929, w_eco148930, w_eco148931, w_eco148932, w_eco148933, w_eco148934, w_eco148935, w_eco148936, w_eco148937, w_eco148938, w_eco148939, w_eco148940, w_eco148941, w_eco148942, w_eco148943, w_eco148944, w_eco148945, w_eco148946, w_eco148947, w_eco148948, w_eco148949, w_eco148950, w_eco148951, w_eco148952, w_eco148953, w_eco148954, w_eco148955, w_eco148956, w_eco148957, w_eco148958, w_eco148959, w_eco148960, w_eco148961, w_eco148962, w_eco148963, w_eco148964, w_eco148965, w_eco148966, w_eco148967, w_eco148968, w_eco148969, w_eco148970, w_eco148971, w_eco148972, w_eco148973, w_eco148974, w_eco148975, w_eco148976, w_eco148977, w_eco148978, w_eco148979, w_eco148980, w_eco148981, w_eco148982, w_eco148983, w_eco148984, w_eco148985, w_eco148986, w_eco148987, w_eco148988, w_eco148989, w_eco148990, w_eco148991, w_eco148992, w_eco148993, w_eco148994, w_eco148995, w_eco148996, w_eco148997, w_eco148998, w_eco148999, w_eco149000, w_eco149001, w_eco149002, w_eco149003, w_eco149004, w_eco149005, w_eco149006, w_eco149007, w_eco149008, w_eco149009, w_eco149010, w_eco149011, w_eco149012, w_eco149013, w_eco149014, w_eco149015, w_eco149016, w_eco149017, w_eco149018, w_eco149019, w_eco149020, w_eco149021, w_eco149022, w_eco149023, w_eco149024, w_eco149025, w_eco149026, w_eco149027, w_eco149028, w_eco149029, w_eco149030, w_eco149031, w_eco149032, w_eco149033, w_eco149034, w_eco149035, w_eco149036, w_eco149037, w_eco149038, w_eco149039, w_eco149040, w_eco149041, w_eco149042, w_eco149043, w_eco149044, w_eco149045, w_eco149046, w_eco149047, w_eco149048, w_eco149049, w_eco149050, w_eco149051, w_eco149052, w_eco149053, w_eco149054, w_eco149055, w_eco149056, w_eco149057, w_eco149058, w_eco149059, w_eco149060, w_eco149061, w_eco149062, w_eco149063, w_eco149064, w_eco149065, w_eco149066, w_eco149067, w_eco149068, w_eco149069, w_eco149070, w_eco149071, w_eco149072, w_eco149073, w_eco149074, w_eco149075, w_eco149076, w_eco149077, w_eco149078, w_eco149079, w_eco149080, w_eco149081, w_eco149082, w_eco149083, w_eco149084, w_eco149085, w_eco149086, w_eco149087, w_eco149088, w_eco149089, w_eco149090, w_eco149091, w_eco149092, w_eco149093, w_eco149094, w_eco149095, w_eco149096, w_eco149097, w_eco149098, w_eco149099, w_eco149100, w_eco149101, w_eco149102, w_eco149103, w_eco149104, w_eco149105, w_eco149106, w_eco149107, w_eco149108, w_eco149109, w_eco149110, w_eco149111, w_eco149112, w_eco149113, w_eco149114, w_eco149115, w_eco149116, w_eco149117, w_eco149118, w_eco149119, w_eco149120, w_eco149121, w_eco149122, w_eco149123, w_eco149124, w_eco149125, w_eco149126, w_eco149127, w_eco149128, w_eco149129, w_eco149130, w_eco149131, w_eco149132, w_eco149133, w_eco149134, w_eco149135, w_eco149136, w_eco149137, w_eco149138, w_eco149139, w_eco149140, w_eco149141, w_eco149142, w_eco149143, w_eco149144, w_eco149145, w_eco149146, w_eco149147, w_eco149148, w_eco149149, w_eco149150, w_eco149151, w_eco149152, w_eco149153, w_eco149154, w_eco149155, w_eco149156, w_eco149157, w_eco149158, w_eco149159, w_eco149160, w_eco149161, w_eco149162, w_eco149163, w_eco149164, w_eco149165, w_eco149166, w_eco149167, w_eco149168, w_eco149169, w_eco149170, w_eco149171, w_eco149172, w_eco149173, w_eco149174, w_eco149175, w_eco149176, w_eco149177, w_eco149178, w_eco149179, w_eco149180, w_eco149181, w_eco149182, w_eco149183, w_eco149184, w_eco149185, w_eco149186, w_eco149187, w_eco149188, w_eco149189, w_eco149190, w_eco149191, w_eco149192, w_eco149193, w_eco149194, w_eco149195, w_eco149196, w_eco149197, w_eco149198, w_eco149199, w_eco149200, w_eco149201, w_eco149202, w_eco149203, w_eco149204, w_eco149205, w_eco149206, w_eco149207, w_eco149208, w_eco149209, w_eco149210, w_eco149211, w_eco149212, w_eco149213, w_eco149214, w_eco149215, w_eco149216, w_eco149217, w_eco149218, w_eco149219, w_eco149220, w_eco149221, w_eco149222, w_eco149223, w_eco149224, w_eco149225, w_eco149226, w_eco149227, w_eco149228, w_eco149229, w_eco149230, w_eco149231, w_eco149232, w_eco149233, w_eco149234, w_eco149235, w_eco149236, w_eco149237, w_eco149238, w_eco149239, w_eco149240, w_eco149241, w_eco149242, w_eco149243, w_eco149244, w_eco149245, w_eco149246, w_eco149247, w_eco149248, w_eco149249, w_eco149250, w_eco149251, w_eco149252, w_eco149253, w_eco149254, w_eco149255, w_eco149256, w_eco149257, w_eco149258, w_eco149259, w_eco149260, w_eco149261, w_eco149262, w_eco149263, w_eco149264, w_eco149265, w_eco149266, w_eco149267, w_eco149268, w_eco149269, w_eco149270, w_eco149271, w_eco149272, w_eco149273, w_eco149274, w_eco149275, w_eco149276, w_eco149277, w_eco149278, w_eco149279, w_eco149280, w_eco149281, w_eco149282, w_eco149283, w_eco149284, w_eco149285, w_eco149286, w_eco149287, w_eco149288, w_eco149289, w_eco149290, w_eco149291, w_eco149292, w_eco149293, w_eco149294, w_eco149295, w_eco149296, w_eco149297, w_eco149298, w_eco149299, w_eco149300, w_eco149301, w_eco149302, w_eco149303, w_eco149304, w_eco149305, w_eco149306, w_eco149307, w_eco149308, w_eco149309, w_eco149310, w_eco149311, w_eco149312, w_eco149313, w_eco149314, w_eco149315, w_eco149316, w_eco149317, w_eco149318, w_eco149319, w_eco149320, w_eco149321, w_eco149322, w_eco149323, w_eco149324, w_eco149325, w_eco149326, w_eco149327, w_eco149328, w_eco149329, w_eco149330, w_eco149331, w_eco149332, w_eco149333, w_eco149334, w_eco149335, w_eco149336, w_eco149337, w_eco149338, w_eco149339, w_eco149340, w_eco149341, w_eco149342, w_eco149343, w_eco149344, w_eco149345, w_eco149346, w_eco149347, w_eco149348, w_eco149349, w_eco149350, w_eco149351, w_eco149352, w_eco149353, w_eco149354, w_eco149355, w_eco149356, w_eco149357, w_eco149358, w_eco149359, w_eco149360, w_eco149361, w_eco149362, w_eco149363, w_eco149364, w_eco149365, w_eco149366, w_eco149367, w_eco149368, w_eco149369, w_eco149370, w_eco149371, w_eco149372, w_eco149373, w_eco149374, w_eco149375, w_eco149376, w_eco149377, w_eco149378, w_eco149379, w_eco149380, w_eco149381, w_eco149382, w_eco149383, w_eco149384, w_eco149385, w_eco149386, w_eco149387, w_eco149388, w_eco149389, w_eco149390, w_eco149391, w_eco149392, w_eco149393, w_eco149394, w_eco149395, w_eco149396, w_eco149397, w_eco149398, w_eco149399, w_eco149400, w_eco149401, w_eco149402, w_eco149403, w_eco149404, w_eco149405, w_eco149406, w_eco149407, w_eco149408, w_eco149409, w_eco149410, w_eco149411, w_eco149412, w_eco149413, w_eco149414, w_eco149415, w_eco149416, w_eco149417, w_eco149418, w_eco149419, w_eco149420, w_eco149421, w_eco149422, w_eco149423, w_eco149424, w_eco149425, w_eco149426, w_eco149427, w_eco149428, w_eco149429, w_eco149430, w_eco149431, w_eco149432, w_eco149433, w_eco149434, w_eco149435, w_eco149436, w_eco149437, w_eco149438, w_eco149439, w_eco149440, w_eco149441, w_eco149442, w_eco149443, w_eco149444, w_eco149445, w_eco149446, w_eco149447, w_eco149448, w_eco149449, w_eco149450, w_eco149451, w_eco149452, w_eco149453, w_eco149454, w_eco149455, w_eco149456, w_eco149457, w_eco149458, w_eco149459, w_eco149460, w_eco149461, w_eco149462, w_eco149463, w_eco149464, w_eco149465, w_eco149466, w_eco149467, w_eco149468, w_eco149469, w_eco149470, w_eco149471, w_eco149472, w_eco149473, w_eco149474, w_eco149475, w_eco149476, w_eco149477, w_eco149478, w_eco149479, w_eco149480, w_eco149481, w_eco149482, w_eco149483, w_eco149484, w_eco149485, w_eco149486, w_eco149487, w_eco149488, w_eco149489, w_eco149490, w_eco149491, w_eco149492, w_eco149493, w_eco149494, w_eco149495, w_eco149496, w_eco149497, w_eco149498, w_eco149499, w_eco149500, w_eco149501, w_eco149502, w_eco149503, w_eco149504, w_eco149505, w_eco149506, w_eco149507, w_eco149508, w_eco149509, w_eco149510, w_eco149511, w_eco149512, w_eco149513, w_eco149514, w_eco149515, w_eco149516, w_eco149517, w_eco149518, w_eco149519, w_eco149520, w_eco149521, w_eco149522, w_eco149523, w_eco149524, w_eco149525, w_eco149526, w_eco149527, w_eco149528, w_eco149529, w_eco149530, w_eco149531, w_eco149532, w_eco149533, w_eco149534, w_eco149535, w_eco149536, w_eco149537, w_eco149538, w_eco149539, w_eco149540, w_eco149541, w_eco149542, w_eco149543, w_eco149544, w_eco149545, w_eco149546, w_eco149547, w_eco149548, w_eco149549, w_eco149550, w_eco149551, w_eco149552, w_eco149553, w_eco149554, w_eco149555, w_eco149556, w_eco149557, w_eco149558, w_eco149559, w_eco149560, w_eco149561, w_eco149562, w_eco149563, w_eco149564, w_eco149565, w_eco149566, w_eco149567, w_eco149568, w_eco149569, w_eco149570, w_eco149571, w_eco149572, w_eco149573, w_eco149574, w_eco149575, w_eco149576, w_eco149577, w_eco149578, w_eco149579, w_eco149580, w_eco149581, w_eco149582, w_eco149583, w_eco149584, w_eco149585, w_eco149586, w_eco149587, w_eco149588, w_eco149589, w_eco149590, w_eco149591, w_eco149592, w_eco149593, w_eco149594, w_eco149595, w_eco149596, w_eco149597, w_eco149598, w_eco149599, w_eco149600, w_eco149601, w_eco149602, w_eco149603, w_eco149604, w_eco149605, w_eco149606, w_eco149607, w_eco149608, w_eco149609, w_eco149610, w_eco149611, w_eco149612, w_eco149613, w_eco149614, w_eco149615, w_eco149616, w_eco149617, w_eco149618, w_eco149619, w_eco149620, w_eco149621, w_eco149622, w_eco149623, w_eco149624, w_eco149625, w_eco149626, w_eco149627, w_eco149628, w_eco149629, w_eco149630, w_eco149631, w_eco149632, w_eco149633, w_eco149634, w_eco149635, w_eco149636, w_eco149637, w_eco149638, w_eco149639, w_eco149640, w_eco149641, w_eco149642, w_eco149643, w_eco149644, w_eco149645, w_eco149646, w_eco149647, w_eco149648, w_eco149649, w_eco149650, w_eco149651, w_eco149652, w_eco149653, w_eco149654, w_eco149655, w_eco149656, w_eco149657, w_eco149658, w_eco149659, w_eco149660, w_eco149661, w_eco149662, w_eco149663, w_eco149664, w_eco149665, w_eco149666, w_eco149667, w_eco149668, w_eco149669, w_eco149670, w_eco149671, w_eco149672, w_eco149673, w_eco149674, w_eco149675, w_eco149676, w_eco149677, w_eco149678, w_eco149679, w_eco149680, w_eco149681, w_eco149682, w_eco149683, w_eco149684, w_eco149685, w_eco149686, w_eco149687, w_eco149688, w_eco149689, w_eco149690, w_eco149691, w_eco149692, w_eco149693, w_eco149694, w_eco149695, w_eco149696, w_eco149697, w_eco149698, w_eco149699, w_eco149700, w_eco149701, w_eco149702, w_eco149703, w_eco149704, w_eco149705, w_eco149706, w_eco149707, w_eco149708, w_eco149709, w_eco149710, w_eco149711, w_eco149712, w_eco149713, w_eco149714, w_eco149715, w_eco149716, w_eco149717, w_eco149718, w_eco149719, w_eco149720, w_eco149721, w_eco149722, w_eco149723, w_eco149724, w_eco149725, w_eco149726, w_eco149727, w_eco149728, w_eco149729, w_eco149730, w_eco149731, w_eco149732, w_eco149733, w_eco149734, w_eco149735, w_eco149736, w_eco149737, w_eco149738, w_eco149739, w_eco149740, w_eco149741, w_eco149742, w_eco149743, w_eco149744, w_eco149745, w_eco149746, w_eco149747, w_eco149748, w_eco149749, w_eco149750, w_eco149751, w_eco149752, w_eco149753, w_eco149754, w_eco149755, w_eco149756, w_eco149757, w_eco149758, w_eco149759, w_eco149760, w_eco149761, w_eco149762, w_eco149763, w_eco149764, w_eco149765, w_eco149766, w_eco149767, w_eco149768, w_eco149769, w_eco149770, w_eco149771, w_eco149772, w_eco149773, w_eco149774, w_eco149775, w_eco149776, w_eco149777, w_eco149778, w_eco149779, w_eco149780, w_eco149781, w_eco149782, w_eco149783, w_eco149784, w_eco149785, w_eco149786, w_eco149787, w_eco149788, w_eco149789, w_eco149790, w_eco149791, w_eco149792, w_eco149793, w_eco149794, w_eco149795, w_eco149796, w_eco149797, w_eco149798, w_eco149799, w_eco149800, w_eco149801, w_eco149802, w_eco149803, w_eco149804, w_eco149805, w_eco149806, w_eco149807, w_eco149808, w_eco149809, w_eco149810, w_eco149811, w_eco149812, w_eco149813, w_eco149814, w_eco149815, w_eco149816, w_eco149817, w_eco149818, w_eco149819, w_eco149820, w_eco149821, w_eco149822, w_eco149823, w_eco149824, w_eco149825, w_eco149826, w_eco149827, w_eco149828, w_eco149829, w_eco149830, w_eco149831, w_eco149832, w_eco149833, w_eco149834, w_eco149835, w_eco149836, w_eco149837, w_eco149838, w_eco149839, w_eco149840, w_eco149841, w_eco149842, w_eco149843, w_eco149844, w_eco149845, w_eco149846, w_eco149847, w_eco149848, w_eco149849, w_eco149850, w_eco149851, w_eco149852, w_eco149853, w_eco149854, w_eco149855, w_eco149856, w_eco149857, w_eco149858, w_eco149859, w_eco149860, w_eco149861, w_eco149862, w_eco149863, w_eco149864, w_eco149865, w_eco149866, w_eco149867, w_eco149868, w_eco149869, w_eco149870, w_eco149871, w_eco149872, w_eco149873, w_eco149874, w_eco149875, w_eco149876, w_eco149877, w_eco149878, w_eco149879, w_eco149880, w_eco149881, w_eco149882, w_eco149883, w_eco149884, w_eco149885, w_eco149886, w_eco149887, w_eco149888, w_eco149889, w_eco149890, w_eco149891, w_eco149892, w_eco149893, w_eco149894, w_eco149895, w_eco149896, w_eco149897, w_eco149898, w_eco149899, w_eco149900, w_eco149901, w_eco149902, w_eco149903, w_eco149904, w_eco149905, w_eco149906, w_eco149907, w_eco149908, w_eco149909, w_eco149910, w_eco149911, w_eco149912, w_eco149913, w_eco149914, w_eco149915, w_eco149916, w_eco149917, w_eco149918, w_eco149919, w_eco149920, w_eco149921, w_eco149922, w_eco149923, w_eco149924, w_eco149925, w_eco149926, w_eco149927, w_eco149928, w_eco149929, w_eco149930, w_eco149931, w_eco149932, w_eco149933, w_eco149934, w_eco149935, w_eco149936, w_eco149937, w_eco149938, w_eco149939, w_eco149940, w_eco149941, w_eco149942, w_eco149943, w_eco149944, w_eco149945, w_eco149946, w_eco149947, w_eco149948, w_eco149949, w_eco149950, w_eco149951, w_eco149952, w_eco149953, w_eco149954, w_eco149955, w_eco149956, w_eco149957, w_eco149958, w_eco149959, w_eco149960, w_eco149961, w_eco149962, w_eco149963, w_eco149964, w_eco149965, w_eco149966, w_eco149967, w_eco149968, w_eco149969, w_eco149970, w_eco149971, w_eco149972, w_eco149973, w_eco149974, w_eco149975, w_eco149976, w_eco149977, w_eco149978, w_eco149979, w_eco149980, w_eco149981, w_eco149982, w_eco149983, w_eco149984, w_eco149985, w_eco149986, w_eco149987, w_eco149988, w_eco149989, w_eco149990, w_eco149991, w_eco149992, w_eco149993, w_eco149994, w_eco149995, w_eco149996, w_eco149997, w_eco149998, w_eco149999, w_eco150000, w_eco150001, w_eco150002, w_eco150003, w_eco150004, w_eco150005, w_eco150006, w_eco150007, w_eco150008, w_eco150009, w_eco150010, w_eco150011, w_eco150012, w_eco150013, w_eco150014, w_eco150015, w_eco150016, w_eco150017, w_eco150018, w_eco150019, w_eco150020, w_eco150021, w_eco150022, w_eco150023, w_eco150024, w_eco150025, w_eco150026, w_eco150027, w_eco150028, w_eco150029, w_eco150030, w_eco150031, w_eco150032, w_eco150033, w_eco150034, w_eco150035, w_eco150036, w_eco150037, w_eco150038, w_eco150039, w_eco150040, w_eco150041, w_eco150042, w_eco150043, w_eco150044, w_eco150045, w_eco150046, w_eco150047, w_eco150048, w_eco150049, w_eco150050, w_eco150051, w_eco150052, w_eco150053, w_eco150054, w_eco150055, w_eco150056, w_eco150057, w_eco150058, w_eco150059, w_eco150060, w_eco150061, w_eco150062, w_eco150063, w_eco150064, w_eco150065, w_eco150066, w_eco150067, w_eco150068, w_eco150069, w_eco150070, w_eco150071, w_eco150072, w_eco150073, w_eco150074, w_eco150075, w_eco150076, w_eco150077, w_eco150078, w_eco150079, w_eco150080, w_eco150081, w_eco150082, w_eco150083, w_eco150084, w_eco150085, w_eco150086, w_eco150087, w_eco150088, w_eco150089, w_eco150090, w_eco150091, w_eco150092, w_eco150093, w_eco150094, w_eco150095, w_eco150096, w_eco150097, w_eco150098, w_eco150099, w_eco150100, w_eco150101, w_eco150102, w_eco150103, w_eco150104, w_eco150105, w_eco150106, w_eco150107, w_eco150108, w_eco150109, w_eco150110, w_eco150111, w_eco150112, w_eco150113, w_eco150114, w_eco150115, w_eco150116, w_eco150117, w_eco150118, w_eco150119, w_eco150120, w_eco150121, w_eco150122, w_eco150123, w_eco150124, w_eco150125, w_eco150126, w_eco150127, w_eco150128, w_eco150129, w_eco150130, w_eco150131, w_eco150132, w_eco150133, w_eco150134, w_eco150135, w_eco150136, w_eco150137, w_eco150138, w_eco150139, w_eco150140, w_eco150141, w_eco150142, w_eco150143, w_eco150144, w_eco150145, w_eco150146, w_eco150147, w_eco150148, w_eco150149, w_eco150150, w_eco150151, w_eco150152, w_eco150153, w_eco150154, w_eco150155, w_eco150156, w_eco150157, w_eco150158, w_eco150159, w_eco150160, w_eco150161, w_eco150162, w_eco150163, w_eco150164, w_eco150165, w_eco150166, w_eco150167, w_eco150168, w_eco150169, w_eco150170, w_eco150171, w_eco150172, w_eco150173, w_eco150174, w_eco150175, w_eco150176, w_eco150177, w_eco150178, w_eco150179, w_eco150180, w_eco150181, w_eco150182, w_eco150183, w_eco150184, w_eco150185, w_eco150186, w_eco150187, w_eco150188, w_eco150189, w_eco150190, w_eco150191, w_eco150192, w_eco150193, w_eco150194, w_eco150195, w_eco150196, w_eco150197, w_eco150198, w_eco150199, w_eco150200, w_eco150201, w_eco150202, w_eco150203, w_eco150204, w_eco150205, w_eco150206, w_eco150207, w_eco150208, w_eco150209, w_eco150210, w_eco150211, w_eco150212, w_eco150213, w_eco150214, w_eco150215, w_eco150216, w_eco150217, w_eco150218, w_eco150219, w_eco150220, w_eco150221, w_eco150222, w_eco150223, w_eco150224, w_eco150225, w_eco150226, w_eco150227, w_eco150228, w_eco150229, w_eco150230, w_eco150231, w_eco150232, w_eco150233, w_eco150234, w_eco150235, w_eco150236, w_eco150237, w_eco150238, w_eco150239, w_eco150240, w_eco150241, w_eco150242, w_eco150243, w_eco150244, w_eco150245, w_eco150246, w_eco150247, w_eco150248, w_eco150249, w_eco150250, w_eco150251, w_eco150252, w_eco150253, w_eco150254, w_eco150255, w_eco150256, w_eco150257, w_eco150258, w_eco150259, w_eco150260, w_eco150261, w_eco150262, w_eco150263, w_eco150264, w_eco150265, w_eco150266, w_eco150267, w_eco150268, w_eco150269, w_eco150270, w_eco150271, w_eco150272, w_eco150273, w_eco150274, w_eco150275, w_eco150276, w_eco150277, w_eco150278, w_eco150279, w_eco150280, w_eco150281, w_eco150282, w_eco150283, w_eco150284, w_eco150285, w_eco150286, w_eco150287, w_eco150288, w_eco150289, w_eco150290, w_eco150291, w_eco150292, w_eco150293, w_eco150294, w_eco150295, w_eco150296, w_eco150297, w_eco150298, w_eco150299, w_eco150300, w_eco150301, w_eco150302, w_eco150303, w_eco150304, w_eco150305, w_eco150306, w_eco150307, w_eco150308, w_eco150309, w_eco150310, w_eco150311, w_eco150312, w_eco150313, w_eco150314, w_eco150315, w_eco150316, w_eco150317, w_eco150318, w_eco150319, w_eco150320, w_eco150321, w_eco150322, w_eco150323, w_eco150324, w_eco150325, w_eco150326, w_eco150327, w_eco150328, w_eco150329, w_eco150330, w_eco150331, w_eco150332, w_eco150333, w_eco150334, w_eco150335, w_eco150336, w_eco150337, w_eco150338, w_eco150339, w_eco150340, w_eco150341, w_eco150342, w_eco150343, w_eco150344, w_eco150345, w_eco150346, w_eco150347, w_eco150348, w_eco150349, w_eco150350, w_eco150351, w_eco150352, w_eco150353, w_eco150354, w_eco150355, w_eco150356, w_eco150357, w_eco150358, w_eco150359, w_eco150360, w_eco150361, w_eco150362, w_eco150363, w_eco150364, w_eco150365, w_eco150366, w_eco150367, w_eco150368, w_eco150369, w_eco150370, w_eco150371, w_eco150372, w_eco150373, w_eco150374, w_eco150375, w_eco150376, w_eco150377, w_eco150378, w_eco150379, w_eco150380, w_eco150381, w_eco150382, w_eco150383, w_eco150384, w_eco150385, w_eco150386, w_eco150387, w_eco150388, w_eco150389, w_eco150390, w_eco150391, w_eco150392, w_eco150393, w_eco150394, w_eco150395, w_eco150396, w_eco150397, w_eco150398, w_eco150399, w_eco150400, w_eco150401, w_eco150402, w_eco150403, w_eco150404, w_eco150405, w_eco150406, w_eco150407, w_eco150408, w_eco150409, w_eco150410, w_eco150411, w_eco150412, w_eco150413, w_eco150414, w_eco150415, w_eco150416, w_eco150417, w_eco150418, w_eco150419, w_eco150420, w_eco150421, w_eco150422, w_eco150423, w_eco150424, w_eco150425, w_eco150426, w_eco150427, w_eco150428, w_eco150429, w_eco150430, w_eco150431, w_eco150432, w_eco150433, w_eco150434, w_eco150435, w_eco150436, w_eco150437, w_eco150438, w_eco150439, w_eco150440, w_eco150441, w_eco150442, w_eco150443, w_eco150444, w_eco150445, w_eco150446, w_eco150447, w_eco150448, w_eco150449, w_eco150450, w_eco150451, w_eco150452, w_eco150453, w_eco150454, w_eco150455, w_eco150456, w_eco150457, w_eco150458, w_eco150459, w_eco150460, w_eco150461, w_eco150462, w_eco150463, w_eco150464, w_eco150465, w_eco150466, w_eco150467, w_eco150468, w_eco150469, w_eco150470, w_eco150471, w_eco150472, w_eco150473, w_eco150474, w_eco150475, w_eco150476, w_eco150477, w_eco150478, w_eco150479, w_eco150480, w_eco150481, w_eco150482, w_eco150483, w_eco150484, w_eco150485, w_eco150486, w_eco150487, w_eco150488, w_eco150489, w_eco150490, w_eco150491, w_eco150492, w_eco150493, w_eco150494, w_eco150495, w_eco150496, w_eco150497, w_eco150498, w_eco150499, w_eco150500, w_eco150501, w_eco150502, w_eco150503, w_eco150504, w_eco150505, w_eco150506, w_eco150507, w_eco150508, w_eco150509, w_eco150510, w_eco150511, w_eco150512, w_eco150513, w_eco150514, w_eco150515, w_eco150516, w_eco150517, w_eco150518, w_eco150519, w_eco150520, w_eco150521, w_eco150522, w_eco150523, w_eco150524, w_eco150525, w_eco150526, w_eco150527, w_eco150528, w_eco150529, w_eco150530, w_eco150531, w_eco150532, w_eco150533, w_eco150534, w_eco150535, w_eco150536, w_eco150537, w_eco150538, w_eco150539, w_eco150540, w_eco150541, w_eco150542, w_eco150543, w_eco150544, w_eco150545, w_eco150546, w_eco150547, w_eco150548, w_eco150549, w_eco150550, w_eco150551, w_eco150552, w_eco150553, w_eco150554, w_eco150555, w_eco150556, w_eco150557, w_eco150558, w_eco150559, w_eco150560, w_eco150561, w_eco150562, w_eco150563, w_eco150564, w_eco150565, w_eco150566, w_eco150567, w_eco150568, w_eco150569, w_eco150570, w_eco150571, w_eco150572, w_eco150573, w_eco150574, w_eco150575, w_eco150576, w_eco150577, w_eco150578, w_eco150579, w_eco150580, w_eco150581, w_eco150582, w_eco150583, w_eco150584, w_eco150585, w_eco150586, w_eco150587, w_eco150588, w_eco150589, w_eco150590, w_eco150591, w_eco150592, w_eco150593, w_eco150594, w_eco150595, w_eco150596, w_eco150597, w_eco150598, w_eco150599, w_eco150600, w_eco150601, w_eco150602, w_eco150603, w_eco150604, w_eco150605, w_eco150606, w_eco150607, w_eco150608, w_eco150609, w_eco150610, w_eco150611, w_eco150612, w_eco150613, w_eco150614, w_eco150615, w_eco150616, w_eco150617, w_eco150618, w_eco150619, w_eco150620, w_eco150621, w_eco150622, w_eco150623, w_eco150624, w_eco150625, w_eco150626, w_eco150627, w_eco150628, w_eco150629, w_eco150630, w_eco150631, w_eco150632, w_eco150633, w_eco150634, w_eco150635, w_eco150636, w_eco150637, w_eco150638, w_eco150639, w_eco150640, w_eco150641, w_eco150642, w_eco150643, w_eco150644, w_eco150645, w_eco150646, w_eco150647, w_eco150648, w_eco150649, w_eco150650, w_eco150651, w_eco150652, w_eco150653, w_eco150654, w_eco150655, w_eco150656, w_eco150657, w_eco150658, w_eco150659, w_eco150660, w_eco150661, w_eco150662, w_eco150663, w_eco150664, w_eco150665, w_eco150666, w_eco150667, w_eco150668, w_eco150669, w_eco150670, w_eco150671, w_eco150672, w_eco150673, w_eco150674, w_eco150675, w_eco150676, w_eco150677, w_eco150678, w_eco150679, w_eco150680, w_eco150681, w_eco150682, w_eco150683, w_eco150684, w_eco150685, w_eco150686, w_eco150687, w_eco150688, w_eco150689, w_eco150690, w_eco150691, w_eco150692, w_eco150693, w_eco150694, w_eco150695, w_eco150696, w_eco150697, w_eco150698, w_eco150699, w_eco150700, w_eco150701, w_eco150702, w_eco150703, w_eco150704, w_eco150705, w_eco150706, w_eco150707, w_eco150708, w_eco150709, w_eco150710, w_eco150711, w_eco150712, w_eco150713, w_eco150714, w_eco150715, w_eco150716, w_eco150717, w_eco150718, w_eco150719, w_eco150720, w_eco150721, w_eco150722, w_eco150723, w_eco150724, w_eco150725, w_eco150726, w_eco150727, w_eco150728, w_eco150729, w_eco150730, w_eco150731, w_eco150732, w_eco150733, w_eco150734, w_eco150735, w_eco150736, w_eco150737, w_eco150738, w_eco150739, w_eco150740, w_eco150741, w_eco150742, w_eco150743, w_eco150744, w_eco150745, w_eco150746, w_eco150747, w_eco150748, w_eco150749, w_eco150750, w_eco150751, w_eco150752, w_eco150753, w_eco150754, w_eco150755, w_eco150756, w_eco150757, w_eco150758, w_eco150759, w_eco150760, w_eco150761, w_eco150762, w_eco150763, w_eco150764, w_eco150765, w_eco150766, w_eco150767, w_eco150768, w_eco150769, w_eco150770, w_eco150771, w_eco150772, w_eco150773, w_eco150774, w_eco150775, w_eco150776, w_eco150777, w_eco150778, w_eco150779, w_eco150780, w_eco150781, w_eco150782, w_eco150783, w_eco150784, w_eco150785, w_eco150786, w_eco150787, w_eco150788, w_eco150789, w_eco150790, w_eco150791, w_eco150792, w_eco150793, w_eco150794, w_eco150795, w_eco150796, w_eco150797, w_eco150798, w_eco150799, w_eco150800, w_eco150801, w_eco150802, w_eco150803, w_eco150804, w_eco150805, w_eco150806, w_eco150807, w_eco150808, w_eco150809, w_eco150810, w_eco150811, w_eco150812, w_eco150813, w_eco150814, w_eco150815, w_eco150816, w_eco150817, w_eco150818, w_eco150819, w_eco150820, w_eco150821, w_eco150822, w_eco150823, w_eco150824, w_eco150825, w_eco150826, w_eco150827, w_eco150828, w_eco150829, w_eco150830, w_eco150831, w_eco150832, w_eco150833, w_eco150834, w_eco150835, w_eco150836, w_eco150837, w_eco150838, w_eco150839, w_eco150840, w_eco150841, w_eco150842, w_eco150843, w_eco150844, w_eco150845, w_eco150846, w_eco150847, w_eco150848, w_eco150849, w_eco150850, w_eco150851, w_eco150852, w_eco150853, w_eco150854, w_eco150855, w_eco150856, w_eco150857, w_eco150858, w_eco150859, w_eco150860, w_eco150861, w_eco150862, w_eco150863, w_eco150864, w_eco150865, w_eco150866, w_eco150867, w_eco150868, w_eco150869, w_eco150870, w_eco150871, w_eco150872, w_eco150873, w_eco150874, w_eco150875, w_eco150876, w_eco150877, w_eco150878, w_eco150879, w_eco150880, w_eco150881, w_eco150882, w_eco150883, w_eco150884, w_eco150885, w_eco150886, w_eco150887, w_eco150888, w_eco150889, w_eco150890, w_eco150891, w_eco150892, w_eco150893, w_eco150894, w_eco150895, w_eco150896, w_eco150897, w_eco150898, w_eco150899, w_eco150900, w_eco150901, w_eco150902, w_eco150903, w_eco150904, w_eco150905, w_eco150906, w_eco150907, w_eco150908, w_eco150909, w_eco150910, w_eco150911, w_eco150912, w_eco150913, w_eco150914, w_eco150915, w_eco150916, w_eco150917, w_eco150918, w_eco150919, w_eco150920, w_eco150921, w_eco150922, w_eco150923, w_eco150924, w_eco150925, w_eco150926, w_eco150927, w_eco150928, w_eco150929, w_eco150930, w_eco150931, w_eco150932, w_eco150933, w_eco150934, w_eco150935, w_eco150936, w_eco150937, w_eco150938, w_eco150939, w_eco150940, w_eco150941, w_eco150942, w_eco150943, w_eco150944, w_eco150945, w_eco150946, w_eco150947, w_eco150948, w_eco150949, w_eco150950, w_eco150951, w_eco150952, w_eco150953, w_eco150954, w_eco150955, w_eco150956, w_eco150957, w_eco150958, w_eco150959, w_eco150960, w_eco150961, w_eco150962, w_eco150963, w_eco150964, w_eco150965, w_eco150966, w_eco150967, w_eco150968, w_eco150969, w_eco150970, w_eco150971, w_eco150972, w_eco150973, w_eco150974, w_eco150975, w_eco150976, w_eco150977, w_eco150978, w_eco150979, w_eco150980, w_eco150981, w_eco150982, w_eco150983, w_eco150984, w_eco150985, w_eco150986, w_eco150987, w_eco150988, w_eco150989, w_eco150990, w_eco150991, w_eco150992, w_eco150993, w_eco150994, w_eco150995, w_eco150996, w_eco150997, w_eco150998, w_eco150999, w_eco151000, w_eco151001, w_eco151002, w_eco151003, w_eco151004, w_eco151005, w_eco151006, w_eco151007, w_eco151008, w_eco151009, w_eco151010, w_eco151011, w_eco151012, w_eco151013, w_eco151014, w_eco151015, w_eco151016, w_eco151017, w_eco151018, w_eco151019, w_eco151020, w_eco151021, w_eco151022, w_eco151023, w_eco151024, w_eco151025, w_eco151026, w_eco151027, w_eco151028, w_eco151029, w_eco151030, w_eco151031, w_eco151032, w_eco151033, w_eco151034, w_eco151035, w_eco151036, w_eco151037, w_eco151038, w_eco151039, w_eco151040, w_eco151041, w_eco151042, w_eco151043, w_eco151044, w_eco151045, w_eco151046, w_eco151047, w_eco151048, w_eco151049, w_eco151050, w_eco151051, w_eco151052, w_eco151053, w_eco151054, w_eco151055, w_eco151056, w_eco151057, w_eco151058, w_eco151059, w_eco151060, w_eco151061, w_eco151062, w_eco151063, w_eco151064, w_eco151065, w_eco151066, w_eco151067, w_eco151068, w_eco151069, w_eco151070, w_eco151071, w_eco151072, w_eco151073, w_eco151074, w_eco151075, w_eco151076, w_eco151077, w_eco151078, w_eco151079, w_eco151080, w_eco151081, w_eco151082, w_eco151083, w_eco151084, w_eco151085, w_eco151086, w_eco151087, w_eco151088, w_eco151089, w_eco151090, w_eco151091, w_eco151092, w_eco151093, w_eco151094, w_eco151095, w_eco151096, w_eco151097, w_eco151098, w_eco151099, w_eco151100, w_eco151101, w_eco151102, w_eco151103, w_eco151104, w_eco151105, w_eco151106, w_eco151107, w_eco151108, w_eco151109, w_eco151110, w_eco151111, w_eco151112, w_eco151113, w_eco151114, w_eco151115, w_eco151116, w_eco151117, w_eco151118, w_eco151119, w_eco151120, w_eco151121, w_eco151122, w_eco151123, w_eco151124, w_eco151125, w_eco151126, w_eco151127, w_eco151128, w_eco151129, w_eco151130, w_eco151131, w_eco151132, w_eco151133, w_eco151134, w_eco151135, w_eco151136, w_eco151137, w_eco151138, w_eco151139, w_eco151140, w_eco151141, w_eco151142, w_eco151143, w_eco151144, w_eco151145, w_eco151146, w_eco151147, w_eco151148, w_eco151149, w_eco151150, w_eco151151, w_eco151152, w_eco151153, w_eco151154, w_eco151155, w_eco151156, w_eco151157, w_eco151158, w_eco151159, w_eco151160, w_eco151161, w_eco151162, w_eco151163, w_eco151164, w_eco151165, w_eco151166, w_eco151167, w_eco151168, w_eco151169, w_eco151170, w_eco151171, w_eco151172, w_eco151173, w_eco151174, w_eco151175, w_eco151176, w_eco151177, w_eco151178, w_eco151179, w_eco151180, w_eco151181, w_eco151182, w_eco151183, w_eco151184, w_eco151185, w_eco151186, w_eco151187, w_eco151188, w_eco151189, w_eco151190, w_eco151191, w_eco151192, w_eco151193, w_eco151194, w_eco151195, w_eco151196, w_eco151197, w_eco151198, w_eco151199, w_eco151200, w_eco151201, w_eco151202, w_eco151203, w_eco151204, w_eco151205, w_eco151206, w_eco151207, w_eco151208, w_eco151209, w_eco151210, w_eco151211, w_eco151212, w_eco151213, w_eco151214, w_eco151215, w_eco151216, w_eco151217, w_eco151218, w_eco151219, w_eco151220, w_eco151221, w_eco151222, w_eco151223, w_eco151224, w_eco151225, w_eco151226, w_eco151227, w_eco151228, w_eco151229, w_eco151230, w_eco151231, w_eco151232, w_eco151233, w_eco151234, w_eco151235, w_eco151236, w_eco151237, w_eco151238, w_eco151239, w_eco151240, w_eco151241, w_eco151242, w_eco151243, w_eco151244, w_eco151245, w_eco151246, w_eco151247, w_eco151248, w_eco151249, w_eco151250, w_eco151251, w_eco151252, w_eco151253, w_eco151254, w_eco151255, w_eco151256, w_eco151257, w_eco151258, w_eco151259, w_eco151260, w_eco151261, w_eco151262, w_eco151263, w_eco151264, w_eco151265, w_eco151266, w_eco151267, w_eco151268, w_eco151269, w_eco151270, w_eco151271, w_eco151272, w_eco151273, w_eco151274, w_eco151275, w_eco151276, w_eco151277, w_eco151278, w_eco151279, w_eco151280, w_eco151281, w_eco151282, w_eco151283, w_eco151284, w_eco151285, w_eco151286, w_eco151287, w_eco151288, w_eco151289, w_eco151290, w_eco151291, w_eco151292, w_eco151293, w_eco151294, w_eco151295, w_eco151296, w_eco151297, w_eco151298, w_eco151299, w_eco151300, w_eco151301, w_eco151302, w_eco151303, w_eco151304, w_eco151305, w_eco151306, w_eco151307, w_eco151308, w_eco151309, w_eco151310, w_eco151311, w_eco151312, w_eco151313, w_eco151314, w_eco151315, w_eco151316, w_eco151317, w_eco151318, w_eco151319, w_eco151320, w_eco151321, w_eco151322, w_eco151323, w_eco151324, w_eco151325, w_eco151326, w_eco151327, w_eco151328, w_eco151329, w_eco151330, w_eco151331, w_eco151332, w_eco151333, w_eco151334, w_eco151335, w_eco151336, w_eco151337, w_eco151338, w_eco151339, w_eco151340, w_eco151341, w_eco151342, w_eco151343, w_eco151344, w_eco151345, w_eco151346, w_eco151347, w_eco151348, w_eco151349, w_eco151350, w_eco151351, w_eco151352, w_eco151353, w_eco151354, w_eco151355, w_eco151356, w_eco151357, w_eco151358, w_eco151359, w_eco151360, w_eco151361, w_eco151362, w_eco151363, w_eco151364, w_eco151365, w_eco151366, w_eco151367, w_eco151368, w_eco151369, w_eco151370, w_eco151371, w_eco151372, w_eco151373, w_eco151374, w_eco151375, w_eco151376, w_eco151377, w_eco151378, w_eco151379, w_eco151380, w_eco151381, w_eco151382, w_eco151383, w_eco151384, w_eco151385, w_eco151386, w_eco151387, w_eco151388, w_eco151389, w_eco151390, w_eco151391, w_eco151392, w_eco151393, w_eco151394, w_eco151395, w_eco151396, w_eco151397, w_eco151398, w_eco151399, w_eco151400, w_eco151401, w_eco151402, w_eco151403, w_eco151404, w_eco151405, w_eco151406, w_eco151407, w_eco151408, w_eco151409, w_eco151410, w_eco151411, w_eco151412, w_eco151413, w_eco151414, w_eco151415, w_eco151416, w_eco151417, w_eco151418, w_eco151419, w_eco151420, w_eco151421, w_eco151422, w_eco151423, w_eco151424, w_eco151425, w_eco151426, w_eco151427, w_eco151428, w_eco151429, w_eco151430, w_eco151431, w_eco151432, w_eco151433, w_eco151434, w_eco151435, w_eco151436, w_eco151437, w_eco151438, w_eco151439, w_eco151440, w_eco151441, w_eco151442, w_eco151443, w_eco151444, w_eco151445, w_eco151446, w_eco151447, w_eco151448, w_eco151449, w_eco151450, w_eco151451, w_eco151452, w_eco151453, w_eco151454, w_eco151455, w_eco151456, w_eco151457, w_eco151458, w_eco151459, w_eco151460, w_eco151461, w_eco151462, w_eco151463, w_eco151464, w_eco151465, w_eco151466, w_eco151467, w_eco151468, w_eco151469, w_eco151470, w_eco151471, w_eco151472, w_eco151473, w_eco151474, w_eco151475, w_eco151476, w_eco151477, w_eco151478, w_eco151479, w_eco151480, w_eco151481, w_eco151482, w_eco151483, w_eco151484, w_eco151485, w_eco151486, w_eco151487, w_eco151488, w_eco151489, w_eco151490, w_eco151491, w_eco151492, w_eco151493, w_eco151494, w_eco151495, w_eco151496, w_eco151497, w_eco151498, w_eco151499, w_eco151500, w_eco151501, w_eco151502, w_eco151503, w_eco151504, w_eco151505, w_eco151506, w_eco151507, w_eco151508, w_eco151509, w_eco151510, w_eco151511, w_eco151512, w_eco151513, w_eco151514, w_eco151515, w_eco151516, w_eco151517, w_eco151518, w_eco151519, w_eco151520, w_eco151521, w_eco151522, w_eco151523, w_eco151524, w_eco151525, w_eco151526, w_eco151527, w_eco151528, w_eco151529, w_eco151530, w_eco151531, w_eco151532, w_eco151533, w_eco151534, w_eco151535, w_eco151536, w_eco151537, w_eco151538, w_eco151539, w_eco151540, w_eco151541, w_eco151542, w_eco151543, w_eco151544, w_eco151545, w_eco151546, w_eco151547, w_eco151548, w_eco151549, w_eco151550, w_eco151551, w_eco151552, w_eco151553, w_eco151554, w_eco151555, w_eco151556, w_eco151557, w_eco151558, w_eco151559, w_eco151560, w_eco151561, w_eco151562, w_eco151563, w_eco151564, w_eco151565, w_eco151566, w_eco151567, w_eco151568, w_eco151569, w_eco151570, w_eco151571, w_eco151572, w_eco151573, w_eco151574, w_eco151575, w_eco151576, w_eco151577, w_eco151578, w_eco151579, w_eco151580, w_eco151581, w_eco151582, w_eco151583, w_eco151584, w_eco151585, w_eco151586, w_eco151587, w_eco151588, w_eco151589, w_eco151590, w_eco151591, w_eco151592, w_eco151593, w_eco151594, w_eco151595, w_eco151596, w_eco151597, w_eco151598, w_eco151599, w_eco151600, w_eco151601, w_eco151602, w_eco151603, w_eco151604, w_eco151605, w_eco151606, w_eco151607, w_eco151608, w_eco151609, w_eco151610, w_eco151611, w_eco151612, w_eco151613, w_eco151614, w_eco151615, w_eco151616, w_eco151617, w_eco151618, w_eco151619, w_eco151620, w_eco151621, w_eco151622, w_eco151623, w_eco151624, w_eco151625, w_eco151626, w_eco151627, w_eco151628, w_eco151629, w_eco151630, w_eco151631, w_eco151632, w_eco151633, w_eco151634, w_eco151635, w_eco151636, w_eco151637, w_eco151638, w_eco151639, w_eco151640, w_eco151641, w_eco151642, w_eco151643, w_eco151644, w_eco151645, w_eco151646, w_eco151647, w_eco151648, w_eco151649, w_eco151650, w_eco151651, w_eco151652, w_eco151653, w_eco151654, w_eco151655, w_eco151656, w_eco151657, w_eco151658, w_eco151659, w_eco151660, w_eco151661, w_eco151662, w_eco151663, w_eco151664, w_eco151665, w_eco151666, w_eco151667, w_eco151668, w_eco151669, w_eco151670, w_eco151671, w_eco151672, w_eco151673, w_eco151674, w_eco151675, w_eco151676, w_eco151677, w_eco151678, w_eco151679, w_eco151680, w_eco151681, w_eco151682, w_eco151683, w_eco151684, w_eco151685, w_eco151686, w_eco151687, w_eco151688, w_eco151689, w_eco151690, w_eco151691, w_eco151692, w_eco151693, w_eco151694, w_eco151695, w_eco151696, w_eco151697, w_eco151698, w_eco151699, w_eco151700, w_eco151701, w_eco151702, w_eco151703, w_eco151704, w_eco151705, w_eco151706, w_eco151707, w_eco151708, w_eco151709, w_eco151710, w_eco151711, w_eco151712, w_eco151713, w_eco151714, w_eco151715, w_eco151716, w_eco151717, w_eco151718, w_eco151719, w_eco151720, w_eco151721, w_eco151722, w_eco151723, w_eco151724, w_eco151725, w_eco151726, w_eco151727, w_eco151728, w_eco151729, w_eco151730, w_eco151731, w_eco151732, w_eco151733, w_eco151734, w_eco151735, w_eco151736, w_eco151737, w_eco151738, w_eco151739, w_eco151740, w_eco151741, w_eco151742, w_eco151743, w_eco151744, w_eco151745, w_eco151746, w_eco151747, w_eco151748, w_eco151749, w_eco151750, w_eco151751, w_eco151752, w_eco151753, w_eco151754, w_eco151755, w_eco151756, w_eco151757, w_eco151758, w_eco151759, w_eco151760, w_eco151761, w_eco151762, w_eco151763, w_eco151764, w_eco151765, w_eco151766, w_eco151767, w_eco151768, w_eco151769, w_eco151770, w_eco151771, w_eco151772, w_eco151773, w_eco151774, w_eco151775, w_eco151776, w_eco151777, w_eco151778, w_eco151779, w_eco151780, w_eco151781, w_eco151782, w_eco151783, w_eco151784, w_eco151785, w_eco151786, w_eco151787, w_eco151788, w_eco151789, w_eco151790, w_eco151791, w_eco151792, w_eco151793, w_eco151794, w_eco151795, w_eco151796, w_eco151797, w_eco151798, w_eco151799, w_eco151800, w_eco151801, w_eco151802, w_eco151803, w_eco151804, w_eco151805, w_eco151806, w_eco151807, w_eco151808, w_eco151809, w_eco151810, w_eco151811, w_eco151812, w_eco151813, w_eco151814, w_eco151815, w_eco151816, w_eco151817, w_eco151818, w_eco151819, w_eco151820, w_eco151821, w_eco151822, w_eco151823, w_eco151824, w_eco151825, w_eco151826, w_eco151827, w_eco151828, w_eco151829, w_eco151830, w_eco151831, w_eco151832, w_eco151833, w_eco151834, w_eco151835, w_eco151836, w_eco151837, w_eco151838, w_eco151839, w_eco151840, w_eco151841, w_eco151842, w_eco151843, w_eco151844, w_eco151845, w_eco151846, w_eco151847, w_eco151848, w_eco151849, w_eco151850, w_eco151851, w_eco151852, w_eco151853, w_eco151854, w_eco151855, w_eco151856, w_eco151857, w_eco151858, w_eco151859, w_eco151860, w_eco151861, w_eco151862, w_eco151863, w_eco151864, w_eco151865, w_eco151866, w_eco151867, w_eco151868, w_eco151869, w_eco151870, w_eco151871, w_eco151872, w_eco151873, w_eco151874, w_eco151875, w_eco151876, w_eco151877, w_eco151878, w_eco151879, w_eco151880, w_eco151881, w_eco151882, w_eco151883, w_eco151884, w_eco151885, w_eco151886, w_eco151887, w_eco151888, w_eco151889, w_eco151890, w_eco151891, w_eco151892, w_eco151893, w_eco151894, w_eco151895, w_eco151896, w_eco151897, w_eco151898, w_eco151899, w_eco151900, w_eco151901, w_eco151902, w_eco151903, w_eco151904, w_eco151905, w_eco151906, w_eco151907, w_eco151908, w_eco151909, w_eco151910, w_eco151911, w_eco151912, w_eco151913, w_eco151914, w_eco151915, w_eco151916, w_eco151917, w_eco151918, w_eco151919, w_eco151920, w_eco151921, w_eco151922, w_eco151923, w_eco151924, w_eco151925, w_eco151926, w_eco151927, w_eco151928, w_eco151929, w_eco151930, w_eco151931, w_eco151932, w_eco151933, w_eco151934, w_eco151935, w_eco151936, w_eco151937, w_eco151938, w_eco151939, w_eco151940, w_eco151941, w_eco151942, w_eco151943, w_eco151944, w_eco151945, w_eco151946, w_eco151947, w_eco151948, w_eco151949, w_eco151950, w_eco151951, w_eco151952, w_eco151953, w_eco151954, w_eco151955, w_eco151956, w_eco151957, w_eco151958, w_eco151959, w_eco151960, w_eco151961, w_eco151962, w_eco151963, w_eco151964, w_eco151965, w_eco151966, w_eco151967, w_eco151968, w_eco151969, w_eco151970, w_eco151971, w_eco151972, w_eco151973, w_eco151974, w_eco151975, w_eco151976, w_eco151977, w_eco151978, w_eco151979, w_eco151980, w_eco151981, w_eco151982, w_eco151983, w_eco151984, w_eco151985, w_eco151986, w_eco151987, w_eco151988, w_eco151989, w_eco151990, w_eco151991, w_eco151992, w_eco151993, w_eco151994, w_eco151995, w_eco151996, w_eco151997, w_eco151998, w_eco151999, w_eco152000, w_eco152001, w_eco152002, w_eco152003, w_eco152004, w_eco152005, w_eco152006, w_eco152007, w_eco152008, w_eco152009, w_eco152010, w_eco152011, w_eco152012, w_eco152013, w_eco152014, w_eco152015, w_eco152016, w_eco152017, w_eco152018, w_eco152019, w_eco152020, w_eco152021, w_eco152022, w_eco152023, w_eco152024, w_eco152025, w_eco152026, w_eco152027, w_eco152028, w_eco152029, w_eco152030, w_eco152031, w_eco152032, w_eco152033, w_eco152034, w_eco152035, w_eco152036, w_eco152037, w_eco152038, w_eco152039, w_eco152040, w_eco152041, w_eco152042, w_eco152043, w_eco152044, w_eco152045, w_eco152046, w_eco152047, w_eco152048, w_eco152049, w_eco152050, w_eco152051, w_eco152052, w_eco152053, w_eco152054, w_eco152055, w_eco152056, w_eco152057, w_eco152058, w_eco152059, w_eco152060, w_eco152061, w_eco152062, w_eco152063, w_eco152064, w_eco152065, w_eco152066, w_eco152067, w_eco152068, w_eco152069, w_eco152070, w_eco152071, w_eco152072, w_eco152073, w_eco152074, w_eco152075, w_eco152076, w_eco152077, w_eco152078, w_eco152079, w_eco152080, w_eco152081, w_eco152082, w_eco152083, w_eco152084, w_eco152085, w_eco152086, w_eco152087, w_eco152088, w_eco152089, w_eco152090, w_eco152091, w_eco152092, w_eco152093, w_eco152094, w_eco152095, w_eco152096, w_eco152097, w_eco152098, w_eco152099, w_eco152100, w_eco152101, w_eco152102, w_eco152103, w_eco152104, w_eco152105, w_eco152106, w_eco152107, w_eco152108, w_eco152109, w_eco152110, w_eco152111, w_eco152112, w_eco152113, w_eco152114, w_eco152115, w_eco152116, w_eco152117, w_eco152118, w_eco152119, w_eco152120, w_eco152121, w_eco152122, w_eco152123, w_eco152124, w_eco152125, w_eco152126, w_eco152127, w_eco152128, w_eco152129, w_eco152130, w_eco152131, w_eco152132, w_eco152133, w_eco152134, w_eco152135, w_eco152136, w_eco152137, w_eco152138, w_eco152139, w_eco152140, w_eco152141, w_eco152142, w_eco152143, w_eco152144, w_eco152145, w_eco152146, w_eco152147, w_eco152148, w_eco152149, w_eco152150, w_eco152151, w_eco152152, w_eco152153, w_eco152154, w_eco152155, w_eco152156, w_eco152157, w_eco152158, w_eco152159, w_eco152160, w_eco152161, w_eco152162, w_eco152163, w_eco152164, w_eco152165, w_eco152166, w_eco152167, w_eco152168, w_eco152169, w_eco152170, w_eco152171, w_eco152172, w_eco152173, w_eco152174, w_eco152175, w_eco152176, w_eco152177, w_eco152178, w_eco152179, w_eco152180, w_eco152181, w_eco152182, w_eco152183, w_eco152184, w_eco152185, w_eco152186, w_eco152187, w_eco152188, w_eco152189, w_eco152190, w_eco152191, w_eco152192, w_eco152193, w_eco152194, w_eco152195, w_eco152196, w_eco152197, w_eco152198, w_eco152199, w_eco152200, w_eco152201, w_eco152202, w_eco152203, w_eco152204, w_eco152205, w_eco152206, w_eco152207, w_eco152208, w_eco152209, w_eco152210, w_eco152211, w_eco152212, w_eco152213, w_eco152214, w_eco152215, w_eco152216, w_eco152217, w_eco152218, w_eco152219, w_eco152220, w_eco152221, w_eco152222, w_eco152223, w_eco152224, w_eco152225, w_eco152226, w_eco152227, w_eco152228, w_eco152229, w_eco152230, w_eco152231, w_eco152232, w_eco152233, w_eco152234, w_eco152235, w_eco152236, w_eco152237, w_eco152238, w_eco152239, w_eco152240, w_eco152241, w_eco152242, w_eco152243, w_eco152244, w_eco152245, w_eco152246, w_eco152247, w_eco152248, w_eco152249, w_eco152250, w_eco152251, w_eco152252, w_eco152253, w_eco152254, w_eco152255, w_eco152256, w_eco152257, w_eco152258, w_eco152259, w_eco152260, w_eco152261, w_eco152262, w_eco152263, w_eco152264, w_eco152265, w_eco152266, w_eco152267, w_eco152268, w_eco152269, w_eco152270, w_eco152271, w_eco152272, w_eco152273, w_eco152274, w_eco152275, w_eco152276, w_eco152277, w_eco152278, w_eco152279, w_eco152280, w_eco152281, w_eco152282, w_eco152283, w_eco152284, w_eco152285, w_eco152286, w_eco152287, w_eco152288, w_eco152289, w_eco152290, w_eco152291, w_eco152292, w_eco152293, w_eco152294, w_eco152295, w_eco152296, w_eco152297, w_eco152298, w_eco152299, w_eco152300, w_eco152301, w_eco152302, w_eco152303, w_eco152304, w_eco152305, w_eco152306, w_eco152307, w_eco152308, w_eco152309, w_eco152310, w_eco152311, w_eco152312, w_eco152313, w_eco152314, w_eco152315, w_eco152316, w_eco152317, w_eco152318, w_eco152319, w_eco152320, w_eco152321, w_eco152322, w_eco152323, w_eco152324, w_eco152325, w_eco152326, w_eco152327, w_eco152328, w_eco152329, w_eco152330, w_eco152331, w_eco152332, w_eco152333, w_eco152334, w_eco152335, w_eco152336, w_eco152337, w_eco152338, w_eco152339, w_eco152340, w_eco152341, w_eco152342, w_eco152343, w_eco152344, w_eco152345, w_eco152346, w_eco152347, w_eco152348, w_eco152349, w_eco152350, w_eco152351, w_eco152352, w_eco152353, w_eco152354, w_eco152355, w_eco152356, w_eco152357, w_eco152358, w_eco152359, w_eco152360, w_eco152361, w_eco152362, w_eco152363, w_eco152364, w_eco152365, w_eco152366, w_eco152367, w_eco152368, w_eco152369, w_eco152370, w_eco152371, w_eco152372, w_eco152373, w_eco152374, w_eco152375, w_eco152376, w_eco152377, w_eco152378, w_eco152379, w_eco152380, w_eco152381, w_eco152382, w_eco152383, w_eco152384, w_eco152385, w_eco152386, w_eco152387, w_eco152388, w_eco152389, w_eco152390, w_eco152391, w_eco152392, w_eco152393, w_eco152394, w_eco152395, w_eco152396, w_eco152397, w_eco152398, w_eco152399, w_eco152400, w_eco152401, w_eco152402, w_eco152403, w_eco152404, w_eco152405, w_eco152406, w_eco152407, w_eco152408, w_eco152409, w_eco152410, w_eco152411, w_eco152412, w_eco152413, w_eco152414, w_eco152415, w_eco152416, w_eco152417, w_eco152418, w_eco152419, w_eco152420, w_eco152421, w_eco152422, w_eco152423, w_eco152424, w_eco152425, w_eco152426, w_eco152427, w_eco152428, w_eco152429, w_eco152430, w_eco152431, w_eco152432, w_eco152433, w_eco152434, w_eco152435, w_eco152436, w_eco152437, w_eco152438, w_eco152439, w_eco152440, w_eco152441, w_eco152442, w_eco152443, w_eco152444, w_eco152445, w_eco152446, w_eco152447, w_eco152448, w_eco152449, w_eco152450, w_eco152451, w_eco152452, w_eco152453, w_eco152454, w_eco152455, w_eco152456, w_eco152457, w_eco152458, w_eco152459, w_eco152460, w_eco152461, w_eco152462, w_eco152463, w_eco152464, w_eco152465, w_eco152466, w_eco152467, w_eco152468, w_eco152469, w_eco152470, w_eco152471, w_eco152472, w_eco152473, w_eco152474, w_eco152475, w_eco152476, w_eco152477, w_eco152478, w_eco152479, w_eco152480, w_eco152481, w_eco152482, w_eco152483, w_eco152484, w_eco152485, w_eco152486, w_eco152487, w_eco152488, w_eco152489, w_eco152490, w_eco152491, w_eco152492, w_eco152493, w_eco152494, w_eco152495, w_eco152496, w_eco152497, w_eco152498, w_eco152499, w_eco152500, w_eco152501, w_eco152502, w_eco152503, w_eco152504, w_eco152505, w_eco152506, w_eco152507, w_eco152508, w_eco152509, w_eco152510, w_eco152511, w_eco152512, w_eco152513, w_eco152514, w_eco152515, w_eco152516, w_eco152517, w_eco152518, w_eco152519, w_eco152520, w_eco152521, w_eco152522, w_eco152523, w_eco152524, w_eco152525, w_eco152526, w_eco152527, w_eco152528, w_eco152529, w_eco152530, w_eco152531, w_eco152532, w_eco152533, w_eco152534, w_eco152535, w_eco152536, w_eco152537, w_eco152538, w_eco152539, w_eco152540, w_eco152541, w_eco152542, w_eco152543, w_eco152544, w_eco152545, w_eco152546, w_eco152547, w_eco152548, w_eco152549, w_eco152550, w_eco152551, w_eco152552, w_eco152553, w_eco152554, w_eco152555, w_eco152556, w_eco152557, w_eco152558, w_eco152559, w_eco152560, w_eco152561, w_eco152562, w_eco152563, w_eco152564, w_eco152565, w_eco152566, w_eco152567, w_eco152568, w_eco152569, w_eco152570, w_eco152571, w_eco152572, w_eco152573, w_eco152574, w_eco152575, w_eco152576, w_eco152577, w_eco152578, w_eco152579, w_eco152580, w_eco152581, w_eco152582, w_eco152583, w_eco152584, w_eco152585, w_eco152586, w_eco152587, w_eco152588, w_eco152589, w_eco152590, w_eco152591, w_eco152592, w_eco152593, w_eco152594, w_eco152595, w_eco152596, w_eco152597, w_eco152598, w_eco152599, w_eco152600, w_eco152601, w_eco152602, w_eco152603, w_eco152604, w_eco152605, w_eco152606, w_eco152607, w_eco152608, w_eco152609, w_eco152610, w_eco152611, w_eco152612, w_eco152613, w_eco152614, w_eco152615, w_eco152616, w_eco152617, w_eco152618, w_eco152619, w_eco152620, w_eco152621, w_eco152622, w_eco152623, w_eco152624, w_eco152625, w_eco152626, w_eco152627, w_eco152628, w_eco152629, w_eco152630, w_eco152631, w_eco152632, w_eco152633, w_eco152634, w_eco152635, w_eco152636, w_eco152637, w_eco152638, w_eco152639, w_eco152640, w_eco152641, w_eco152642, w_eco152643, w_eco152644, w_eco152645, w_eco152646, w_eco152647, w_eco152648, w_eco152649, w_eco152650, w_eco152651, w_eco152652, w_eco152653, w_eco152654, w_eco152655, w_eco152656, w_eco152657, w_eco152658, w_eco152659, w_eco152660, w_eco152661, w_eco152662, w_eco152663, w_eco152664, w_eco152665, w_eco152666, w_eco152667, w_eco152668, w_eco152669, w_eco152670, w_eco152671, w_eco152672, w_eco152673, w_eco152674, w_eco152675, w_eco152676, w_eco152677, w_eco152678, w_eco152679, w_eco152680, w_eco152681, w_eco152682, w_eco152683, w_eco152684, w_eco152685, w_eco152686, w_eco152687, w_eco152688, w_eco152689, w_eco152690, w_eco152691, w_eco152692, w_eco152693, w_eco152694, w_eco152695, w_eco152696, w_eco152697, w_eco152698, w_eco152699, w_eco152700, w_eco152701, w_eco152702, w_eco152703, w_eco152704, w_eco152705, w_eco152706, w_eco152707, w_eco152708, w_eco152709, w_eco152710, w_eco152711, w_eco152712, w_eco152713, w_eco152714, w_eco152715, w_eco152716, w_eco152717, w_eco152718, w_eco152719, w_eco152720, w_eco152721, w_eco152722, w_eco152723, w_eco152724, w_eco152725, w_eco152726, w_eco152727, w_eco152728, w_eco152729, w_eco152730, w_eco152731, w_eco152732, w_eco152733, w_eco152734, w_eco152735, w_eco152736, w_eco152737, w_eco152738, w_eco152739, w_eco152740, w_eco152741, w_eco152742, w_eco152743, w_eco152744, w_eco152745, w_eco152746, w_eco152747, w_eco152748, w_eco152749, w_eco152750, w_eco152751, w_eco152752, w_eco152753, w_eco152754, w_eco152755, w_eco152756, w_eco152757, w_eco152758, w_eco152759, w_eco152760, w_eco152761, w_eco152762, w_eco152763, w_eco152764, w_eco152765, w_eco152766, w_eco152767, w_eco152768, w_eco152769, w_eco152770, w_eco152771, w_eco152772, w_eco152773, w_eco152774, w_eco152775, w_eco152776, w_eco152777, w_eco152778, w_eco152779, w_eco152780, w_eco152781, w_eco152782, w_eco152783, w_eco152784, w_eco152785, w_eco152786, w_eco152787, w_eco152788, w_eco152789, w_eco152790, w_eco152791, w_eco152792, w_eco152793, w_eco152794, w_eco152795, w_eco152796, w_eco152797, w_eco152798, w_eco152799, w_eco152800, w_eco152801, w_eco152802, w_eco152803, w_eco152804, w_eco152805, w_eco152806, w_eco152807, w_eco152808, w_eco152809, w_eco152810, w_eco152811, w_eco152812, w_eco152813, w_eco152814, w_eco152815, w_eco152816, w_eco152817, w_eco152818, w_eco152819, w_eco152820, w_eco152821, w_eco152822, w_eco152823, w_eco152824, w_eco152825, w_eco152826, w_eco152827, w_eco152828, w_eco152829, w_eco152830, w_eco152831, w_eco152832, w_eco152833, w_eco152834, w_eco152835, w_eco152836, w_eco152837, w_eco152838, w_eco152839, w_eco152840, w_eco152841, w_eco152842, w_eco152843, w_eco152844, w_eco152845, w_eco152846, w_eco152847, w_eco152848, w_eco152849, w_eco152850, w_eco152851, w_eco152852, w_eco152853, w_eco152854, w_eco152855, w_eco152856, w_eco152857, w_eco152858, w_eco152859, w_eco152860, w_eco152861, w_eco152862, w_eco152863, w_eco152864, w_eco152865, w_eco152866, w_eco152867, w_eco152868, w_eco152869, w_eco152870, w_eco152871, w_eco152872, w_eco152873, w_eco152874, w_eco152875, w_eco152876, w_eco152877, w_eco152878, w_eco152879, w_eco152880, w_eco152881, w_eco152882, w_eco152883, w_eco152884, w_eco152885, w_eco152886, w_eco152887, w_eco152888, w_eco152889, w_eco152890, w_eco152891, w_eco152892, w_eco152893, w_eco152894, w_eco152895, w_eco152896, w_eco152897, w_eco152898, w_eco152899, w_eco152900, w_eco152901, w_eco152902, w_eco152903, w_eco152904, w_eco152905, w_eco152906, w_eco152907, w_eco152908, w_eco152909, w_eco152910, w_eco152911, w_eco152912, w_eco152913, w_eco152914, w_eco152915, w_eco152916, w_eco152917, w_eco152918, w_eco152919, w_eco152920, w_eco152921, w_eco152922, w_eco152923, w_eco152924, w_eco152925, w_eco152926, w_eco152927, w_eco152928, w_eco152929, w_eco152930, w_eco152931, w_eco152932, w_eco152933, w_eco152934, w_eco152935, w_eco152936, w_eco152937, w_eco152938, w_eco152939, w_eco152940, w_eco152941, w_eco152942, w_eco152943, w_eco152944, w_eco152945, w_eco152946, w_eco152947, w_eco152948, w_eco152949, w_eco152950, w_eco152951, w_eco152952, w_eco152953, w_eco152954, w_eco152955, w_eco152956, w_eco152957, w_eco152958, w_eco152959, w_eco152960, w_eco152961, w_eco152962, w_eco152963, w_eco152964, w_eco152965, w_eco152966, w_eco152967, w_eco152968, w_eco152969, w_eco152970, w_eco152971, w_eco152972, w_eco152973, w_eco152974, w_eco152975, w_eco152976, w_eco152977, w_eco152978, w_eco152979, w_eco152980, w_eco152981, w_eco152982, w_eco152983, w_eco152984, w_eco152985, w_eco152986, w_eco152987, w_eco152988, w_eco152989, w_eco152990, w_eco152991, w_eco152992, w_eco152993, w_eco152994, w_eco152995, w_eco152996, w_eco152997, w_eco152998, w_eco152999, w_eco153000, w_eco153001, w_eco153002, w_eco153003, w_eco153004, w_eco153005, w_eco153006, w_eco153007, w_eco153008, w_eco153009, w_eco153010, w_eco153011, w_eco153012, w_eco153013, w_eco153014, w_eco153015, w_eco153016, w_eco153017, w_eco153018, w_eco153019, w_eco153020, w_eco153021, w_eco153022, w_eco153023, w_eco153024, w_eco153025, w_eco153026, w_eco153027, w_eco153028, w_eco153029, w_eco153030, w_eco153031, w_eco153032, w_eco153033, w_eco153034, w_eco153035, w_eco153036, w_eco153037, w_eco153038, w_eco153039, w_eco153040, w_eco153041, w_eco153042, w_eco153043, w_eco153044, w_eco153045, w_eco153046, w_eco153047, w_eco153048, w_eco153049, w_eco153050, w_eco153051, w_eco153052, w_eco153053, w_eco153054, w_eco153055, w_eco153056, w_eco153057, w_eco153058, w_eco153059, w_eco153060, w_eco153061, w_eco153062, w_eco153063, w_eco153064, w_eco153065, w_eco153066, w_eco153067, w_eco153068, w_eco153069, w_eco153070, w_eco153071, w_eco153072, w_eco153073, w_eco153074, w_eco153075, w_eco153076, w_eco153077, w_eco153078, w_eco153079, w_eco153080, w_eco153081, w_eco153082, w_eco153083, w_eco153084, w_eco153085, w_eco153086, w_eco153087, w_eco153088, w_eco153089, w_eco153090, w_eco153091, w_eco153092, w_eco153093, w_eco153094, w_eco153095, w_eco153096, w_eco153097, w_eco153098, w_eco153099, w_eco153100, w_eco153101, w_eco153102, w_eco153103, w_eco153104, w_eco153105, w_eco153106, w_eco153107, w_eco153108, w_eco153109, w_eco153110, w_eco153111, w_eco153112, w_eco153113, w_eco153114, w_eco153115, w_eco153116, w_eco153117, w_eco153118, w_eco153119, w_eco153120, w_eco153121, w_eco153122, w_eco153123, w_eco153124, w_eco153125, w_eco153126, w_eco153127, w_eco153128, w_eco153129, w_eco153130, w_eco153131, w_eco153132, w_eco153133, w_eco153134, w_eco153135, w_eco153136, w_eco153137, w_eco153138, w_eco153139, w_eco153140, w_eco153141, w_eco153142, w_eco153143, w_eco153144, w_eco153145, w_eco153146, w_eco153147, w_eco153148, w_eco153149, w_eco153150, w_eco153151, w_eco153152, w_eco153153, w_eco153154, w_eco153155, w_eco153156, w_eco153157, w_eco153158, w_eco153159, w_eco153160, w_eco153161, w_eco153162, w_eco153163, w_eco153164, w_eco153165, w_eco153166, w_eco153167, w_eco153168, w_eco153169, w_eco153170, w_eco153171, w_eco153172, w_eco153173, w_eco153174, w_eco153175, w_eco153176, w_eco153177, w_eco153178, w_eco153179, w_eco153180, w_eco153181, w_eco153182, w_eco153183, w_eco153184, w_eco153185, w_eco153186, w_eco153187, w_eco153188, w_eco153189, w_eco153190, w_eco153191, w_eco153192, w_eco153193, w_eco153194, w_eco153195, w_eco153196, w_eco153197, w_eco153198, w_eco153199, w_eco153200, w_eco153201, w_eco153202, w_eco153203, w_eco153204, w_eco153205, w_eco153206, w_eco153207, w_eco153208, w_eco153209, w_eco153210, w_eco153211, w_eco153212, w_eco153213, w_eco153214, w_eco153215, w_eco153216, w_eco153217, w_eco153218, w_eco153219, w_eco153220, w_eco153221, w_eco153222, w_eco153223, w_eco153224, w_eco153225, w_eco153226, w_eco153227, w_eco153228, w_eco153229, w_eco153230, w_eco153231, w_eco153232, w_eco153233, w_eco153234, w_eco153235, w_eco153236, w_eco153237, w_eco153238, w_eco153239, w_eco153240, w_eco153241, w_eco153242, w_eco153243, w_eco153244, w_eco153245, w_eco153246, w_eco153247, w_eco153248, w_eco153249, w_eco153250, w_eco153251, w_eco153252, w_eco153253, w_eco153254, w_eco153255, w_eco153256, w_eco153257, w_eco153258, w_eco153259, w_eco153260, w_eco153261, w_eco153262, w_eco153263, w_eco153264, w_eco153265, w_eco153266, w_eco153267, w_eco153268, w_eco153269, w_eco153270, w_eco153271, w_eco153272, w_eco153273, w_eco153274, w_eco153275, w_eco153276, w_eco153277, w_eco153278, w_eco153279, w_eco153280, w_eco153281, w_eco153282, w_eco153283, w_eco153284, w_eco153285, w_eco153286, w_eco153287, w_eco153288, w_eco153289, w_eco153290, w_eco153291, w_eco153292, w_eco153293, w_eco153294, w_eco153295, w_eco153296, w_eco153297, w_eco153298, w_eco153299, w_eco153300, w_eco153301, w_eco153302, w_eco153303, w_eco153304, w_eco153305, w_eco153306, w_eco153307, w_eco153308, w_eco153309, w_eco153310, w_eco153311, w_eco153312, w_eco153313, w_eco153314, w_eco153315, w_eco153316, w_eco153317, w_eco153318, w_eco153319, w_eco153320, w_eco153321, w_eco153322, w_eco153323, w_eco153324, w_eco153325, w_eco153326, w_eco153327, w_eco153328, w_eco153329, w_eco153330, w_eco153331, w_eco153332, w_eco153333, w_eco153334, w_eco153335, w_eco153336, w_eco153337, w_eco153338, w_eco153339, w_eco153340, w_eco153341, w_eco153342, w_eco153343, w_eco153344, w_eco153345, w_eco153346, w_eco153347, w_eco153348, w_eco153349, w_eco153350, w_eco153351, w_eco153352, w_eco153353, w_eco153354, w_eco153355, w_eco153356, w_eco153357, w_eco153358, w_eco153359, w_eco153360, w_eco153361, w_eco153362, w_eco153363, w_eco153364, w_eco153365, w_eco153366, w_eco153367, w_eco153368, w_eco153369, w_eco153370, w_eco153371, w_eco153372, w_eco153373, w_eco153374, w_eco153375, w_eco153376, w_eco153377, w_eco153378, w_eco153379, w_eco153380, w_eco153381, w_eco153382, w_eco153383, w_eco153384, w_eco153385, w_eco153386, w_eco153387, w_eco153388, w_eco153389, w_eco153390, w_eco153391, w_eco153392, w_eco153393, w_eco153394, w_eco153395, w_eco153396, w_eco153397, w_eco153398, w_eco153399, w_eco153400, w_eco153401, w_eco153402, w_eco153403, w_eco153404, w_eco153405, w_eco153406, w_eco153407, w_eco153408, w_eco153409, w_eco153410, w_eco153411, w_eco153412, w_eco153413, w_eco153414, w_eco153415, w_eco153416, w_eco153417, w_eco153418, w_eco153419, w_eco153420, w_eco153421, w_eco153422, w_eco153423, w_eco153424, w_eco153425, w_eco153426, w_eco153427, w_eco153428, w_eco153429, w_eco153430, w_eco153431, w_eco153432, w_eco153433, w_eco153434, w_eco153435, w_eco153436, w_eco153437, w_eco153438, w_eco153439, w_eco153440, w_eco153441, w_eco153442, w_eco153443, w_eco153444, w_eco153445, w_eco153446, w_eco153447, w_eco153448, w_eco153449, w_eco153450, w_eco153451, w_eco153452, w_eco153453, w_eco153454, w_eco153455, w_eco153456, w_eco153457, w_eco153458, w_eco153459, w_eco153460, w_eco153461, w_eco153462, w_eco153463, w_eco153464, w_eco153465, w_eco153466, w_eco153467, w_eco153468, w_eco153469, w_eco153470, w_eco153471, w_eco153472, w_eco153473, w_eco153474, w_eco153475, w_eco153476, w_eco153477, w_eco153478, w_eco153479, w_eco153480, w_eco153481, w_eco153482, w_eco153483, w_eco153484, w_eco153485, w_eco153486, w_eco153487, w_eco153488, w_eco153489, w_eco153490, w_eco153491, w_eco153492, w_eco153493, w_eco153494, w_eco153495, w_eco153496, w_eco153497, w_eco153498, w_eco153499, w_eco153500, w_eco153501, w_eco153502, w_eco153503, w_eco153504, w_eco153505, w_eco153506, w_eco153507, w_eco153508, w_eco153509, w_eco153510, w_eco153511, w_eco153512, w_eco153513, w_eco153514, w_eco153515, w_eco153516, w_eco153517, w_eco153518, w_eco153519, w_eco153520, w_eco153521, w_eco153522, w_eco153523, w_eco153524, w_eco153525, w_eco153526, w_eco153527, w_eco153528, w_eco153529, w_eco153530, w_eco153531, w_eco153532, w_eco153533, w_eco153534, w_eco153535, w_eco153536, w_eco153537, w_eco153538, w_eco153539, w_eco153540, w_eco153541, w_eco153542, w_eco153543, w_eco153544, w_eco153545, w_eco153546, w_eco153547, w_eco153548, w_eco153549, w_eco153550, w_eco153551, w_eco153552, w_eco153553, w_eco153554, w_eco153555, w_eco153556, w_eco153557, w_eco153558, w_eco153559, w_eco153560, w_eco153561, w_eco153562, w_eco153563, w_eco153564, w_eco153565, w_eco153566, w_eco153567, w_eco153568, w_eco153569, w_eco153570, w_eco153571, w_eco153572, w_eco153573, w_eco153574, w_eco153575, w_eco153576, w_eco153577, w_eco153578, w_eco153579, w_eco153580, w_eco153581, w_eco153582, w_eco153583, w_eco153584, w_eco153585, w_eco153586, w_eco153587, w_eco153588, w_eco153589, w_eco153590, w_eco153591, w_eco153592, w_eco153593, w_eco153594, w_eco153595, w_eco153596, w_eco153597, w_eco153598, w_eco153599, w_eco153600, w_eco153601, w_eco153602, w_eco153603, w_eco153604, w_eco153605, w_eco153606, w_eco153607, w_eco153608, w_eco153609, w_eco153610, w_eco153611, w_eco153612, w_eco153613, w_eco153614, w_eco153615, w_eco153616, w_eco153617, w_eco153618, w_eco153619, w_eco153620, w_eco153621, w_eco153622, w_eco153623, w_eco153624, w_eco153625, w_eco153626, w_eco153627, w_eco153628, w_eco153629, w_eco153630, w_eco153631, w_eco153632, w_eco153633, w_eco153634, w_eco153635, w_eco153636, w_eco153637, w_eco153638, w_eco153639, w_eco153640, w_eco153641, w_eco153642, w_eco153643, w_eco153644, w_eco153645, w_eco153646, w_eco153647, w_eco153648, w_eco153649, w_eco153650, w_eco153651, w_eco153652, w_eco153653, w_eco153654, w_eco153655, w_eco153656, w_eco153657, w_eco153658, w_eco153659, w_eco153660, w_eco153661, w_eco153662, w_eco153663, w_eco153664, w_eco153665, w_eco153666, w_eco153667, w_eco153668, w_eco153669, w_eco153670, w_eco153671, w_eco153672, w_eco153673, w_eco153674, w_eco153675, w_eco153676, w_eco153677, w_eco153678, w_eco153679, w_eco153680, w_eco153681, w_eco153682, w_eco153683, w_eco153684, w_eco153685, w_eco153686, w_eco153687, w_eco153688, w_eco153689, w_eco153690, w_eco153691, w_eco153692, w_eco153693, w_eco153694, w_eco153695, w_eco153696, w_eco153697, w_eco153698, w_eco153699, w_eco153700, w_eco153701, w_eco153702, w_eco153703, w_eco153704, w_eco153705, w_eco153706, w_eco153707, w_eco153708, w_eco153709, w_eco153710, w_eco153711, w_eco153712, w_eco153713, w_eco153714, w_eco153715, w_eco153716, w_eco153717, w_eco153718, w_eco153719, w_eco153720, w_eco153721, w_eco153722, w_eco153723, w_eco153724, w_eco153725, w_eco153726, w_eco153727, w_eco153728, w_eco153729, w_eco153730, w_eco153731, w_eco153732, w_eco153733, w_eco153734, w_eco153735, w_eco153736, w_eco153737, w_eco153738, w_eco153739, w_eco153740, w_eco153741, w_eco153742, w_eco153743, w_eco153744, w_eco153745, w_eco153746, w_eco153747, w_eco153748, w_eco153749, w_eco153750, w_eco153751, w_eco153752, w_eco153753, w_eco153754, w_eco153755, w_eco153756, w_eco153757, w_eco153758, w_eco153759, w_eco153760, w_eco153761, w_eco153762, w_eco153763, w_eco153764, w_eco153765, w_eco153766, w_eco153767, w_eco153768, w_eco153769, w_eco153770, w_eco153771, w_eco153772, w_eco153773, w_eco153774, w_eco153775, w_eco153776, w_eco153777, w_eco153778, w_eco153779, w_eco153780, w_eco153781, w_eco153782, w_eco153783, w_eco153784, w_eco153785, w_eco153786, w_eco153787, w_eco153788, w_eco153789, w_eco153790, w_eco153791, w_eco153792, w_eco153793, w_eco153794, w_eco153795, w_eco153796, w_eco153797, w_eco153798, w_eco153799, w_eco153800, w_eco153801, w_eco153802, w_eco153803, w_eco153804, w_eco153805, w_eco153806, w_eco153807, w_eco153808, w_eco153809, w_eco153810, w_eco153811, w_eco153812, w_eco153813, w_eco153814, w_eco153815, w_eco153816, w_eco153817, w_eco153818, w_eco153819, w_eco153820, w_eco153821, w_eco153822, w_eco153823, w_eco153824, w_eco153825, w_eco153826, w_eco153827, w_eco153828, w_eco153829, w_eco153830, w_eco153831, w_eco153832, w_eco153833, w_eco153834, w_eco153835, w_eco153836, w_eco153837, w_eco153838, w_eco153839, w_eco153840, w_eco153841, w_eco153842, w_eco153843, w_eco153844, w_eco153845, w_eco153846, w_eco153847, w_eco153848, w_eco153849, w_eco153850, w_eco153851, w_eco153852, w_eco153853, w_eco153854, w_eco153855, w_eco153856, w_eco153857, w_eco153858, w_eco153859, w_eco153860, w_eco153861, w_eco153862, w_eco153863, w_eco153864, w_eco153865, w_eco153866, w_eco153867, w_eco153868, w_eco153869, w_eco153870, w_eco153871, w_eco153872, w_eco153873, w_eco153874, w_eco153875, w_eco153876, w_eco153877, w_eco153878, w_eco153879, w_eco153880, w_eco153881, w_eco153882, w_eco153883, w_eco153884, w_eco153885, w_eco153886, w_eco153887, w_eco153888, w_eco153889, w_eco153890, w_eco153891, w_eco153892, w_eco153893, w_eco153894, w_eco153895, w_eco153896, w_eco153897, w_eco153898, w_eco153899, w_eco153900, w_eco153901, w_eco153902, w_eco153903, w_eco153904, w_eco153905, w_eco153906, w_eco153907, w_eco153908, w_eco153909, w_eco153910, w_eco153911, w_eco153912, w_eco153913, w_eco153914, w_eco153915, w_eco153916, w_eco153917, w_eco153918, w_eco153919, w_eco153920, w_eco153921, w_eco153922, w_eco153923, w_eco153924, w_eco153925, w_eco153926, w_eco153927, w_eco153928, w_eco153929, w_eco153930, w_eco153931, w_eco153932, w_eco153933, w_eco153934, w_eco153935, w_eco153936, w_eco153937, w_eco153938, w_eco153939, w_eco153940, w_eco153941, w_eco153942, w_eco153943, w_eco153944, w_eco153945, w_eco153946, w_eco153947, w_eco153948, w_eco153949, w_eco153950, w_eco153951, w_eco153952, w_eco153953, w_eco153954, w_eco153955, w_eco153956, w_eco153957, w_eco153958, w_eco153959, w_eco153960, w_eco153961, w_eco153962, w_eco153963, w_eco153964, w_eco153965, w_eco153966, w_eco153967, w_eco153968, w_eco153969, w_eco153970, w_eco153971, w_eco153972, w_eco153973, w_eco153974, w_eco153975, w_eco153976, w_eco153977, w_eco153978, w_eco153979, w_eco153980, w_eco153981, w_eco153982, w_eco153983, w_eco153984, w_eco153985, w_eco153986, w_eco153987, w_eco153988, w_eco153989, w_eco153990, w_eco153991, w_eco153992, w_eco153993, w_eco153994, w_eco153995, w_eco153996, w_eco153997, w_eco153998, w_eco153999, w_eco154000, w_eco154001, w_eco154002, w_eco154003, w_eco154004, w_eco154005, w_eco154006, w_eco154007, w_eco154008, w_eco154009, w_eco154010, w_eco154011, w_eco154012, w_eco154013, w_eco154014, w_eco154015, w_eco154016, w_eco154017, w_eco154018, w_eco154019, w_eco154020, w_eco154021, w_eco154022, w_eco154023, w_eco154024, w_eco154025, w_eco154026, w_eco154027, w_eco154028, w_eco154029, w_eco154030, w_eco154031, w_eco154032, w_eco154033, w_eco154034, w_eco154035, w_eco154036, w_eco154037, w_eco154038, w_eco154039, w_eco154040, w_eco154041, w_eco154042, w_eco154043, w_eco154044, w_eco154045, w_eco154046, w_eco154047, w_eco154048, w_eco154049, w_eco154050, w_eco154051, w_eco154052, w_eco154053, w_eco154054, w_eco154055, w_eco154056, w_eco154057, w_eco154058, w_eco154059, w_eco154060, w_eco154061, w_eco154062, w_eco154063, w_eco154064, w_eco154065, w_eco154066, w_eco154067, w_eco154068, w_eco154069, w_eco154070, w_eco154071, w_eco154072, w_eco154073, w_eco154074, w_eco154075, w_eco154076, w_eco154077, w_eco154078, w_eco154079, w_eco154080, w_eco154081, w_eco154082, w_eco154083, w_eco154084, w_eco154085, w_eco154086, w_eco154087, w_eco154088, w_eco154089, w_eco154090, w_eco154091, w_eco154092, w_eco154093, w_eco154094, w_eco154095, w_eco154096, w_eco154097, w_eco154098, w_eco154099, w_eco154100, w_eco154101, w_eco154102, w_eco154103, w_eco154104, w_eco154105, w_eco154106, w_eco154107, w_eco154108, w_eco154109, w_eco154110, w_eco154111, w_eco154112, w_eco154113, w_eco154114, w_eco154115, w_eco154116, w_eco154117, w_eco154118, w_eco154119, w_eco154120, w_eco154121, w_eco154122, w_eco154123, w_eco154124, w_eco154125, w_eco154126, w_eco154127, w_eco154128, w_eco154129, w_eco154130, w_eco154131, w_eco154132, w_eco154133, w_eco154134, w_eco154135, w_eco154136, w_eco154137, w_eco154138, w_eco154139, w_eco154140, w_eco154141, w_eco154142, w_eco154143, w_eco154144, w_eco154145, w_eco154146, w_eco154147, w_eco154148, w_eco154149, w_eco154150, w_eco154151, w_eco154152, w_eco154153, w_eco154154, w_eco154155, w_eco154156, w_eco154157, w_eco154158, w_eco154159, w_eco154160, w_eco154161, w_eco154162, w_eco154163, w_eco154164, w_eco154165, w_eco154166, w_eco154167, w_eco154168, w_eco154169, w_eco154170, w_eco154171, w_eco154172, w_eco154173, w_eco154174, w_eco154175, w_eco154176, w_eco154177, w_eco154178, w_eco154179, w_eco154180, w_eco154181, w_eco154182, w_eco154183, w_eco154184, w_eco154185, w_eco154186, w_eco154187, w_eco154188, w_eco154189, w_eco154190, w_eco154191, w_eco154192, w_eco154193, w_eco154194, w_eco154195, w_eco154196, w_eco154197, w_eco154198, w_eco154199, w_eco154200, w_eco154201, w_eco154202, w_eco154203, w_eco154204, w_eco154205, w_eco154206, w_eco154207, w_eco154208, w_eco154209, w_eco154210, w_eco154211, w_eco154212, w_eco154213, w_eco154214, w_eco154215, w_eco154216, w_eco154217, w_eco154218, w_eco154219, w_eco154220, w_eco154221, w_eco154222, w_eco154223, w_eco154224, w_eco154225, w_eco154226, w_eco154227, w_eco154228, w_eco154229, w_eco154230, w_eco154231, w_eco154232, w_eco154233, w_eco154234, w_eco154235, w_eco154236, w_eco154237, w_eco154238, w_eco154239, w_eco154240, w_eco154241, w_eco154242, w_eco154243, w_eco154244, w_eco154245, w_eco154246, w_eco154247, w_eco154248, w_eco154249, w_eco154250, w_eco154251, w_eco154252, w_eco154253, w_eco154254, w_eco154255, w_eco154256, w_eco154257, w_eco154258, w_eco154259, w_eco154260, w_eco154261, w_eco154262, w_eco154263, w_eco154264, w_eco154265, w_eco154266, w_eco154267, w_eco154268, w_eco154269, w_eco154270, w_eco154271, w_eco154272, w_eco154273, w_eco154274, w_eco154275, w_eco154276, w_eco154277, w_eco154278, w_eco154279, w_eco154280, w_eco154281, w_eco154282, w_eco154283, w_eco154284, w_eco154285, w_eco154286, w_eco154287, w_eco154288, w_eco154289, w_eco154290, w_eco154291, w_eco154292, w_eco154293, w_eco154294, w_eco154295, w_eco154296, w_eco154297, w_eco154298, w_eco154299, w_eco154300, w_eco154301, w_eco154302, w_eco154303, w_eco154304, w_eco154305, w_eco154306, w_eco154307, w_eco154308, w_eco154309, w_eco154310, w_eco154311, w_eco154312, w_eco154313, w_eco154314, w_eco154315, w_eco154316, w_eco154317, w_eco154318, w_eco154319, w_eco154320, w_eco154321, w_eco154322, w_eco154323, w_eco154324, w_eco154325, w_eco154326, w_eco154327, w_eco154328, w_eco154329, w_eco154330, w_eco154331, w_eco154332, w_eco154333, w_eco154334, w_eco154335, w_eco154336, w_eco154337, w_eco154338, w_eco154339, w_eco154340, w_eco154341, w_eco154342, w_eco154343, w_eco154344, w_eco154345, w_eco154346, w_eco154347, w_eco154348, w_eco154349, w_eco154350, w_eco154351, w_eco154352, w_eco154353, w_eco154354, w_eco154355, w_eco154356, w_eco154357, w_eco154358, w_eco154359, w_eco154360, w_eco154361, w_eco154362, w_eco154363, w_eco154364, w_eco154365, w_eco154366, w_eco154367, w_eco154368, w_eco154369, w_eco154370, w_eco154371, w_eco154372, w_eco154373, w_eco154374, w_eco154375, w_eco154376, w_eco154377, w_eco154378, w_eco154379, w_eco154380, w_eco154381, w_eco154382, w_eco154383, w_eco154384, w_eco154385, w_eco154386, w_eco154387, w_eco154388, w_eco154389, w_eco154390, w_eco154391, w_eco154392, w_eco154393, w_eco154394, w_eco154395, w_eco154396, w_eco154397, w_eco154398, w_eco154399, w_eco154400, w_eco154401, w_eco154402, w_eco154403, w_eco154404, w_eco154405, w_eco154406, w_eco154407, w_eco154408, w_eco154409, w_eco154410, w_eco154411, w_eco154412, w_eco154413, w_eco154414, w_eco154415, w_eco154416, w_eco154417, w_eco154418, w_eco154419, w_eco154420, w_eco154421, w_eco154422, w_eco154423, w_eco154424, w_eco154425, w_eco154426, w_eco154427, w_eco154428, w_eco154429, w_eco154430, w_eco154431, w_eco154432, w_eco154433, w_eco154434, w_eco154435, w_eco154436, w_eco154437, w_eco154438, w_eco154439, w_eco154440, w_eco154441, w_eco154442, w_eco154443, w_eco154444, w_eco154445, w_eco154446, w_eco154447, w_eco154448, w_eco154449, w_eco154450, w_eco154451, w_eco154452, w_eco154453, w_eco154454, w_eco154455, w_eco154456, w_eco154457, w_eco154458, w_eco154459, w_eco154460, w_eco154461, w_eco154462, w_eco154463, w_eco154464, w_eco154465, w_eco154466, w_eco154467, w_eco154468, w_eco154469, w_eco154470, w_eco154471, w_eco154472, w_eco154473, w_eco154474, w_eco154475, w_eco154476, w_eco154477, w_eco154478, w_eco154479, w_eco154480, w_eco154481, w_eco154482, w_eco154483, w_eco154484, w_eco154485, w_eco154486, w_eco154487, w_eco154488, w_eco154489, w_eco154490, w_eco154491, w_eco154492, w_eco154493, w_eco154494, w_eco154495, w_eco154496, w_eco154497, w_eco154498, w_eco154499, w_eco154500, w_eco154501, w_eco154502, w_eco154503, w_eco154504, w_eco154505, w_eco154506, w_eco154507, w_eco154508, w_eco154509, w_eco154510, w_eco154511, w_eco154512, w_eco154513, w_eco154514, w_eco154515, w_eco154516, w_eco154517, w_eco154518, w_eco154519, w_eco154520, w_eco154521, w_eco154522, w_eco154523, w_eco154524, w_eco154525, w_eco154526, w_eco154527, w_eco154528, w_eco154529, w_eco154530, w_eco154531, w_eco154532, w_eco154533, w_eco154534, w_eco154535, w_eco154536, w_eco154537, w_eco154538, w_eco154539, w_eco154540, w_eco154541, w_eco154542, w_eco154543, w_eco154544, w_eco154545, w_eco154546, w_eco154547, w_eco154548, w_eco154549, w_eco154550, w_eco154551, w_eco154552, w_eco154553, w_eco154554, w_eco154555, w_eco154556, w_eco154557, w_eco154558, w_eco154559, w_eco154560, w_eco154561, w_eco154562, w_eco154563, w_eco154564, w_eco154565, w_eco154566, w_eco154567, w_eco154568, w_eco154569, w_eco154570, w_eco154571, w_eco154572, w_eco154573, w_eco154574, w_eco154575, w_eco154576, w_eco154577, w_eco154578, w_eco154579, w_eco154580, w_eco154581, w_eco154582, w_eco154583, w_eco154584, w_eco154585, w_eco154586, w_eco154587, w_eco154588, w_eco154589, w_eco154590, w_eco154591, w_eco154592, w_eco154593, w_eco154594, w_eco154595, w_eco154596, w_eco154597, w_eco154598, w_eco154599, w_eco154600, w_eco154601, w_eco154602, w_eco154603, w_eco154604, w_eco154605, w_eco154606, w_eco154607, w_eco154608, w_eco154609, w_eco154610, w_eco154611, w_eco154612, w_eco154613, w_eco154614, w_eco154615, w_eco154616, w_eco154617, w_eco154618, w_eco154619, w_eco154620, w_eco154621, w_eco154622, w_eco154623, w_eco154624, w_eco154625, w_eco154626, w_eco154627, w_eco154628, w_eco154629, w_eco154630, w_eco154631, w_eco154632, w_eco154633, w_eco154634, w_eco154635, w_eco154636, w_eco154637, w_eco154638, w_eco154639, w_eco154640, w_eco154641, w_eco154642, w_eco154643, w_eco154644, w_eco154645, w_eco154646, w_eco154647, w_eco154648, w_eco154649, w_eco154650, w_eco154651, w_eco154652, w_eco154653, w_eco154654, w_eco154655, w_eco154656, w_eco154657, w_eco154658, w_eco154659, w_eco154660, w_eco154661, w_eco154662, w_eco154663, w_eco154664, w_eco154665, w_eco154666, w_eco154667, w_eco154668, w_eco154669, w_eco154670, w_eco154671, w_eco154672, w_eco154673, w_eco154674, w_eco154675, w_eco154676, w_eco154677, w_eco154678, w_eco154679, w_eco154680, w_eco154681, w_eco154682, w_eco154683, w_eco154684, w_eco154685, w_eco154686, w_eco154687, w_eco154688, w_eco154689, w_eco154690, w_eco154691, w_eco154692, w_eco154693, w_eco154694, w_eco154695, w_eco154696, w_eco154697, w_eco154698, w_eco154699, w_eco154700, w_eco154701, w_eco154702, w_eco154703, w_eco154704, w_eco154705, w_eco154706, w_eco154707, w_eco154708, w_eco154709, w_eco154710, w_eco154711, w_eco154712, w_eco154713, w_eco154714, w_eco154715, w_eco154716, w_eco154717, w_eco154718, w_eco154719, w_eco154720, w_eco154721, w_eco154722, w_eco154723, w_eco154724, w_eco154725, w_eco154726, w_eco154727, w_eco154728, w_eco154729, w_eco154730, w_eco154731, w_eco154732, w_eco154733, w_eco154734, w_eco154735, w_eco154736, w_eco154737, w_eco154738, w_eco154739, w_eco154740, w_eco154741, w_eco154742, w_eco154743, w_eco154744, w_eco154745, w_eco154746, w_eco154747, w_eco154748, w_eco154749, w_eco154750, w_eco154751, w_eco154752, w_eco154753, w_eco154754, w_eco154755, w_eco154756, w_eco154757, w_eco154758, w_eco154759, w_eco154760, w_eco154761, w_eco154762, w_eco154763, w_eco154764, w_eco154765, w_eco154766, w_eco154767, w_eco154768, w_eco154769, w_eco154770, w_eco154771, w_eco154772, w_eco154773, w_eco154774, w_eco154775, w_eco154776, w_eco154777, w_eco154778, w_eco154779, w_eco154780, w_eco154781, w_eco154782, w_eco154783, w_eco154784, w_eco154785, w_eco154786, w_eco154787, w_eco154788, w_eco154789, w_eco154790, w_eco154791, w_eco154792, w_eco154793, w_eco154794, w_eco154795, w_eco154796, w_eco154797, w_eco154798, w_eco154799, w_eco154800, w_eco154801, w_eco154802, w_eco154803, w_eco154804, w_eco154805, w_eco154806, w_eco154807, w_eco154808, w_eco154809, w_eco154810, w_eco154811, w_eco154812, w_eco154813, w_eco154814, w_eco154815, w_eco154816, w_eco154817, w_eco154818, w_eco154819, w_eco154820, w_eco154821, w_eco154822, w_eco154823, w_eco154824, w_eco154825, w_eco154826, w_eco154827, w_eco154828, w_eco154829, w_eco154830, w_eco154831, w_eco154832, w_eco154833, w_eco154834, w_eco154835, w_eco154836, w_eco154837, w_eco154838, w_eco154839, w_eco154840, w_eco154841, w_eco154842, w_eco154843, w_eco154844, w_eco154845, w_eco154846, w_eco154847, w_eco154848, w_eco154849, w_eco154850, w_eco154851, w_eco154852, w_eco154853, w_eco154854, w_eco154855, w_eco154856, w_eco154857, w_eco154858, w_eco154859, w_eco154860, w_eco154861, w_eco154862, w_eco154863, w_eco154864, w_eco154865, w_eco154866, w_eco154867, w_eco154868, w_eco154869, w_eco154870, w_eco154871, w_eco154872, w_eco154873, w_eco154874, w_eco154875, w_eco154876, w_eco154877, w_eco154878, w_eco154879, w_eco154880, w_eco154881, w_eco154882, w_eco154883, w_eco154884, w_eco154885, w_eco154886, w_eco154887, w_eco154888, w_eco154889, w_eco154890, w_eco154891, w_eco154892, w_eco154893, w_eco154894, w_eco154895, w_eco154896, w_eco154897, w_eco154898, w_eco154899, w_eco154900, w_eco154901, w_eco154902, w_eco154903, w_eco154904, w_eco154905, w_eco154906, w_eco154907, w_eco154908, w_eco154909, w_eco154910, w_eco154911, w_eco154912, w_eco154913, w_eco154914, w_eco154915, w_eco154916, w_eco154917, w_eco154918, w_eco154919, w_eco154920, w_eco154921, w_eco154922, w_eco154923, w_eco154924, w_eco154925, w_eco154926, w_eco154927, w_eco154928, w_eco154929, w_eco154930, w_eco154931, w_eco154932, w_eco154933, w_eco154934, w_eco154935, w_eco154936, w_eco154937, w_eco154938, w_eco154939, w_eco154940, w_eco154941, w_eco154942, w_eco154943, w_eco154944, w_eco154945, w_eco154946, w_eco154947, w_eco154948, w_eco154949, w_eco154950, w_eco154951, w_eco154952, w_eco154953, w_eco154954, w_eco154955, w_eco154956, w_eco154957, w_eco154958, w_eco154959, w_eco154960, w_eco154961, w_eco154962, w_eco154963, w_eco154964, w_eco154965, w_eco154966, w_eco154967, w_eco154968, w_eco154969, w_eco154970, w_eco154971, w_eco154972, w_eco154973, w_eco154974, w_eco154975, w_eco154976, w_eco154977, w_eco154978, w_eco154979, w_eco154980, w_eco154981, w_eco154982, w_eco154983, w_eco154984, w_eco154985, w_eco154986, w_eco154987, w_eco154988, w_eco154989, w_eco154990, w_eco154991, w_eco154992, w_eco154993, w_eco154994, w_eco154995, w_eco154996, w_eco154997, w_eco154998, w_eco154999, w_eco155000, w_eco155001, w_eco155002, w_eco155003, w_eco155004, w_eco155005, w_eco155006, w_eco155007, w_eco155008, w_eco155009, w_eco155010, w_eco155011, w_eco155012, w_eco155013, w_eco155014, w_eco155015, w_eco155016, w_eco155017, w_eco155018, w_eco155019, w_eco155020, w_eco155021, w_eco155022, w_eco155023, w_eco155024, w_eco155025, w_eco155026, w_eco155027, w_eco155028, w_eco155029, w_eco155030, w_eco155031, w_eco155032, w_eco155033, w_eco155034, w_eco155035, w_eco155036, w_eco155037, w_eco155038, w_eco155039, w_eco155040, w_eco155041, w_eco155042, w_eco155043, w_eco155044, w_eco155045, w_eco155046, w_eco155047, w_eco155048, w_eco155049, w_eco155050, w_eco155051, w_eco155052, w_eco155053, w_eco155054, w_eco155055, w_eco155056, w_eco155057, w_eco155058, w_eco155059, w_eco155060, w_eco155061, w_eco155062, w_eco155063, w_eco155064, w_eco155065, w_eco155066, w_eco155067, w_eco155068, w_eco155069, w_eco155070, w_eco155071, w_eco155072, w_eco155073, w_eco155074, w_eco155075, w_eco155076, w_eco155077, w_eco155078, w_eco155079, w_eco155080, w_eco155081, w_eco155082, w_eco155083, w_eco155084, w_eco155085, w_eco155086, w_eco155087, w_eco155088, w_eco155089, w_eco155090, w_eco155091, w_eco155092, w_eco155093, w_eco155094, w_eco155095, w_eco155096, w_eco155097, w_eco155098, w_eco155099, w_eco155100, w_eco155101, w_eco155102, w_eco155103, w_eco155104, w_eco155105, w_eco155106, w_eco155107, w_eco155108, w_eco155109, w_eco155110, w_eco155111, w_eco155112, w_eco155113, w_eco155114, w_eco155115, w_eco155116, w_eco155117, w_eco155118, w_eco155119, w_eco155120, w_eco155121, w_eco155122, w_eco155123, w_eco155124, w_eco155125, w_eco155126, w_eco155127, w_eco155128, w_eco155129, w_eco155130, w_eco155131, w_eco155132, w_eco155133, w_eco155134, w_eco155135, w_eco155136, w_eco155137, w_eco155138, w_eco155139, w_eco155140, w_eco155141, w_eco155142, w_eco155143, w_eco155144, w_eco155145, w_eco155146, w_eco155147, w_eco155148, w_eco155149, w_eco155150, w_eco155151, w_eco155152, w_eco155153, w_eco155154, w_eco155155, w_eco155156, w_eco155157, w_eco155158, w_eco155159, w_eco155160, w_eco155161, w_eco155162, w_eco155163, w_eco155164, w_eco155165, w_eco155166, w_eco155167, w_eco155168, w_eco155169, w_eco155170, w_eco155171, w_eco155172, w_eco155173, w_eco155174, w_eco155175, w_eco155176, w_eco155177, w_eco155178, w_eco155179, w_eco155180, w_eco155181, w_eco155182, w_eco155183, w_eco155184, w_eco155185, w_eco155186, w_eco155187, w_eco155188, w_eco155189, w_eco155190, w_eco155191, w_eco155192, w_eco155193, w_eco155194, w_eco155195, w_eco155196, w_eco155197, w_eco155198, w_eco155199, w_eco155200, w_eco155201, w_eco155202, w_eco155203, w_eco155204, w_eco155205, w_eco155206, w_eco155207, w_eco155208, w_eco155209, w_eco155210, w_eco155211, w_eco155212, w_eco155213, w_eco155214, w_eco155215, w_eco155216, w_eco155217, w_eco155218, w_eco155219, w_eco155220, w_eco155221, w_eco155222, w_eco155223, w_eco155224, w_eco155225, w_eco155226, w_eco155227, w_eco155228, w_eco155229, w_eco155230, w_eco155231, w_eco155232, w_eco155233, w_eco155234, w_eco155235, w_eco155236, w_eco155237, w_eco155238, w_eco155239, w_eco155240, w_eco155241, w_eco155242, w_eco155243, w_eco155244, w_eco155245, w_eco155246, w_eco155247, w_eco155248, w_eco155249, w_eco155250, w_eco155251, w_eco155252, w_eco155253, w_eco155254, w_eco155255, w_eco155256, w_eco155257, w_eco155258, w_eco155259, w_eco155260, w_eco155261, w_eco155262, w_eco155263, w_eco155264, w_eco155265, w_eco155266, w_eco155267, w_eco155268, w_eco155269, w_eco155270, w_eco155271, w_eco155272, w_eco155273, w_eco155274, w_eco155275, w_eco155276, w_eco155277, w_eco155278, w_eco155279, w_eco155280, w_eco155281, w_eco155282, w_eco155283, w_eco155284, w_eco155285, w_eco155286, w_eco155287, w_eco155288, w_eco155289, w_eco155290, w_eco155291, w_eco155292, w_eco155293, w_eco155294, w_eco155295, w_eco155296, w_eco155297, w_eco155298, w_eco155299, w_eco155300, w_eco155301, w_eco155302, w_eco155303, w_eco155304, w_eco155305, w_eco155306, w_eco155307, w_eco155308, w_eco155309, w_eco155310, w_eco155311, w_eco155312, w_eco155313, w_eco155314, w_eco155315, w_eco155316, w_eco155317, w_eco155318, w_eco155319, w_eco155320, w_eco155321, w_eco155322, w_eco155323, w_eco155324, w_eco155325, w_eco155326, w_eco155327, w_eco155328, w_eco155329, w_eco155330, w_eco155331, w_eco155332, w_eco155333, w_eco155334, w_eco155335, w_eco155336, w_eco155337, w_eco155338, w_eco155339, w_eco155340, w_eco155341, w_eco155342, w_eco155343, w_eco155344, w_eco155345, w_eco155346, w_eco155347, w_eco155348, w_eco155349, w_eco155350, w_eco155351, w_eco155352, w_eco155353, w_eco155354, w_eco155355, w_eco155356, w_eco155357, w_eco155358, w_eco155359, w_eco155360, w_eco155361, w_eco155362, w_eco155363, w_eco155364, w_eco155365, w_eco155366, w_eco155367, w_eco155368, w_eco155369, w_eco155370, w_eco155371, w_eco155372, w_eco155373, w_eco155374, w_eco155375, w_eco155376, w_eco155377, w_eco155378, w_eco155379, w_eco155380, w_eco155381, w_eco155382, w_eco155383, w_eco155384, w_eco155385, w_eco155386, w_eco155387, w_eco155388, w_eco155389, w_eco155390, w_eco155391, w_eco155392, w_eco155393, w_eco155394, w_eco155395, w_eco155396, w_eco155397, w_eco155398, w_eco155399, w_eco155400, w_eco155401, w_eco155402, w_eco155403, w_eco155404, w_eco155405, w_eco155406, w_eco155407, w_eco155408, w_eco155409, w_eco155410, w_eco155411, w_eco155412, w_eco155413, w_eco155414, w_eco155415, w_eco155416, w_eco155417, w_eco155418, w_eco155419, w_eco155420, w_eco155421, w_eco155422, w_eco155423, w_eco155424, w_eco155425, w_eco155426, w_eco155427, w_eco155428, w_eco155429, w_eco155430, w_eco155431, w_eco155432, w_eco155433, w_eco155434, w_eco155435, w_eco155436, w_eco155437, w_eco155438, w_eco155439, w_eco155440, w_eco155441, w_eco155442, w_eco155443, w_eco155444, w_eco155445, w_eco155446, w_eco155447, w_eco155448, w_eco155449, w_eco155450, w_eco155451, w_eco155452, w_eco155453, w_eco155454, w_eco155455, w_eco155456, w_eco155457, w_eco155458, w_eco155459, w_eco155460, w_eco155461, w_eco155462, w_eco155463, w_eco155464, w_eco155465, w_eco155466, w_eco155467, w_eco155468, w_eco155469, w_eco155470, w_eco155471, w_eco155472, w_eco155473, w_eco155474, w_eco155475, w_eco155476, w_eco155477, w_eco155478, w_eco155479, w_eco155480, w_eco155481, w_eco155482, w_eco155483, w_eco155484, w_eco155485, w_eco155486, w_eco155487, w_eco155488, w_eco155489, w_eco155490, w_eco155491, w_eco155492, w_eco155493, w_eco155494, w_eco155495, w_eco155496, w_eco155497, w_eco155498, w_eco155499, w_eco155500, w_eco155501, w_eco155502, w_eco155503, w_eco155504, w_eco155505, w_eco155506, w_eco155507, w_eco155508, w_eco155509, w_eco155510, w_eco155511, w_eco155512, w_eco155513, w_eco155514, w_eco155515, w_eco155516, w_eco155517, w_eco155518, w_eco155519, w_eco155520, w_eco155521, w_eco155522, w_eco155523, w_eco155524, w_eco155525, w_eco155526, w_eco155527, w_eco155528, w_eco155529, w_eco155530, w_eco155531, w_eco155532, w_eco155533, w_eco155534, w_eco155535, w_eco155536, w_eco155537, w_eco155538, w_eco155539, w_eco155540, w_eco155541, w_eco155542, w_eco155543, w_eco155544, w_eco155545, w_eco155546, w_eco155547, w_eco155548, w_eco155549, w_eco155550, w_eco155551, w_eco155552, w_eco155553, w_eco155554, w_eco155555, w_eco155556, w_eco155557, w_eco155558, w_eco155559, w_eco155560, w_eco155561, w_eco155562, w_eco155563, w_eco155564, w_eco155565, w_eco155566, w_eco155567, w_eco155568, w_eco155569, w_eco155570, w_eco155571, w_eco155572, w_eco155573, w_eco155574, w_eco155575, w_eco155576, w_eco155577, w_eco155578, w_eco155579, w_eco155580, w_eco155581, w_eco155582, w_eco155583, w_eco155584, w_eco155585, w_eco155586, w_eco155587, w_eco155588, w_eco155589, w_eco155590, w_eco155591, w_eco155592, w_eco155593, w_eco155594, w_eco155595, w_eco155596, w_eco155597, w_eco155598, w_eco155599, w_eco155600, w_eco155601, w_eco155602, w_eco155603, w_eco155604, w_eco155605, w_eco155606, w_eco155607, w_eco155608, w_eco155609, w_eco155610, w_eco155611, w_eco155612, w_eco155613, w_eco155614, w_eco155615, w_eco155616, w_eco155617, w_eco155618, w_eco155619, w_eco155620, w_eco155621, w_eco155622, w_eco155623, w_eco155624, w_eco155625, w_eco155626, w_eco155627, w_eco155628, w_eco155629, w_eco155630, w_eco155631, w_eco155632, w_eco155633, w_eco155634, w_eco155635, w_eco155636, w_eco155637, w_eco155638, w_eco155639, w_eco155640, w_eco155641, w_eco155642, w_eco155643, w_eco155644, w_eco155645, w_eco155646, w_eco155647, w_eco155648, w_eco155649, w_eco155650, w_eco155651, w_eco155652, w_eco155653, w_eco155654, w_eco155655, w_eco155656, w_eco155657, w_eco155658, w_eco155659, w_eco155660, w_eco155661, w_eco155662, w_eco155663, w_eco155664, w_eco155665, w_eco155666, w_eco155667, w_eco155668, w_eco155669, w_eco155670, w_eco155671, w_eco155672, w_eco155673, w_eco155674, w_eco155675, w_eco155676, w_eco155677, w_eco155678, w_eco155679, w_eco155680, w_eco155681, w_eco155682, w_eco155683, w_eco155684, w_eco155685, w_eco155686, w_eco155687, w_eco155688, w_eco155689, w_eco155690, w_eco155691, w_eco155692, w_eco155693, w_eco155694, w_eco155695, w_eco155696, w_eco155697, w_eco155698, w_eco155699, w_eco155700, w_eco155701, w_eco155702, w_eco155703, w_eco155704, w_eco155705, w_eco155706, w_eco155707, w_eco155708, w_eco155709, w_eco155710, w_eco155711, w_eco155712, w_eco155713, w_eco155714, w_eco155715, w_eco155716, w_eco155717, w_eco155718, w_eco155719, w_eco155720, w_eco155721, w_eco155722, w_eco155723, w_eco155724, w_eco155725, w_eco155726, w_eco155727, w_eco155728, w_eco155729, w_eco155730, w_eco155731, w_eco155732, w_eco155733, w_eco155734, w_eco155735, w_eco155736, w_eco155737, w_eco155738, w_eco155739, w_eco155740, w_eco155741, w_eco155742, w_eco155743, w_eco155744, w_eco155745, w_eco155746, w_eco155747, w_eco155748, w_eco155749, w_eco155750, w_eco155751, w_eco155752, w_eco155753, w_eco155754, w_eco155755, w_eco155756, w_eco155757, w_eco155758, w_eco155759, w_eco155760, w_eco155761, w_eco155762, w_eco155763, w_eco155764, w_eco155765, w_eco155766, w_eco155767, w_eco155768, w_eco155769, w_eco155770, w_eco155771, w_eco155772, w_eco155773, w_eco155774, w_eco155775, w_eco155776, w_eco155777, w_eco155778, w_eco155779, w_eco155780, w_eco155781, w_eco155782, w_eco155783, w_eco155784, w_eco155785, w_eco155786, w_eco155787, w_eco155788, w_eco155789, w_eco155790, w_eco155791, w_eco155792, w_eco155793, w_eco155794, w_eco155795, w_eco155796, w_eco155797, w_eco155798, w_eco155799, w_eco155800, w_eco155801, w_eco155802, w_eco155803, w_eco155804, w_eco155805, w_eco155806, w_eco155807, w_eco155808, w_eco155809, w_eco155810, w_eco155811, w_eco155812, w_eco155813, w_eco155814, w_eco155815, w_eco155816, w_eco155817, w_eco155818, w_eco155819, w_eco155820, w_eco155821, w_eco155822, w_eco155823, w_eco155824, w_eco155825, w_eco155826, w_eco155827, w_eco155828, w_eco155829, w_eco155830, w_eco155831, w_eco155832, w_eco155833, w_eco155834, w_eco155835, w_eco155836, w_eco155837, w_eco155838, w_eco155839, w_eco155840, w_eco155841, w_eco155842, w_eco155843, w_eco155844, w_eco155845, w_eco155846, w_eco155847, w_eco155848, w_eco155849, w_eco155850, w_eco155851, w_eco155852, w_eco155853, w_eco155854, w_eco155855, w_eco155856, w_eco155857, w_eco155858, w_eco155859, w_eco155860, w_eco155861, w_eco155862, w_eco155863, w_eco155864, w_eco155865, w_eco155866, w_eco155867, w_eco155868, w_eco155869, w_eco155870, w_eco155871, w_eco155872, w_eco155873, w_eco155874, w_eco155875, w_eco155876, w_eco155877, w_eco155878, w_eco155879, w_eco155880, w_eco155881, w_eco155882, w_eco155883, w_eco155884, w_eco155885, w_eco155886, w_eco155887, w_eco155888, w_eco155889, w_eco155890, w_eco155891, w_eco155892, w_eco155893, w_eco155894, w_eco155895, w_eco155896, w_eco155897, w_eco155898, w_eco155899, w_eco155900, w_eco155901, w_eco155902, w_eco155903, w_eco155904, w_eco155905, w_eco155906, w_eco155907, w_eco155908, w_eco155909, w_eco155910, w_eco155911, w_eco155912, w_eco155913, w_eco155914, w_eco155915, w_eco155916, w_eco155917, w_eco155918, w_eco155919, w_eco155920, w_eco155921, w_eco155922, w_eco155923, w_eco155924, w_eco155925, w_eco155926, w_eco155927, w_eco155928, w_eco155929, w_eco155930, w_eco155931, w_eco155932, w_eco155933, w_eco155934, w_eco155935, w_eco155936, w_eco155937, w_eco155938, w_eco155939, w_eco155940, w_eco155941, w_eco155942, w_eco155943, w_eco155944, w_eco155945, w_eco155946, w_eco155947, w_eco155948, w_eco155949, w_eco155950, w_eco155951, w_eco155952, w_eco155953, w_eco155954, w_eco155955, w_eco155956, w_eco155957, w_eco155958, w_eco155959, w_eco155960, w_eco155961, w_eco155962, w_eco155963, w_eco155964, w_eco155965, w_eco155966, w_eco155967, w_eco155968, w_eco155969, w_eco155970, w_eco155971, w_eco155972, w_eco155973, w_eco155974, w_eco155975, w_eco155976, w_eco155977, w_eco155978, w_eco155979, w_eco155980, w_eco155981, w_eco155982, w_eco155983, w_eco155984, w_eco155985, w_eco155986, w_eco155987, w_eco155988, w_eco155989, w_eco155990, w_eco155991, w_eco155992, w_eco155993, w_eco155994, w_eco155995, w_eco155996, w_eco155997, w_eco155998, w_eco155999, w_eco156000, w_eco156001, w_eco156002, w_eco156003, w_eco156004, w_eco156005, w_eco156006, w_eco156007, w_eco156008, w_eco156009, w_eco156010, w_eco156011, w_eco156012, w_eco156013, w_eco156014, w_eco156015, w_eco156016, w_eco156017, w_eco156018, w_eco156019, w_eco156020, w_eco156021, w_eco156022, w_eco156023, w_eco156024, w_eco156025, w_eco156026, w_eco156027, w_eco156028, w_eco156029, w_eco156030, w_eco156031, w_eco156032, w_eco156033, w_eco156034, w_eco156035, w_eco156036, w_eco156037, w_eco156038, w_eco156039, w_eco156040, w_eco156041, w_eco156042, w_eco156043, w_eco156044, w_eco156045, w_eco156046, w_eco156047, w_eco156048, w_eco156049, w_eco156050, w_eco156051, w_eco156052, w_eco156053, w_eco156054, w_eco156055, w_eco156056, w_eco156057, w_eco156058, w_eco156059, w_eco156060, w_eco156061, w_eco156062, w_eco156063, w_eco156064, w_eco156065, w_eco156066, w_eco156067, w_eco156068, w_eco156069, w_eco156070, w_eco156071, w_eco156072, w_eco156073, w_eco156074, w_eco156075, w_eco156076, w_eco156077, w_eco156078, w_eco156079, w_eco156080, w_eco156081, w_eco156082, w_eco156083, w_eco156084, w_eco156085, w_eco156086, w_eco156087, w_eco156088, w_eco156089, w_eco156090, w_eco156091, w_eco156092, w_eco156093, w_eco156094, w_eco156095, w_eco156096, w_eco156097, w_eco156098, w_eco156099, w_eco156100, w_eco156101, w_eco156102, w_eco156103, w_eco156104, w_eco156105, w_eco156106, w_eco156107, w_eco156108, w_eco156109, w_eco156110, w_eco156111, w_eco156112, w_eco156113, w_eco156114, w_eco156115, w_eco156116, w_eco156117, w_eco156118, w_eco156119, w_eco156120, w_eco156121, w_eco156122, w_eco156123, w_eco156124, w_eco156125, w_eco156126, w_eco156127, w_eco156128, w_eco156129, w_eco156130, w_eco156131, w_eco156132, w_eco156133, w_eco156134, w_eco156135, w_eco156136, w_eco156137, w_eco156138, w_eco156139, w_eco156140, w_eco156141, w_eco156142, w_eco156143, w_eco156144, w_eco156145, w_eco156146, w_eco156147, w_eco156148, w_eco156149, w_eco156150, w_eco156151, w_eco156152, w_eco156153, w_eco156154, w_eco156155, w_eco156156, w_eco156157, w_eco156158, w_eco156159, w_eco156160, w_eco156161, w_eco156162, w_eco156163, w_eco156164, w_eco156165, w_eco156166, w_eco156167, w_eco156168, w_eco156169, w_eco156170, w_eco156171, w_eco156172, w_eco156173, w_eco156174, w_eco156175, w_eco156176, w_eco156177, w_eco156178, w_eco156179, w_eco156180, w_eco156181, w_eco156182, w_eco156183, w_eco156184, w_eco156185, w_eco156186, w_eco156187, w_eco156188, w_eco156189, w_eco156190, w_eco156191, w_eco156192, w_eco156193, w_eco156194, w_eco156195, w_eco156196, w_eco156197, w_eco156198, w_eco156199, w_eco156200, w_eco156201, w_eco156202, w_eco156203, w_eco156204, w_eco156205, w_eco156206, w_eco156207, w_eco156208, w_eco156209, w_eco156210, w_eco156211, w_eco156212, w_eco156213, w_eco156214, w_eco156215, w_eco156216, w_eco156217, w_eco156218, w_eco156219, w_eco156220, w_eco156221, w_eco156222, w_eco156223, w_eco156224, w_eco156225, w_eco156226, w_eco156227, w_eco156228, w_eco156229, w_eco156230, w_eco156231, w_eco156232, w_eco156233, w_eco156234, w_eco156235, w_eco156236, w_eco156237, w_eco156238, w_eco156239, w_eco156240, w_eco156241, w_eco156242, w_eco156243, w_eco156244, w_eco156245, w_eco156246, w_eco156247, w_eco156248, w_eco156249, w_eco156250, w_eco156251, w_eco156252, w_eco156253, w_eco156254, w_eco156255, w_eco156256, w_eco156257, w_eco156258, w_eco156259, w_eco156260, w_eco156261, w_eco156262, w_eco156263, w_eco156264, w_eco156265, w_eco156266, w_eco156267, w_eco156268, w_eco156269, w_eco156270, w_eco156271, w_eco156272, w_eco156273, w_eco156274, w_eco156275, w_eco156276, w_eco156277, w_eco156278, w_eco156279, w_eco156280, w_eco156281, w_eco156282, w_eco156283, w_eco156284, w_eco156285, w_eco156286, w_eco156287, w_eco156288, w_eco156289, w_eco156290, w_eco156291, w_eco156292, w_eco156293, w_eco156294, w_eco156295, w_eco156296, w_eco156297, w_eco156298, w_eco156299, w_eco156300, w_eco156301, w_eco156302, w_eco156303, w_eco156304, w_eco156305, w_eco156306, w_eco156307, w_eco156308, w_eco156309, w_eco156310, w_eco156311, w_eco156312, w_eco156313, w_eco156314, w_eco156315, w_eco156316, w_eco156317, w_eco156318, w_eco156319, w_eco156320, w_eco156321, w_eco156322, w_eco156323, w_eco156324, w_eco156325, w_eco156326, w_eco156327, w_eco156328, w_eco156329, w_eco156330, w_eco156331, w_eco156332, w_eco156333, w_eco156334, w_eco156335, w_eco156336, w_eco156337, w_eco156338, w_eco156339, w_eco156340, w_eco156341, w_eco156342, w_eco156343, w_eco156344, w_eco156345, w_eco156346, w_eco156347, w_eco156348, w_eco156349, w_eco156350, w_eco156351, w_eco156352, w_eco156353, w_eco156354, w_eco156355, w_eco156356, w_eco156357, w_eco156358, w_eco156359, w_eco156360, w_eco156361, w_eco156362, w_eco156363, w_eco156364, w_eco156365, w_eco156366, w_eco156367, w_eco156368, w_eco156369, w_eco156370, w_eco156371, w_eco156372, w_eco156373, w_eco156374, w_eco156375, w_eco156376, w_eco156377, w_eco156378, w_eco156379, w_eco156380, w_eco156381, w_eco156382, w_eco156383, w_eco156384, w_eco156385, w_eco156386, w_eco156387, w_eco156388, w_eco156389, w_eco156390, w_eco156391, w_eco156392, w_eco156393, w_eco156394, w_eco156395, w_eco156396, w_eco156397, w_eco156398, w_eco156399, w_eco156400, w_eco156401, w_eco156402, w_eco156403, w_eco156404, w_eco156405, w_eco156406, w_eco156407, w_eco156408, w_eco156409, w_eco156410, w_eco156411, w_eco156412, w_eco156413, w_eco156414, w_eco156415, w_eco156416, w_eco156417, w_eco156418, w_eco156419, w_eco156420, w_eco156421, w_eco156422, w_eco156423, w_eco156424, w_eco156425, w_eco156426, w_eco156427, w_eco156428, w_eco156429, w_eco156430, w_eco156431, w_eco156432, w_eco156433, w_eco156434, w_eco156435, w_eco156436, w_eco156437, w_eco156438, w_eco156439, w_eco156440, w_eco156441, w_eco156442, w_eco156443, w_eco156444, w_eco156445, w_eco156446, w_eco156447, w_eco156448, w_eco156449, w_eco156450, w_eco156451, w_eco156452, w_eco156453, w_eco156454, w_eco156455, w_eco156456, w_eco156457, w_eco156458, w_eco156459, w_eco156460, w_eco156461, w_eco156462, w_eco156463, w_eco156464, w_eco156465, w_eco156466, w_eco156467, w_eco156468, w_eco156469, w_eco156470, w_eco156471, w_eco156472, w_eco156473, w_eco156474, w_eco156475, w_eco156476, w_eco156477, w_eco156478, w_eco156479, w_eco156480, w_eco156481, w_eco156482, w_eco156483, w_eco156484, w_eco156485, w_eco156486, w_eco156487, w_eco156488, w_eco156489, w_eco156490, w_eco156491, w_eco156492, w_eco156493, w_eco156494, w_eco156495, w_eco156496, w_eco156497, w_eco156498, w_eco156499, w_eco156500, w_eco156501, w_eco156502, w_eco156503, w_eco156504, w_eco156505, w_eco156506, w_eco156507, w_eco156508, w_eco156509, w_eco156510, w_eco156511, w_eco156512, w_eco156513, w_eco156514, w_eco156515, w_eco156516, w_eco156517, w_eco156518, w_eco156519, w_eco156520, w_eco156521, w_eco156522, w_eco156523, w_eco156524, w_eco156525, w_eco156526, w_eco156527, w_eco156528, w_eco156529, w_eco156530, w_eco156531, w_eco156532, w_eco156533, w_eco156534, w_eco156535, w_eco156536, w_eco156537, w_eco156538, w_eco156539, w_eco156540, w_eco156541, w_eco156542, w_eco156543, w_eco156544, w_eco156545, w_eco156546, w_eco156547, w_eco156548, w_eco156549, w_eco156550, w_eco156551, w_eco156552, w_eco156553, w_eco156554, w_eco156555, w_eco156556, w_eco156557, w_eco156558, w_eco156559, w_eco156560, w_eco156561, w_eco156562, w_eco156563, w_eco156564, w_eco156565, w_eco156566, w_eco156567, w_eco156568, w_eco156569, w_eco156570, w_eco156571, w_eco156572, w_eco156573, w_eco156574, w_eco156575, w_eco156576, w_eco156577, w_eco156578, w_eco156579, w_eco156580, w_eco156581, w_eco156582, w_eco156583, w_eco156584, w_eco156585, w_eco156586, w_eco156587, w_eco156588, w_eco156589, w_eco156590, w_eco156591, w_eco156592, w_eco156593, w_eco156594, w_eco156595, w_eco156596, w_eco156597, w_eco156598, w_eco156599, w_eco156600, w_eco156601, w_eco156602, w_eco156603, w_eco156604, w_eco156605, w_eco156606, w_eco156607, w_eco156608, w_eco156609, w_eco156610, w_eco156611, w_eco156612, w_eco156613, w_eco156614, w_eco156615, w_eco156616, w_eco156617, w_eco156618, w_eco156619, w_eco156620, w_eco156621, w_eco156622, w_eco156623, w_eco156624, w_eco156625, w_eco156626, w_eco156627, w_eco156628, w_eco156629, w_eco156630, w_eco156631, w_eco156632, w_eco156633, w_eco156634, w_eco156635, w_eco156636, w_eco156637, w_eco156638, w_eco156639, w_eco156640, w_eco156641, w_eco156642, w_eco156643, w_eco156644, w_eco156645, w_eco156646, w_eco156647, w_eco156648, w_eco156649, w_eco156650, w_eco156651, w_eco156652, w_eco156653, w_eco156654, w_eco156655, w_eco156656, w_eco156657, w_eco156658, w_eco156659, w_eco156660, w_eco156661, w_eco156662, w_eco156663, w_eco156664, w_eco156665, w_eco156666, w_eco156667, w_eco156668, w_eco156669, w_eco156670, w_eco156671, w_eco156672, w_eco156673, w_eco156674, w_eco156675, w_eco156676, w_eco156677, w_eco156678, w_eco156679, w_eco156680, w_eco156681, w_eco156682, w_eco156683, w_eco156684, w_eco156685, w_eco156686, w_eco156687, w_eco156688, w_eco156689, w_eco156690, w_eco156691, w_eco156692, w_eco156693, w_eco156694, w_eco156695, w_eco156696, w_eco156697, w_eco156698, w_eco156699, w_eco156700, w_eco156701, w_eco156702, w_eco156703, w_eco156704, w_eco156705, w_eco156706, w_eco156707, w_eco156708, w_eco156709, w_eco156710, w_eco156711, w_eco156712, w_eco156713, w_eco156714, w_eco156715, w_eco156716, w_eco156717, w_eco156718, w_eco156719, w_eco156720, w_eco156721, w_eco156722, w_eco156723, w_eco156724, w_eco156725, w_eco156726, w_eco156727, w_eco156728, w_eco156729, w_eco156730, w_eco156731, w_eco156732, w_eco156733, w_eco156734, w_eco156735, w_eco156736, w_eco156737, w_eco156738, w_eco156739, w_eco156740, w_eco156741, w_eco156742, w_eco156743, w_eco156744, w_eco156745, w_eco156746, w_eco156747, w_eco156748, w_eco156749, w_eco156750, w_eco156751, w_eco156752, w_eco156753, w_eco156754, w_eco156755, w_eco156756, w_eco156757, w_eco156758, w_eco156759, w_eco156760, w_eco156761, w_eco156762, w_eco156763, w_eco156764, w_eco156765, w_eco156766, w_eco156767, w_eco156768, w_eco156769, w_eco156770, w_eco156771, w_eco156772, w_eco156773, w_eco156774, w_eco156775, w_eco156776, w_eco156777, w_eco156778, w_eco156779, w_eco156780, w_eco156781, w_eco156782, w_eco156783, w_eco156784, w_eco156785, w_eco156786, w_eco156787, w_eco156788, w_eco156789, w_eco156790, w_eco156791, w_eco156792, w_eco156793, w_eco156794, w_eco156795, w_eco156796, w_eco156797, w_eco156798, w_eco156799, w_eco156800, w_eco156801, w_eco156802, w_eco156803, w_eco156804, w_eco156805, w_eco156806, w_eco156807, w_eco156808, w_eco156809, w_eco156810, w_eco156811, w_eco156812, w_eco156813, w_eco156814, w_eco156815, w_eco156816, w_eco156817, w_eco156818, w_eco156819, w_eco156820, w_eco156821, w_eco156822, w_eco156823, w_eco156824, w_eco156825, w_eco156826, w_eco156827, w_eco156828, w_eco156829, w_eco156830, w_eco156831, w_eco156832, w_eco156833, w_eco156834, w_eco156835, w_eco156836, w_eco156837, w_eco156838, w_eco156839, w_eco156840, w_eco156841, w_eco156842, w_eco156843, w_eco156844, w_eco156845, w_eco156846, w_eco156847, w_eco156848, w_eco156849, w_eco156850, w_eco156851, w_eco156852, w_eco156853, w_eco156854, w_eco156855, w_eco156856, w_eco156857, w_eco156858, w_eco156859, w_eco156860, w_eco156861, w_eco156862, w_eco156863, w_eco156864, w_eco156865, w_eco156866, w_eco156867, w_eco156868, w_eco156869, w_eco156870, w_eco156871, w_eco156872, w_eco156873, w_eco156874, w_eco156875, w_eco156876, w_eco156877, w_eco156878, w_eco156879, w_eco156880, w_eco156881, w_eco156882, w_eco156883, w_eco156884, w_eco156885, w_eco156886, w_eco156887, w_eco156888, w_eco156889, w_eco156890, w_eco156891, w_eco156892, w_eco156893, w_eco156894, w_eco156895, w_eco156896, w_eco156897, w_eco156898, w_eco156899, w_eco156900, w_eco156901, w_eco156902, w_eco156903, w_eco156904, w_eco156905, w_eco156906, w_eco156907, w_eco156908, w_eco156909, w_eco156910, w_eco156911, w_eco156912, w_eco156913, w_eco156914, w_eco156915, w_eco156916, w_eco156917, w_eco156918, w_eco156919, w_eco156920, w_eco156921, w_eco156922, w_eco156923, w_eco156924, w_eco156925, w_eco156926, w_eco156927, w_eco156928, w_eco156929, w_eco156930, w_eco156931, w_eco156932, w_eco156933, w_eco156934, w_eco156935, w_eco156936, w_eco156937, w_eco156938, w_eco156939, w_eco156940, w_eco156941, w_eco156942, w_eco156943, w_eco156944, w_eco156945, w_eco156946, w_eco156947, w_eco156948, w_eco156949, w_eco156950, w_eco156951, w_eco156952, w_eco156953, w_eco156954, w_eco156955, w_eco156956, w_eco156957, w_eco156958, w_eco156959, w_eco156960, w_eco156961, w_eco156962, w_eco156963, w_eco156964, w_eco156965, w_eco156966, w_eco156967, w_eco156968, w_eco156969, w_eco156970, w_eco156971, w_eco156972, w_eco156973, w_eco156974, w_eco156975, w_eco156976, w_eco156977, w_eco156978, w_eco156979, w_eco156980, w_eco156981, w_eco156982, w_eco156983, w_eco156984, w_eco156985, w_eco156986, w_eco156987, w_eco156988, w_eco156989, w_eco156990, w_eco156991, w_eco156992, w_eco156993, w_eco156994, w_eco156995, w_eco156996, w_eco156997, w_eco156998, w_eco156999, w_eco157000, w_eco157001, w_eco157002, w_eco157003, w_eco157004, w_eco157005, w_eco157006, w_eco157007, w_eco157008, w_eco157009, w_eco157010, w_eco157011, w_eco157012, w_eco157013, w_eco157014, w_eco157015, w_eco157016, w_eco157017, w_eco157018, w_eco157019, w_eco157020, w_eco157021, w_eco157022, w_eco157023, w_eco157024, w_eco157025, w_eco157026, w_eco157027, w_eco157028, w_eco157029, w_eco157030, w_eco157031, w_eco157032, w_eco157033, w_eco157034, w_eco157035, w_eco157036, w_eco157037, w_eco157038, w_eco157039, w_eco157040, w_eco157041, w_eco157042, w_eco157043, w_eco157044, w_eco157045, w_eco157046, w_eco157047, w_eco157048, w_eco157049, w_eco157050, w_eco157051, w_eco157052, w_eco157053, w_eco157054, w_eco157055, w_eco157056, w_eco157057, w_eco157058, w_eco157059, w_eco157060, w_eco157061, w_eco157062, w_eco157063, w_eco157064, w_eco157065, w_eco157066, w_eco157067, w_eco157068, w_eco157069, w_eco157070, w_eco157071, w_eco157072, w_eco157073, w_eco157074, w_eco157075, w_eco157076, w_eco157077, w_eco157078, w_eco157079, w_eco157080, w_eco157081, w_eco157082, w_eco157083, w_eco157084, w_eco157085, w_eco157086, w_eco157087, w_eco157088, w_eco157089, w_eco157090, w_eco157091, w_eco157092, w_eco157093, w_eco157094, w_eco157095, w_eco157096, w_eco157097, w_eco157098, w_eco157099, w_eco157100, w_eco157101, w_eco157102, w_eco157103, w_eco157104, w_eco157105, w_eco157106, w_eco157107, w_eco157108, w_eco157109, w_eco157110, w_eco157111, w_eco157112, w_eco157113, w_eco157114, w_eco157115, w_eco157116, w_eco157117, w_eco157118, w_eco157119, w_eco157120, w_eco157121, w_eco157122, w_eco157123, w_eco157124, w_eco157125, w_eco157126, w_eco157127, w_eco157128, w_eco157129, w_eco157130, w_eco157131, w_eco157132, w_eco157133, w_eco157134, w_eco157135, w_eco157136, w_eco157137, w_eco157138, w_eco157139, w_eco157140, w_eco157141, w_eco157142, w_eco157143, w_eco157144, w_eco157145, w_eco157146, w_eco157147, w_eco157148, w_eco157149, w_eco157150, w_eco157151, w_eco157152, w_eco157153, w_eco157154, w_eco157155, w_eco157156, w_eco157157, w_eco157158, w_eco157159, w_eco157160, w_eco157161, w_eco157162, w_eco157163, w_eco157164, w_eco157165, w_eco157166, w_eco157167, w_eco157168, w_eco157169, w_eco157170, w_eco157171, w_eco157172, w_eco157173, w_eco157174, w_eco157175, w_eco157176, w_eco157177, w_eco157178, w_eco157179, w_eco157180, w_eco157181, w_eco157182, w_eco157183, w_eco157184, w_eco157185, w_eco157186, w_eco157187, w_eco157188, w_eco157189, w_eco157190, w_eco157191, w_eco157192, w_eco157193, w_eco157194, w_eco157195, w_eco157196, w_eco157197, w_eco157198, w_eco157199, w_eco157200, w_eco157201, w_eco157202, w_eco157203, w_eco157204, w_eco157205, w_eco157206, w_eco157207, w_eco157208, w_eco157209, w_eco157210, w_eco157211, w_eco157212, w_eco157213, w_eco157214, w_eco157215, w_eco157216, w_eco157217, w_eco157218, w_eco157219, w_eco157220, w_eco157221, w_eco157222, w_eco157223, w_eco157224, w_eco157225, w_eco157226, w_eco157227, w_eco157228, w_eco157229, w_eco157230, w_eco157231, w_eco157232, w_eco157233, w_eco157234, w_eco157235, w_eco157236, w_eco157237, w_eco157238, w_eco157239, w_eco157240, w_eco157241, w_eco157242, w_eco157243, w_eco157244, w_eco157245, w_eco157246, w_eco157247, w_eco157248, w_eco157249, w_eco157250, w_eco157251, w_eco157252, w_eco157253, w_eco157254, w_eco157255, w_eco157256, w_eco157257, w_eco157258, w_eco157259, w_eco157260, w_eco157261, w_eco157262, w_eco157263, w_eco157264, w_eco157265, w_eco157266, w_eco157267, w_eco157268, w_eco157269, w_eco157270, w_eco157271, w_eco157272, w_eco157273, w_eco157274, w_eco157275, w_eco157276, w_eco157277, w_eco157278, w_eco157279, w_eco157280, w_eco157281, w_eco157282, w_eco157283, w_eco157284, w_eco157285, w_eco157286, w_eco157287, w_eco157288, w_eco157289, w_eco157290, w_eco157291, w_eco157292, w_eco157293, w_eco157294, w_eco157295, w_eco157296, w_eco157297, w_eco157298, w_eco157299, w_eco157300, w_eco157301, w_eco157302, w_eco157303, w_eco157304, w_eco157305, w_eco157306, w_eco157307, w_eco157308, w_eco157309, w_eco157310, w_eco157311, w_eco157312, w_eco157313, w_eco157314, w_eco157315, w_eco157316, w_eco157317, w_eco157318, w_eco157319, w_eco157320, w_eco157321, w_eco157322, w_eco157323, w_eco157324, w_eco157325, w_eco157326, w_eco157327, w_eco157328, w_eco157329, w_eco157330, w_eco157331, w_eco157332, w_eco157333, w_eco157334, w_eco157335, w_eco157336, w_eco157337, w_eco157338, w_eco157339, w_eco157340, w_eco157341, w_eco157342, w_eco157343, w_eco157344, w_eco157345, w_eco157346, w_eco157347, w_eco157348, w_eco157349, w_eco157350, w_eco157351, w_eco157352, w_eco157353, w_eco157354, w_eco157355, w_eco157356, w_eco157357, w_eco157358, w_eco157359, w_eco157360, w_eco157361, w_eco157362, w_eco157363, w_eco157364, w_eco157365, w_eco157366, w_eco157367, w_eco157368, w_eco157369, w_eco157370, w_eco157371, w_eco157372, w_eco157373, w_eco157374, w_eco157375, w_eco157376, w_eco157377, w_eco157378, w_eco157379, w_eco157380, w_eco157381, w_eco157382, w_eco157383, w_eco157384, w_eco157385, w_eco157386, w_eco157387, w_eco157388, w_eco157389, w_eco157390, w_eco157391, w_eco157392, w_eco157393, w_eco157394, w_eco157395, w_eco157396, w_eco157397, w_eco157398, w_eco157399, w_eco157400, w_eco157401, w_eco157402, w_eco157403, w_eco157404, w_eco157405, w_eco157406, w_eco157407, w_eco157408, w_eco157409, w_eco157410, w_eco157411, w_eco157412, w_eco157413, w_eco157414, w_eco157415, w_eco157416, w_eco157417, w_eco157418, w_eco157419, w_eco157420, w_eco157421, w_eco157422, w_eco157423, w_eco157424, w_eco157425, w_eco157426, w_eco157427, w_eco157428, w_eco157429, w_eco157430, w_eco157431, w_eco157432, w_eco157433, w_eco157434, w_eco157435, w_eco157436, w_eco157437, w_eco157438, w_eco157439, w_eco157440, w_eco157441, w_eco157442, w_eco157443, w_eco157444, w_eco157445, w_eco157446, w_eco157447, w_eco157448, w_eco157449, w_eco157450, w_eco157451, w_eco157452, w_eco157453, w_eco157454, w_eco157455, w_eco157456, w_eco157457, w_eco157458, w_eco157459, w_eco157460, w_eco157461, w_eco157462, w_eco157463, w_eco157464, w_eco157465, w_eco157466, w_eco157467, w_eco157468, w_eco157469, w_eco157470, w_eco157471, w_eco157472, w_eco157473, w_eco157474, w_eco157475, w_eco157476, w_eco157477, w_eco157478, w_eco157479, w_eco157480, w_eco157481, w_eco157482, w_eco157483, w_eco157484, w_eco157485, w_eco157486, w_eco157487, w_eco157488, w_eco157489, w_eco157490, w_eco157491, w_eco157492, w_eco157493, w_eco157494, w_eco157495, w_eco157496, w_eco157497, w_eco157498, w_eco157499, w_eco157500, w_eco157501, w_eco157502, w_eco157503, w_eco157504, w_eco157505, w_eco157506, w_eco157507, w_eco157508, w_eco157509, w_eco157510, w_eco157511, w_eco157512, w_eco157513, w_eco157514, w_eco157515, w_eco157516, w_eco157517, w_eco157518, w_eco157519, w_eco157520, w_eco157521, w_eco157522, w_eco157523, w_eco157524, w_eco157525, w_eco157526, w_eco157527, w_eco157528, w_eco157529, w_eco157530, w_eco157531, w_eco157532, w_eco157533, w_eco157534, w_eco157535, w_eco157536, w_eco157537, w_eco157538, w_eco157539, w_eco157540, w_eco157541, w_eco157542, w_eco157543, w_eco157544, w_eco157545, w_eco157546, w_eco157547, w_eco157548, w_eco157549, w_eco157550, w_eco157551, w_eco157552, w_eco157553, w_eco157554, w_eco157555, w_eco157556, w_eco157557, w_eco157558, w_eco157559, w_eco157560, w_eco157561, w_eco157562, w_eco157563, w_eco157564, w_eco157565, w_eco157566, w_eco157567, w_eco157568, w_eco157569, w_eco157570, w_eco157571, w_eco157572, w_eco157573, w_eco157574, w_eco157575, w_eco157576, w_eco157577, w_eco157578, w_eco157579, w_eco157580, w_eco157581, w_eco157582, w_eco157583, w_eco157584, w_eco157585, w_eco157586, w_eco157587, w_eco157588, w_eco157589, w_eco157590, w_eco157591, w_eco157592, w_eco157593, w_eco157594, w_eco157595, w_eco157596, w_eco157597, w_eco157598, w_eco157599, w_eco157600, w_eco157601, w_eco157602, w_eco157603, w_eco157604, w_eco157605, w_eco157606, w_eco157607, w_eco157608, w_eco157609, w_eco157610, w_eco157611, w_eco157612, w_eco157613, w_eco157614, w_eco157615, w_eco157616, w_eco157617, w_eco157618, w_eco157619, w_eco157620, w_eco157621, w_eco157622, w_eco157623, w_eco157624, w_eco157625, w_eco157626, w_eco157627, w_eco157628, w_eco157629, w_eco157630, w_eco157631, w_eco157632, w_eco157633, w_eco157634, w_eco157635, w_eco157636, w_eco157637, w_eco157638, w_eco157639, w_eco157640, w_eco157641, w_eco157642, w_eco157643, w_eco157644, w_eco157645, w_eco157646, w_eco157647, w_eco157648, w_eco157649, w_eco157650, w_eco157651, w_eco157652, w_eco157653, w_eco157654, w_eco157655, w_eco157656, w_eco157657, w_eco157658, w_eco157659, w_eco157660, w_eco157661, w_eco157662, w_eco157663, w_eco157664, w_eco157665, w_eco157666, w_eco157667, w_eco157668, w_eco157669, w_eco157670, w_eco157671, w_eco157672, w_eco157673, w_eco157674, w_eco157675, w_eco157676, w_eco157677, w_eco157678, w_eco157679, w_eco157680, w_eco157681, w_eco157682, w_eco157683, w_eco157684, w_eco157685, w_eco157686, w_eco157687, w_eco157688, w_eco157689, w_eco157690, w_eco157691, w_eco157692, w_eco157693, w_eco157694, w_eco157695, w_eco157696, w_eco157697, w_eco157698, w_eco157699, w_eco157700, w_eco157701, w_eco157702, w_eco157703, w_eco157704, w_eco157705, w_eco157706, w_eco157707, w_eco157708, w_eco157709, w_eco157710, w_eco157711, w_eco157712, w_eco157713, w_eco157714, w_eco157715, w_eco157716, w_eco157717, w_eco157718, w_eco157719, w_eco157720, w_eco157721, w_eco157722, w_eco157723, w_eco157724, w_eco157725, w_eco157726, w_eco157727, w_eco157728, w_eco157729, w_eco157730, w_eco157731, w_eco157732, w_eco157733, w_eco157734, w_eco157735, w_eco157736, w_eco157737, w_eco157738, w_eco157739, w_eco157740, w_eco157741, w_eco157742, w_eco157743, w_eco157744, w_eco157745, w_eco157746, w_eco157747, w_eco157748, w_eco157749, w_eco157750, w_eco157751, w_eco157752, w_eco157753, w_eco157754, w_eco157755, w_eco157756, w_eco157757, w_eco157758, w_eco157759, w_eco157760, w_eco157761, w_eco157762, w_eco157763, w_eco157764, w_eco157765, w_eco157766, w_eco157767, w_eco157768, w_eco157769, w_eco157770, w_eco157771, w_eco157772, w_eco157773, w_eco157774, w_eco157775, w_eco157776, w_eco157777, w_eco157778, w_eco157779, w_eco157780, w_eco157781, w_eco157782, w_eco157783, w_eco157784, w_eco157785, w_eco157786, w_eco157787, w_eco157788, w_eco157789, w_eco157790, w_eco157791, w_eco157792, w_eco157793, w_eco157794, w_eco157795, w_eco157796, w_eco157797, w_eco157798, w_eco157799, w_eco157800, w_eco157801, w_eco157802, w_eco157803, w_eco157804, w_eco157805, w_eco157806, w_eco157807, w_eco157808, w_eco157809, w_eco157810, w_eco157811, w_eco157812, w_eco157813, w_eco157814, w_eco157815, w_eco157816, w_eco157817, w_eco157818, w_eco157819, w_eco157820, w_eco157821, w_eco157822, w_eco157823, w_eco157824, w_eco157825, w_eco157826, w_eco157827, w_eco157828, w_eco157829, w_eco157830, w_eco157831, w_eco157832, w_eco157833, w_eco157834, w_eco157835, w_eco157836, w_eco157837, w_eco157838, w_eco157839, w_eco157840, w_eco157841, w_eco157842, w_eco157843, w_eco157844, w_eco157845, w_eco157846, w_eco157847, w_eco157848, w_eco157849, w_eco157850, w_eco157851, w_eco157852, w_eco157853, w_eco157854, w_eco157855, w_eco157856, w_eco157857, w_eco157858, w_eco157859, w_eco157860, w_eco157861, w_eco157862, w_eco157863, w_eco157864, w_eco157865, w_eco157866, w_eco157867, w_eco157868, w_eco157869, w_eco157870, w_eco157871, w_eco157872, w_eco157873, w_eco157874, w_eco157875, w_eco157876, w_eco157877, w_eco157878, w_eco157879, w_eco157880, w_eco157881, w_eco157882, w_eco157883, w_eco157884, w_eco157885, w_eco157886, w_eco157887, w_eco157888, w_eco157889, w_eco157890, w_eco157891, w_eco157892, w_eco157893, w_eco157894, w_eco157895, w_eco157896, w_eco157897, w_eco157898, w_eco157899, w_eco157900, w_eco157901, w_eco157902, w_eco157903, w_eco157904, w_eco157905, w_eco157906, w_eco157907, w_eco157908, w_eco157909, w_eco157910, w_eco157911, w_eco157912, w_eco157913, w_eco157914, w_eco157915, w_eco157916, w_eco157917, w_eco157918, w_eco157919, w_eco157920, w_eco157921, w_eco157922, w_eco157923, w_eco157924, w_eco157925, w_eco157926, w_eco157927, w_eco157928, w_eco157929, w_eco157930, w_eco157931, w_eco157932, w_eco157933, w_eco157934, w_eco157935, w_eco157936, w_eco157937, w_eco157938, w_eco157939, w_eco157940, w_eco157941, w_eco157942, w_eco157943, w_eco157944, w_eco157945, w_eco157946, w_eco157947, w_eco157948, w_eco157949, w_eco157950, w_eco157951, w_eco157952, w_eco157953, w_eco157954, w_eco157955, w_eco157956, w_eco157957, w_eco157958, w_eco157959, w_eco157960, w_eco157961, w_eco157962, w_eco157963, w_eco157964, w_eco157965, w_eco157966, w_eco157967, w_eco157968, w_eco157969, w_eco157970, w_eco157971, w_eco157972, w_eco157973, w_eco157974, w_eco157975, w_eco157976, w_eco157977, w_eco157978, w_eco157979, w_eco157980, w_eco157981, w_eco157982, w_eco157983, w_eco157984, w_eco157985, w_eco157986, w_eco157987, w_eco157988, w_eco157989, w_eco157990, w_eco157991, w_eco157992, w_eco157993, w_eco157994, w_eco157995, w_eco157996, w_eco157997, w_eco157998, w_eco157999, w_eco158000, w_eco158001, w_eco158002, w_eco158003, w_eco158004, w_eco158005, w_eco158006, w_eco158007, w_eco158008, w_eco158009, w_eco158010, w_eco158011, w_eco158012, w_eco158013, w_eco158014, w_eco158015, w_eco158016, w_eco158017, w_eco158018, w_eco158019, w_eco158020, w_eco158021, w_eco158022, w_eco158023, w_eco158024, w_eco158025, w_eco158026, w_eco158027, w_eco158028, w_eco158029, w_eco158030, w_eco158031, w_eco158032, w_eco158033, w_eco158034, w_eco158035, w_eco158036, w_eco158037, w_eco158038, w_eco158039, w_eco158040, w_eco158041, w_eco158042, w_eco158043, w_eco158044, w_eco158045, w_eco158046, w_eco158047, w_eco158048, w_eco158049, w_eco158050, w_eco158051, w_eco158052, w_eco158053, w_eco158054, w_eco158055, w_eco158056, w_eco158057, w_eco158058, w_eco158059, w_eco158060, w_eco158061, w_eco158062, w_eco158063, w_eco158064, w_eco158065, w_eco158066, w_eco158067, w_eco158068, w_eco158069, w_eco158070, w_eco158071, w_eco158072, w_eco158073, w_eco158074, w_eco158075, w_eco158076, w_eco158077, w_eco158078, w_eco158079, w_eco158080, w_eco158081, w_eco158082, w_eco158083, w_eco158084, w_eco158085, w_eco158086, w_eco158087, w_eco158088, w_eco158089, w_eco158090, w_eco158091, w_eco158092, w_eco158093, w_eco158094, w_eco158095, w_eco158096, w_eco158097, w_eco158098, w_eco158099, w_eco158100, w_eco158101, w_eco158102, w_eco158103, w_eco158104, w_eco158105, w_eco158106, w_eco158107, w_eco158108, w_eco158109, w_eco158110, w_eco158111, w_eco158112, w_eco158113, w_eco158114, w_eco158115, w_eco158116, w_eco158117, w_eco158118, w_eco158119, w_eco158120, w_eco158121, w_eco158122, w_eco158123, w_eco158124, w_eco158125, w_eco158126, w_eco158127, w_eco158128, w_eco158129, w_eco158130, w_eco158131, w_eco158132, w_eco158133, w_eco158134, w_eco158135, w_eco158136, w_eco158137, w_eco158138, w_eco158139, w_eco158140, w_eco158141, w_eco158142, w_eco158143, w_eco158144, w_eco158145, w_eco158146, w_eco158147, w_eco158148, w_eco158149, w_eco158150, w_eco158151, w_eco158152, w_eco158153, w_eco158154, w_eco158155, w_eco158156, w_eco158157, w_eco158158, w_eco158159, w_eco158160, w_eco158161, w_eco158162, w_eco158163, w_eco158164, w_eco158165, w_eco158166, w_eco158167, w_eco158168, w_eco158169, w_eco158170, w_eco158171, w_eco158172, w_eco158173, w_eco158174, w_eco158175, w_eco158176, w_eco158177, w_eco158178, w_eco158179, w_eco158180, w_eco158181, w_eco158182, w_eco158183, w_eco158184, w_eco158185, w_eco158186, w_eco158187, w_eco158188, w_eco158189, w_eco158190, w_eco158191, w_eco158192, w_eco158193, w_eco158194, w_eco158195, w_eco158196, w_eco158197, w_eco158198, w_eco158199, w_eco158200, w_eco158201, w_eco158202, w_eco158203, w_eco158204, w_eco158205, w_eco158206, w_eco158207, w_eco158208, w_eco158209, w_eco158210, w_eco158211, w_eco158212, w_eco158213, w_eco158214, w_eco158215, w_eco158216, w_eco158217, w_eco158218, w_eco158219, w_eco158220, w_eco158221, w_eco158222, w_eco158223, w_eco158224, w_eco158225, w_eco158226, w_eco158227, w_eco158228, w_eco158229, w_eco158230, w_eco158231, w_eco158232, w_eco158233, w_eco158234, w_eco158235, w_eco158236, w_eco158237, w_eco158238, w_eco158239, w_eco158240, w_eco158241, w_eco158242, w_eco158243, w_eco158244, w_eco158245, w_eco158246, w_eco158247, w_eco158248, w_eco158249, w_eco158250, w_eco158251, w_eco158252, w_eco158253, w_eco158254, w_eco158255, w_eco158256, w_eco158257, w_eco158258, w_eco158259, w_eco158260, w_eco158261, w_eco158262, w_eco158263, w_eco158264, w_eco158265, w_eco158266, w_eco158267, w_eco158268, w_eco158269, w_eco158270, w_eco158271, w_eco158272, w_eco158273, w_eco158274, w_eco158275, w_eco158276, w_eco158277, w_eco158278, w_eco158279, w_eco158280, w_eco158281, w_eco158282, w_eco158283, w_eco158284, w_eco158285, w_eco158286, w_eco158287, w_eco158288, w_eco158289, w_eco158290, w_eco158291, w_eco158292, w_eco158293, w_eco158294, w_eco158295, w_eco158296, w_eco158297, w_eco158298, w_eco158299, w_eco158300, w_eco158301, w_eco158302, w_eco158303, w_eco158304, w_eco158305, w_eco158306, w_eco158307, w_eco158308, w_eco158309, w_eco158310, w_eco158311, w_eco158312, w_eco158313, w_eco158314, w_eco158315, w_eco158316, w_eco158317, w_eco158318, w_eco158319, w_eco158320, w_eco158321, w_eco158322, w_eco158323, w_eco158324, w_eco158325, w_eco158326, w_eco158327, w_eco158328, w_eco158329, w_eco158330, w_eco158331, w_eco158332, w_eco158333, w_eco158334, w_eco158335, w_eco158336, w_eco158337, w_eco158338, w_eco158339, w_eco158340, w_eco158341, w_eco158342, w_eco158343, w_eco158344, w_eco158345, w_eco158346, w_eco158347, w_eco158348, w_eco158349, w_eco158350, w_eco158351, w_eco158352, w_eco158353, w_eco158354, w_eco158355, w_eco158356, w_eco158357, w_eco158358, w_eco158359, w_eco158360, w_eco158361, w_eco158362, w_eco158363, w_eco158364, w_eco158365, w_eco158366, w_eco158367, w_eco158368, w_eco158369, w_eco158370, w_eco158371, w_eco158372, w_eco158373, w_eco158374, w_eco158375, w_eco158376, w_eco158377, w_eco158378, w_eco158379, w_eco158380, w_eco158381, w_eco158382, w_eco158383, w_eco158384, w_eco158385, w_eco158386, w_eco158387, w_eco158388, w_eco158389, w_eco158390, w_eco158391, w_eco158392, w_eco158393, w_eco158394, w_eco158395, w_eco158396, w_eco158397, w_eco158398, w_eco158399, w_eco158400, w_eco158401, w_eco158402, w_eco158403, w_eco158404, w_eco158405, w_eco158406, w_eco158407, w_eco158408, w_eco158409, w_eco158410, w_eco158411, w_eco158412, w_eco158413, w_eco158414, w_eco158415, w_eco158416, w_eco158417, w_eco158418, w_eco158419, w_eco158420, w_eco158421, w_eco158422, w_eco158423, w_eco158424, w_eco158425, w_eco158426, w_eco158427, w_eco158428, w_eco158429, w_eco158430, w_eco158431, w_eco158432, w_eco158433, w_eco158434, w_eco158435, w_eco158436, w_eco158437, w_eco158438, w_eco158439, w_eco158440, w_eco158441, w_eco158442, w_eco158443, w_eco158444, w_eco158445, w_eco158446, w_eco158447, w_eco158448, w_eco158449, w_eco158450, w_eco158451, w_eco158452, w_eco158453, w_eco158454, w_eco158455, w_eco158456, w_eco158457, w_eco158458, w_eco158459, w_eco158460, w_eco158461, w_eco158462, w_eco158463, w_eco158464, w_eco158465, w_eco158466, w_eco158467, w_eco158468, w_eco158469, w_eco158470, w_eco158471, w_eco158472, w_eco158473, w_eco158474, w_eco158475, w_eco158476, w_eco158477, w_eco158478, w_eco158479, w_eco158480, w_eco158481, w_eco158482, w_eco158483, w_eco158484, w_eco158485, w_eco158486, w_eco158487, w_eco158488, w_eco158489, w_eco158490, w_eco158491, w_eco158492, w_eco158493, w_eco158494, w_eco158495, w_eco158496, w_eco158497, w_eco158498, w_eco158499, w_eco158500, w_eco158501, w_eco158502, w_eco158503, w_eco158504, w_eco158505, w_eco158506, w_eco158507, w_eco158508, w_eco158509, w_eco158510, w_eco158511, w_eco158512, w_eco158513, w_eco158514, w_eco158515, w_eco158516, w_eco158517, w_eco158518, w_eco158519, w_eco158520, w_eco158521, w_eco158522, w_eco158523, w_eco158524, w_eco158525, w_eco158526, w_eco158527, w_eco158528, w_eco158529, w_eco158530, w_eco158531, w_eco158532, w_eco158533, w_eco158534, w_eco158535, w_eco158536, w_eco158537, w_eco158538, w_eco158539, w_eco158540, w_eco158541, w_eco158542, w_eco158543, w_eco158544, w_eco158545, w_eco158546, w_eco158547, w_eco158548, w_eco158549, w_eco158550, w_eco158551, w_eco158552, w_eco158553, w_eco158554, w_eco158555, w_eco158556, w_eco158557, w_eco158558, w_eco158559, w_eco158560, w_eco158561, w_eco158562, w_eco158563, w_eco158564, w_eco158565, w_eco158566, w_eco158567, w_eco158568, w_eco158569, w_eco158570, w_eco158571, w_eco158572, w_eco158573, w_eco158574, w_eco158575, w_eco158576, w_eco158577, w_eco158578, w_eco158579, w_eco158580, w_eco158581, w_eco158582, w_eco158583, w_eco158584, w_eco158585, w_eco158586, w_eco158587, w_eco158588, w_eco158589, w_eco158590, w_eco158591, w_eco158592, w_eco158593, w_eco158594, w_eco158595, w_eco158596, w_eco158597, w_eco158598, w_eco158599, w_eco158600, w_eco158601, w_eco158602, w_eco158603, w_eco158604, w_eco158605, w_eco158606, w_eco158607, w_eco158608, w_eco158609, w_eco158610, w_eco158611, w_eco158612, w_eco158613, w_eco158614, w_eco158615, w_eco158616, w_eco158617, w_eco158618, w_eco158619, w_eco158620, w_eco158621, w_eco158622, w_eco158623, w_eco158624, w_eco158625, w_eco158626, w_eco158627, w_eco158628, w_eco158629, w_eco158630, w_eco158631, w_eco158632, w_eco158633, w_eco158634, w_eco158635, w_eco158636, w_eco158637, w_eco158638, w_eco158639, w_eco158640, w_eco158641, w_eco158642, w_eco158643, w_eco158644, w_eco158645, w_eco158646, w_eco158647, w_eco158648, w_eco158649, w_eco158650, w_eco158651, w_eco158652, w_eco158653, w_eco158654, w_eco158655, w_eco158656, w_eco158657, w_eco158658, w_eco158659, w_eco158660, w_eco158661, w_eco158662, w_eco158663, w_eco158664, w_eco158665, w_eco158666, w_eco158667, w_eco158668, w_eco158669, w_eco158670, w_eco158671, w_eco158672, w_eco158673, w_eco158674, w_eco158675, w_eco158676, w_eco158677, w_eco158678, w_eco158679, w_eco158680, w_eco158681, w_eco158682, w_eco158683, w_eco158684, w_eco158685, w_eco158686, w_eco158687, w_eco158688, w_eco158689, w_eco158690, w_eco158691, w_eco158692, w_eco158693, w_eco158694, w_eco158695, w_eco158696, w_eco158697, w_eco158698, w_eco158699, w_eco158700, w_eco158701, w_eco158702, w_eco158703, w_eco158704, w_eco158705, w_eco158706, w_eco158707, w_eco158708, w_eco158709, w_eco158710, w_eco158711, w_eco158712, w_eco158713, w_eco158714, w_eco158715, w_eco158716, w_eco158717, w_eco158718, w_eco158719, w_eco158720, w_eco158721, w_eco158722, w_eco158723, w_eco158724, w_eco158725, w_eco158726, w_eco158727, w_eco158728, w_eco158729, w_eco158730, w_eco158731, w_eco158732, w_eco158733, w_eco158734, w_eco158735, w_eco158736, w_eco158737, w_eco158738, w_eco158739, w_eco158740, w_eco158741, w_eco158742, w_eco158743, w_eco158744, w_eco158745, w_eco158746, w_eco158747, w_eco158748, w_eco158749, w_eco158750, w_eco158751, w_eco158752, w_eco158753, w_eco158754, w_eco158755, w_eco158756, w_eco158757, w_eco158758, w_eco158759, w_eco158760, w_eco158761, w_eco158762, w_eco158763, w_eco158764, w_eco158765, w_eco158766, w_eco158767, w_eco158768, w_eco158769, w_eco158770, w_eco158771, w_eco158772, w_eco158773, w_eco158774, w_eco158775, w_eco158776, w_eco158777, w_eco158778, w_eco158779, w_eco158780, w_eco158781, w_eco158782, w_eco158783, w_eco158784, w_eco158785, w_eco158786, w_eco158787, w_eco158788, w_eco158789, w_eco158790, w_eco158791, w_eco158792, w_eco158793, w_eco158794, w_eco158795, w_eco158796, w_eco158797, w_eco158798, w_eco158799, w_eco158800, w_eco158801, w_eco158802, w_eco158803, w_eco158804, w_eco158805, w_eco158806, w_eco158807, w_eco158808, w_eco158809, w_eco158810, w_eco158811, w_eco158812, w_eco158813, w_eco158814, w_eco158815, w_eco158816, w_eco158817, w_eco158818, w_eco158819, w_eco158820, w_eco158821, w_eco158822, w_eco158823, w_eco158824, w_eco158825, w_eco158826, w_eco158827, w_eco158828, w_eco158829, w_eco158830, w_eco158831, w_eco158832, w_eco158833, w_eco158834, w_eco158835, w_eco158836, w_eco158837, w_eco158838, w_eco158839, w_eco158840, w_eco158841, w_eco158842, w_eco158843, w_eco158844, w_eco158845, w_eco158846, w_eco158847, w_eco158848, w_eco158849, w_eco158850, w_eco158851, w_eco158852, w_eco158853, w_eco158854, w_eco158855, w_eco158856, w_eco158857, w_eco158858, w_eco158859, w_eco158860, w_eco158861, w_eco158862, w_eco158863, w_eco158864, w_eco158865, w_eco158866, w_eco158867, w_eco158868, w_eco158869, w_eco158870, w_eco158871, w_eco158872, w_eco158873, w_eco158874, w_eco158875, w_eco158876, w_eco158877, w_eco158878, w_eco158879, w_eco158880, w_eco158881, w_eco158882, w_eco158883, w_eco158884, w_eco158885, w_eco158886, w_eco158887, w_eco158888, w_eco158889, w_eco158890, w_eco158891, w_eco158892, w_eco158893, w_eco158894, w_eco158895, w_eco158896, w_eco158897, w_eco158898, w_eco158899, w_eco158900, w_eco158901, w_eco158902, w_eco158903, w_eco158904, w_eco158905, w_eco158906, w_eco158907, w_eco158908, w_eco158909, w_eco158910, w_eco158911, w_eco158912, w_eco158913, w_eco158914, w_eco158915, w_eco158916, w_eco158917, w_eco158918, w_eco158919, w_eco158920, w_eco158921, w_eco158922, w_eco158923, w_eco158924, w_eco158925, w_eco158926, w_eco158927, w_eco158928, w_eco158929, w_eco158930, w_eco158931, w_eco158932, w_eco158933, w_eco158934, w_eco158935, w_eco158936, w_eco158937, w_eco158938, w_eco158939, w_eco158940, w_eco158941, w_eco158942, w_eco158943, w_eco158944, w_eco158945, w_eco158946, w_eco158947, w_eco158948, w_eco158949, w_eco158950, w_eco158951, w_eco158952, w_eco158953, w_eco158954, w_eco158955, w_eco158956, w_eco158957, w_eco158958, w_eco158959, w_eco158960, w_eco158961, w_eco158962, w_eco158963, w_eco158964, w_eco158965, w_eco158966, w_eco158967, w_eco158968, w_eco158969, w_eco158970, w_eco158971, w_eco158972, w_eco158973, w_eco158974, w_eco158975, w_eco158976, w_eco158977, w_eco158978, w_eco158979, w_eco158980, w_eco158981, w_eco158982, w_eco158983, w_eco158984, w_eco158985, w_eco158986, w_eco158987, w_eco158988, w_eco158989, w_eco158990, w_eco158991, w_eco158992, w_eco158993, w_eco158994, w_eco158995, w_eco158996, w_eco158997, w_eco158998, w_eco158999, w_eco159000, w_eco159001, w_eco159002, w_eco159003, w_eco159004, w_eco159005, w_eco159006, w_eco159007, w_eco159008, w_eco159009, w_eco159010, w_eco159011, w_eco159012, w_eco159013, w_eco159014, w_eco159015, w_eco159016, w_eco159017, w_eco159018, w_eco159019, w_eco159020, w_eco159021, w_eco159022, w_eco159023, w_eco159024, w_eco159025, w_eco159026, w_eco159027, w_eco159028, w_eco159029, w_eco159030, w_eco159031, w_eco159032, w_eco159033, w_eco159034, w_eco159035, w_eco159036, w_eco159037, w_eco159038, w_eco159039, w_eco159040, w_eco159041, w_eco159042, w_eco159043, w_eco159044, w_eco159045, w_eco159046, w_eco159047, w_eco159048, w_eco159049, w_eco159050, w_eco159051, w_eco159052, w_eco159053, w_eco159054, w_eco159055, w_eco159056, w_eco159057, w_eco159058, w_eco159059, w_eco159060, w_eco159061, w_eco159062, w_eco159063, w_eco159064, w_eco159065, w_eco159066, w_eco159067, w_eco159068, w_eco159069, w_eco159070, w_eco159071, w_eco159072, w_eco159073, w_eco159074, w_eco159075, w_eco159076, w_eco159077, w_eco159078, w_eco159079, w_eco159080, w_eco159081, w_eco159082, w_eco159083, w_eco159084, w_eco159085, w_eco159086, w_eco159087, w_eco159088, w_eco159089, w_eco159090, w_eco159091, w_eco159092, w_eco159093, w_eco159094, w_eco159095, w_eco159096, w_eco159097, w_eco159098, w_eco159099, w_eco159100, w_eco159101, w_eco159102, w_eco159103, w_eco159104, w_eco159105, w_eco159106, w_eco159107, w_eco159108, w_eco159109, w_eco159110, w_eco159111, w_eco159112, w_eco159113, w_eco159114, w_eco159115, w_eco159116, w_eco159117, w_eco159118, w_eco159119, w_eco159120, w_eco159121, w_eco159122, w_eco159123, w_eco159124, w_eco159125, w_eco159126, w_eco159127, w_eco159128, w_eco159129, w_eco159130, w_eco159131, w_eco159132, w_eco159133, w_eco159134, w_eco159135, w_eco159136, w_eco159137, w_eco159138, w_eco159139, w_eco159140, w_eco159141, w_eco159142, w_eco159143, w_eco159144, w_eco159145, w_eco159146, w_eco159147, w_eco159148, w_eco159149, w_eco159150, w_eco159151, w_eco159152, w_eco159153, w_eco159154, w_eco159155, w_eco159156, w_eco159157, w_eco159158, w_eco159159, w_eco159160, w_eco159161, w_eco159162, w_eco159163, w_eco159164, w_eco159165, w_eco159166, w_eco159167, w_eco159168, w_eco159169, w_eco159170, w_eco159171, w_eco159172, w_eco159173, w_eco159174, w_eco159175, w_eco159176, w_eco159177, w_eco159178, w_eco159179, w_eco159180, w_eco159181, w_eco159182, w_eco159183, w_eco159184, w_eco159185, w_eco159186, w_eco159187, w_eco159188, w_eco159189, w_eco159190, w_eco159191, w_eco159192, w_eco159193, w_eco159194, w_eco159195, w_eco159196, w_eco159197, w_eco159198, w_eco159199, w_eco159200, w_eco159201, w_eco159202, w_eco159203, w_eco159204, w_eco159205, w_eco159206, w_eco159207, w_eco159208, w_eco159209, w_eco159210, w_eco159211, w_eco159212, w_eco159213, w_eco159214, w_eco159215, w_eco159216, w_eco159217, w_eco159218, w_eco159219, w_eco159220, w_eco159221, w_eco159222, w_eco159223, w_eco159224, w_eco159225, w_eco159226, w_eco159227, w_eco159228, w_eco159229, w_eco159230, w_eco159231, w_eco159232, w_eco159233, w_eco159234, w_eco159235, w_eco159236, w_eco159237, w_eco159238, w_eco159239, w_eco159240, w_eco159241, w_eco159242, w_eco159243, w_eco159244, w_eco159245, w_eco159246, w_eco159247, w_eco159248, w_eco159249, w_eco159250, w_eco159251, w_eco159252, w_eco159253, w_eco159254, w_eco159255, w_eco159256, w_eco159257, w_eco159258, w_eco159259, w_eco159260, w_eco159261, w_eco159262, w_eco159263, w_eco159264, w_eco159265, w_eco159266, w_eco159267, w_eco159268, w_eco159269, w_eco159270, w_eco159271, w_eco159272, w_eco159273, w_eco159274, w_eco159275, w_eco159276, w_eco159277, w_eco159278, w_eco159279, w_eco159280, w_eco159281, w_eco159282, w_eco159283, w_eco159284, w_eco159285, w_eco159286, w_eco159287, w_eco159288, w_eco159289, w_eco159290, w_eco159291, w_eco159292, w_eco159293, w_eco159294, w_eco159295, w_eco159296, w_eco159297, w_eco159298, w_eco159299, w_eco159300, w_eco159301, w_eco159302, w_eco159303, w_eco159304, w_eco159305, w_eco159306, w_eco159307, w_eco159308, w_eco159309, w_eco159310, w_eco159311, w_eco159312, w_eco159313, w_eco159314, w_eco159315, w_eco159316, w_eco159317, w_eco159318, w_eco159319, w_eco159320, w_eco159321, w_eco159322, w_eco159323, w_eco159324, w_eco159325, w_eco159326, w_eco159327, w_eco159328, w_eco159329, w_eco159330, w_eco159331, w_eco159332, w_eco159333, w_eco159334, w_eco159335, w_eco159336, w_eco159337, w_eco159338, w_eco159339, w_eco159340, w_eco159341, w_eco159342, w_eco159343, w_eco159344, w_eco159345, w_eco159346, w_eco159347, w_eco159348, w_eco159349, w_eco159350, w_eco159351, w_eco159352, w_eco159353, w_eco159354, w_eco159355, w_eco159356, w_eco159357, w_eco159358, w_eco159359, w_eco159360, w_eco159361, w_eco159362, w_eco159363, w_eco159364, w_eco159365, w_eco159366, w_eco159367, w_eco159368, w_eco159369, w_eco159370, w_eco159371, w_eco159372, w_eco159373, w_eco159374, w_eco159375, w_eco159376, w_eco159377, w_eco159378, w_eco159379, w_eco159380, w_eco159381, w_eco159382, w_eco159383, w_eco159384, w_eco159385, w_eco159386, w_eco159387, w_eco159388, w_eco159389, w_eco159390, w_eco159391, w_eco159392, w_eco159393, w_eco159394, w_eco159395, w_eco159396, w_eco159397, w_eco159398, w_eco159399, w_eco159400, w_eco159401, w_eco159402, w_eco159403, w_eco159404, w_eco159405, w_eco159406, w_eco159407, w_eco159408, w_eco159409, w_eco159410, w_eco159411, w_eco159412, w_eco159413, w_eco159414, w_eco159415, w_eco159416, w_eco159417, w_eco159418, w_eco159419, w_eco159420, w_eco159421, w_eco159422, w_eco159423, w_eco159424, w_eco159425, w_eco159426, w_eco159427, w_eco159428, w_eco159429, w_eco159430, w_eco159431, w_eco159432, w_eco159433, w_eco159434, w_eco159435, w_eco159436, w_eco159437, w_eco159438, w_eco159439, w_eco159440, w_eco159441, w_eco159442, w_eco159443, w_eco159444, w_eco159445, w_eco159446, w_eco159447, w_eco159448, w_eco159449, w_eco159450, w_eco159451, w_eco159452, w_eco159453, w_eco159454, w_eco159455, w_eco159456, w_eco159457, w_eco159458, w_eco159459, w_eco159460, w_eco159461, w_eco159462, w_eco159463, w_eco159464, w_eco159465, w_eco159466, w_eco159467, w_eco159468, w_eco159469, w_eco159470, w_eco159471, w_eco159472, w_eco159473, w_eco159474, w_eco159475, w_eco159476, w_eco159477, w_eco159478, w_eco159479, w_eco159480, w_eco159481, w_eco159482, w_eco159483, w_eco159484, w_eco159485, w_eco159486, w_eco159487, w_eco159488, w_eco159489, w_eco159490, w_eco159491, w_eco159492, w_eco159493, w_eco159494, w_eco159495, w_eco159496, w_eco159497, w_eco159498, w_eco159499, w_eco159500, w_eco159501, w_eco159502, w_eco159503, w_eco159504, w_eco159505, w_eco159506, w_eco159507, w_eco159508, w_eco159509, w_eco159510, w_eco159511, w_eco159512, w_eco159513, w_eco159514, w_eco159515, w_eco159516, w_eco159517, w_eco159518, w_eco159519, w_eco159520, w_eco159521, w_eco159522, w_eco159523, w_eco159524, w_eco159525, w_eco159526, w_eco159527, w_eco159528, w_eco159529, w_eco159530, w_eco159531, w_eco159532, w_eco159533, w_eco159534, w_eco159535, w_eco159536, w_eco159537, w_eco159538, w_eco159539, w_eco159540, w_eco159541, w_eco159542, w_eco159543, w_eco159544, w_eco159545, w_eco159546, w_eco159547, w_eco159548, w_eco159549, w_eco159550, w_eco159551, w_eco159552, w_eco159553, w_eco159554, w_eco159555, w_eco159556, w_eco159557, w_eco159558, w_eco159559, w_eco159560, w_eco159561, w_eco159562, w_eco159563, w_eco159564, w_eco159565, w_eco159566, w_eco159567, w_eco159568, w_eco159569, w_eco159570, w_eco159571, w_eco159572, w_eco159573, w_eco159574, w_eco159575, w_eco159576, w_eco159577, w_eco159578, w_eco159579, w_eco159580, w_eco159581, w_eco159582, w_eco159583, w_eco159584, w_eco159585, w_eco159586, w_eco159587, w_eco159588, w_eco159589, w_eco159590, w_eco159591, w_eco159592, w_eco159593, w_eco159594, w_eco159595, w_eco159596, w_eco159597, w_eco159598, w_eco159599, w_eco159600, w_eco159601, w_eco159602, w_eco159603, w_eco159604, w_eco159605, w_eco159606, w_eco159607, w_eco159608, w_eco159609, w_eco159610, w_eco159611, w_eco159612, w_eco159613, w_eco159614, w_eco159615, w_eco159616, w_eco159617, w_eco159618, w_eco159619, w_eco159620, w_eco159621, w_eco159622, w_eco159623, w_eco159624, w_eco159625, w_eco159626, w_eco159627, w_eco159628, w_eco159629, w_eco159630, w_eco159631, w_eco159632, w_eco159633, w_eco159634, w_eco159635, w_eco159636, w_eco159637, w_eco159638, w_eco159639, w_eco159640, w_eco159641, w_eco159642, w_eco159643, w_eco159644, w_eco159645, w_eco159646, w_eco159647, w_eco159648, w_eco159649, w_eco159650, w_eco159651, w_eco159652, w_eco159653, w_eco159654, w_eco159655, w_eco159656, w_eco159657, w_eco159658, w_eco159659, w_eco159660, w_eco159661, w_eco159662, w_eco159663, w_eco159664, w_eco159665, w_eco159666, w_eco159667, w_eco159668, w_eco159669, w_eco159670, w_eco159671, w_eco159672, w_eco159673, w_eco159674, w_eco159675, w_eco159676, w_eco159677, w_eco159678, w_eco159679, w_eco159680, w_eco159681, w_eco159682, w_eco159683, w_eco159684, w_eco159685, w_eco159686, w_eco159687, w_eco159688, w_eco159689, w_eco159690, w_eco159691, w_eco159692, w_eco159693, w_eco159694, w_eco159695, w_eco159696, w_eco159697, w_eco159698, w_eco159699, w_eco159700, w_eco159701, w_eco159702, w_eco159703, w_eco159704, w_eco159705, w_eco159706, w_eco159707, w_eco159708, w_eco159709, w_eco159710, w_eco159711, w_eco159712, w_eco159713, w_eco159714, w_eco159715, w_eco159716, w_eco159717, w_eco159718, w_eco159719, w_eco159720, w_eco159721, w_eco159722, w_eco159723, w_eco159724, w_eco159725, w_eco159726, w_eco159727, w_eco159728, w_eco159729, w_eco159730, w_eco159731, w_eco159732, w_eco159733, w_eco159734, w_eco159735, w_eco159736, w_eco159737, w_eco159738, w_eco159739, w_eco159740, w_eco159741, w_eco159742, w_eco159743, w_eco159744, w_eco159745, w_eco159746, w_eco159747, w_eco159748, w_eco159749, w_eco159750, w_eco159751, w_eco159752, w_eco159753, w_eco159754, w_eco159755, w_eco159756, w_eco159757, w_eco159758, w_eco159759, w_eco159760, w_eco159761, w_eco159762, w_eco159763, w_eco159764, w_eco159765, w_eco159766, w_eco159767, w_eco159768, w_eco159769, w_eco159770, w_eco159771, w_eco159772, w_eco159773, w_eco159774, w_eco159775, w_eco159776, w_eco159777, w_eco159778, w_eco159779, w_eco159780, w_eco159781, w_eco159782, w_eco159783, w_eco159784, w_eco159785, w_eco159786, w_eco159787, w_eco159788, w_eco159789, w_eco159790, w_eco159791, w_eco159792, w_eco159793, w_eco159794, w_eco159795, w_eco159796, w_eco159797, w_eco159798, w_eco159799, w_eco159800, w_eco159801, w_eco159802, w_eco159803, w_eco159804, w_eco159805, w_eco159806, w_eco159807, w_eco159808, w_eco159809, w_eco159810, w_eco159811, w_eco159812, w_eco159813, w_eco159814, w_eco159815, w_eco159816, w_eco159817, w_eco159818, w_eco159819, w_eco159820, w_eco159821, w_eco159822, w_eco159823, w_eco159824, w_eco159825, w_eco159826, w_eco159827, w_eco159828, w_eco159829, w_eco159830, w_eco159831, w_eco159832, w_eco159833, w_eco159834, w_eco159835, w_eco159836, w_eco159837, w_eco159838, w_eco159839, w_eco159840, w_eco159841, w_eco159842, w_eco159843, w_eco159844, w_eco159845, w_eco159846, w_eco159847, w_eco159848, w_eco159849, w_eco159850, w_eco159851, w_eco159852, w_eco159853, w_eco159854, w_eco159855, w_eco159856, w_eco159857, w_eco159858, w_eco159859, w_eco159860, w_eco159861, w_eco159862, w_eco159863, w_eco159864, w_eco159865, w_eco159866, w_eco159867, w_eco159868, w_eco159869, w_eco159870, w_eco159871, w_eco159872, w_eco159873, w_eco159874, w_eco159875, w_eco159876, w_eco159877, w_eco159878, w_eco159879, w_eco159880, w_eco159881, w_eco159882, w_eco159883, w_eco159884, w_eco159885, w_eco159886, w_eco159887, w_eco159888, w_eco159889, w_eco159890, w_eco159891, w_eco159892, w_eco159893, w_eco159894, w_eco159895, w_eco159896, w_eco159897, w_eco159898, w_eco159899, w_eco159900, w_eco159901, w_eco159902, w_eco159903, w_eco159904, w_eco159905, w_eco159906, w_eco159907, w_eco159908, w_eco159909, w_eco159910, w_eco159911, w_eco159912, w_eco159913, w_eco159914, w_eco159915, w_eco159916, w_eco159917, w_eco159918, w_eco159919, w_eco159920, w_eco159921, w_eco159922, w_eco159923, w_eco159924, w_eco159925, w_eco159926, w_eco159927, w_eco159928, w_eco159929, w_eco159930, w_eco159931, w_eco159932, w_eco159933, w_eco159934, w_eco159935, w_eco159936, w_eco159937, w_eco159938, w_eco159939, w_eco159940, w_eco159941, w_eco159942, w_eco159943, w_eco159944, w_eco159945, w_eco159946, w_eco159947, w_eco159948, w_eco159949, w_eco159950, w_eco159951, w_eco159952, w_eco159953, w_eco159954, w_eco159955, w_eco159956, w_eco159957, w_eco159958, w_eco159959, w_eco159960, w_eco159961, w_eco159962, w_eco159963, w_eco159964, w_eco159965, w_eco159966, w_eco159967, w_eco159968, w_eco159969, w_eco159970, w_eco159971, w_eco159972, w_eco159973, w_eco159974, w_eco159975, w_eco159976, w_eco159977, w_eco159978, w_eco159979, w_eco159980, w_eco159981, w_eco159982, w_eco159983, w_eco159984, w_eco159985, w_eco159986, w_eco159987, w_eco159988, w_eco159989, w_eco159990, w_eco159991, w_eco159992, w_eco159993, w_eco159994, w_eco159995, w_eco159996, w_eco159997, w_eco159998, w_eco159999, w_eco160000, w_eco160001, w_eco160002, w_eco160003, w_eco160004, w_eco160005, w_eco160006, w_eco160007, w_eco160008, w_eco160009, w_eco160010, w_eco160011, w_eco160012, w_eco160013, w_eco160014, w_eco160015, w_eco160016, w_eco160017, w_eco160018, w_eco160019, w_eco160020, w_eco160021, w_eco160022, w_eco160023, w_eco160024, w_eco160025, w_eco160026, w_eco160027, w_eco160028, w_eco160029, w_eco160030, w_eco160031, w_eco160032, w_eco160033, w_eco160034, w_eco160035, w_eco160036, w_eco160037, w_eco160038, w_eco160039, w_eco160040, w_eco160041, w_eco160042, w_eco160043, w_eco160044, w_eco160045, w_eco160046, w_eco160047, w_eco160048, w_eco160049, w_eco160050, w_eco160051, w_eco160052, w_eco160053, w_eco160054, w_eco160055, w_eco160056, w_eco160057, w_eco160058, w_eco160059, w_eco160060, w_eco160061, w_eco160062, w_eco160063, w_eco160064, w_eco160065, w_eco160066, w_eco160067, w_eco160068, w_eco160069, w_eco160070, w_eco160071, w_eco160072, w_eco160073, w_eco160074, w_eco160075, w_eco160076, w_eco160077, w_eco160078, w_eco160079, w_eco160080, w_eco160081, w_eco160082, w_eco160083, w_eco160084, w_eco160085, w_eco160086, w_eco160087, w_eco160088, w_eco160089, w_eco160090, w_eco160091, w_eco160092, w_eco160093, w_eco160094, w_eco160095, w_eco160096, w_eco160097, w_eco160098, w_eco160099, w_eco160100, w_eco160101, w_eco160102, w_eco160103, w_eco160104, w_eco160105, w_eco160106, w_eco160107, w_eco160108, w_eco160109, w_eco160110, w_eco160111, w_eco160112, w_eco160113, w_eco160114, w_eco160115, w_eco160116, w_eco160117, w_eco160118, w_eco160119, w_eco160120, w_eco160121, w_eco160122, w_eco160123, w_eco160124, w_eco160125, w_eco160126, w_eco160127, w_eco160128, w_eco160129, w_eco160130, w_eco160131, w_eco160132, w_eco160133, w_eco160134, w_eco160135, w_eco160136, w_eco160137, w_eco160138, w_eco160139, w_eco160140, w_eco160141, w_eco160142, w_eco160143, w_eco160144, w_eco160145, w_eco160146, w_eco160147, w_eco160148, w_eco160149, w_eco160150, w_eco160151, w_eco160152, w_eco160153, w_eco160154, w_eco160155, w_eco160156, w_eco160157, w_eco160158, w_eco160159, w_eco160160, w_eco160161, w_eco160162, w_eco160163, w_eco160164, w_eco160165, w_eco160166, w_eco160167, w_eco160168, w_eco160169, w_eco160170, w_eco160171, w_eco160172, w_eco160173, w_eco160174, w_eco160175, w_eco160176, w_eco160177, w_eco160178, w_eco160179, w_eco160180, w_eco160181, w_eco160182, w_eco160183, w_eco160184, w_eco160185, w_eco160186, w_eco160187, w_eco160188, w_eco160189, w_eco160190, w_eco160191, w_eco160192, w_eco160193, w_eco160194, w_eco160195, w_eco160196, w_eco160197, w_eco160198, w_eco160199, w_eco160200, w_eco160201, w_eco160202, w_eco160203, w_eco160204, w_eco160205, w_eco160206, w_eco160207, w_eco160208, w_eco160209, w_eco160210, w_eco160211, w_eco160212, w_eco160213, w_eco160214, w_eco160215, w_eco160216, w_eco160217, w_eco160218, w_eco160219, w_eco160220, w_eco160221, w_eco160222, w_eco160223, w_eco160224, w_eco160225, w_eco160226, w_eco160227, w_eco160228, w_eco160229, w_eco160230, w_eco160231, w_eco160232, w_eco160233, w_eco160234, w_eco160235, w_eco160236, w_eco160237, w_eco160238, w_eco160239, w_eco160240, w_eco160241, w_eco160242, w_eco160243, w_eco160244, w_eco160245, w_eco160246, w_eco160247, w_eco160248, w_eco160249, w_eco160250, w_eco160251, w_eco160252, w_eco160253, w_eco160254, w_eco160255, w_eco160256, w_eco160257, w_eco160258, w_eco160259, w_eco160260, w_eco160261, w_eco160262, w_eco160263, w_eco160264, w_eco160265, w_eco160266, w_eco160267, w_eco160268, w_eco160269, w_eco160270, w_eco160271, w_eco160272, w_eco160273, w_eco160274, w_eco160275, w_eco160276, w_eco160277, w_eco160278, w_eco160279, w_eco160280, w_eco160281, w_eco160282, w_eco160283, w_eco160284, w_eco160285, w_eco160286, w_eco160287, w_eco160288, w_eco160289, w_eco160290, w_eco160291, w_eco160292, w_eco160293, w_eco160294, w_eco160295, w_eco160296, w_eco160297, w_eco160298, w_eco160299, w_eco160300, w_eco160301, w_eco160302, w_eco160303, w_eco160304, w_eco160305, w_eco160306, w_eco160307, w_eco160308, w_eco160309, w_eco160310, w_eco160311, w_eco160312, w_eco160313, w_eco160314, w_eco160315, w_eco160316, w_eco160317, w_eco160318, w_eco160319, w_eco160320, w_eco160321, w_eco160322, w_eco160323, w_eco160324, w_eco160325, w_eco160326, w_eco160327, w_eco160328, w_eco160329, w_eco160330, w_eco160331, w_eco160332, w_eco160333, w_eco160334, w_eco160335, w_eco160336, w_eco160337, w_eco160338, w_eco160339, w_eco160340, w_eco160341, w_eco160342, w_eco160343, w_eco160344, w_eco160345, w_eco160346, w_eco160347, w_eco160348, w_eco160349, w_eco160350, w_eco160351, w_eco160352, w_eco160353, w_eco160354, w_eco160355, w_eco160356, w_eco160357, w_eco160358, w_eco160359, w_eco160360, w_eco160361, w_eco160362, w_eco160363, w_eco160364, w_eco160365, w_eco160366, w_eco160367, w_eco160368, w_eco160369, w_eco160370, w_eco160371, w_eco160372, w_eco160373, w_eco160374, w_eco160375, w_eco160376, w_eco160377, w_eco160378, w_eco160379, w_eco160380, w_eco160381, w_eco160382, w_eco160383, w_eco160384, w_eco160385, w_eco160386, w_eco160387, w_eco160388, w_eco160389, w_eco160390, w_eco160391, w_eco160392, w_eco160393, w_eco160394, w_eco160395, w_eco160396, w_eco160397, w_eco160398, w_eco160399, w_eco160400, w_eco160401, w_eco160402, w_eco160403, w_eco160404, w_eco160405, w_eco160406, w_eco160407, w_eco160408, w_eco160409, w_eco160410, w_eco160411, w_eco160412, w_eco160413, w_eco160414, w_eco160415, w_eco160416, w_eco160417, w_eco160418, w_eco160419, w_eco160420, w_eco160421, w_eco160422, w_eco160423, w_eco160424, w_eco160425, w_eco160426, w_eco160427, w_eco160428, w_eco160429, w_eco160430, w_eco160431, w_eco160432, w_eco160433, w_eco160434, w_eco160435, w_eco160436, w_eco160437, w_eco160438, w_eco160439, w_eco160440, w_eco160441, w_eco160442, w_eco160443, w_eco160444, w_eco160445, w_eco160446, w_eco160447, w_eco160448, w_eco160449, w_eco160450, w_eco160451, w_eco160452, w_eco160453, w_eco160454, w_eco160455, w_eco160456, w_eco160457, w_eco160458, w_eco160459, w_eco160460, w_eco160461, w_eco160462, w_eco160463, w_eco160464, w_eco160465, w_eco160466, w_eco160467, w_eco160468, w_eco160469, w_eco160470, w_eco160471, w_eco160472, w_eco160473, w_eco160474, w_eco160475, w_eco160476, w_eco160477, w_eco160478, w_eco160479, w_eco160480, w_eco160481, w_eco160482, w_eco160483, w_eco160484, w_eco160485, w_eco160486, w_eco160487, w_eco160488, w_eco160489, w_eco160490, w_eco160491, w_eco160492, w_eco160493, w_eco160494, w_eco160495, w_eco160496, w_eco160497, w_eco160498, w_eco160499, w_eco160500, w_eco160501, w_eco160502, w_eco160503, w_eco160504, w_eco160505, w_eco160506, w_eco160507, w_eco160508, w_eco160509, w_eco160510, w_eco160511, w_eco160512, w_eco160513, w_eco160514, w_eco160515, w_eco160516, w_eco160517, w_eco160518, w_eco160519, w_eco160520, w_eco160521, w_eco160522, w_eco160523, w_eco160524, w_eco160525, w_eco160526, w_eco160527, w_eco160528, w_eco160529, w_eco160530, w_eco160531, w_eco160532, w_eco160533, w_eco160534, w_eco160535, w_eco160536, w_eco160537, w_eco160538, w_eco160539, w_eco160540, w_eco160541, w_eco160542, w_eco160543, w_eco160544, w_eco160545, w_eco160546, w_eco160547, w_eco160548, w_eco160549, w_eco160550, w_eco160551, w_eco160552, w_eco160553, w_eco160554, w_eco160555, w_eco160556, w_eco160557, w_eco160558, w_eco160559, w_eco160560, w_eco160561, w_eco160562, w_eco160563, w_eco160564, w_eco160565, w_eco160566, w_eco160567, w_eco160568, w_eco160569, w_eco160570, w_eco160571, w_eco160572, w_eco160573, w_eco160574, w_eco160575, w_eco160576, w_eco160577, w_eco160578, w_eco160579, w_eco160580, w_eco160581, w_eco160582, w_eco160583, w_eco160584, w_eco160585, w_eco160586, w_eco160587, w_eco160588, w_eco160589, w_eco160590, w_eco160591, w_eco160592, w_eco160593, w_eco160594, w_eco160595, w_eco160596, w_eco160597, w_eco160598, w_eco160599, w_eco160600, w_eco160601, w_eco160602, w_eco160603, w_eco160604, w_eco160605, w_eco160606, w_eco160607, w_eco160608, w_eco160609, w_eco160610, w_eco160611, w_eco160612, w_eco160613, w_eco160614, w_eco160615, w_eco160616, w_eco160617, w_eco160618, w_eco160619, w_eco160620, w_eco160621, w_eco160622, w_eco160623, w_eco160624, w_eco160625, w_eco160626, w_eco160627, w_eco160628, w_eco160629, w_eco160630, w_eco160631, w_eco160632, w_eco160633, w_eco160634, w_eco160635, w_eco160636, w_eco160637, w_eco160638, w_eco160639, w_eco160640, w_eco160641, w_eco160642, w_eco160643, w_eco160644, w_eco160645, w_eco160646, w_eco160647, w_eco160648, w_eco160649, w_eco160650, w_eco160651, w_eco160652, w_eco160653, w_eco160654, w_eco160655, w_eco160656, w_eco160657, w_eco160658, w_eco160659, w_eco160660, w_eco160661, w_eco160662, w_eco160663, w_eco160664, w_eco160665, w_eco160666, w_eco160667, w_eco160668, w_eco160669, w_eco160670, w_eco160671, w_eco160672, w_eco160673, w_eco160674, w_eco160675, w_eco160676, w_eco160677, w_eco160678, w_eco160679, w_eco160680, w_eco160681, w_eco160682, w_eco160683, w_eco160684, w_eco160685, w_eco160686, w_eco160687, w_eco160688, w_eco160689, w_eco160690, w_eco160691, w_eco160692, w_eco160693, w_eco160694, w_eco160695, w_eco160696, w_eco160697, w_eco160698, w_eco160699, w_eco160700, w_eco160701, w_eco160702, w_eco160703, w_eco160704, w_eco160705, w_eco160706, w_eco160707, w_eco160708, w_eco160709, w_eco160710, w_eco160711, w_eco160712, w_eco160713, w_eco160714, w_eco160715, w_eco160716, w_eco160717, w_eco160718, w_eco160719, w_eco160720, w_eco160721, w_eco160722, w_eco160723, w_eco160724, w_eco160725, w_eco160726, w_eco160727, w_eco160728, w_eco160729, w_eco160730, w_eco160731, w_eco160732, w_eco160733, w_eco160734, w_eco160735, w_eco160736, w_eco160737, w_eco160738, w_eco160739, w_eco160740, w_eco160741, w_eco160742, w_eco160743, w_eco160744, w_eco160745, w_eco160746, w_eco160747, w_eco160748, w_eco160749, w_eco160750, w_eco160751, w_eco160752, w_eco160753, w_eco160754, w_eco160755, w_eco160756, w_eco160757, w_eco160758, w_eco160759, w_eco160760, w_eco160761, w_eco160762, w_eco160763, w_eco160764, w_eco160765, w_eco160766, w_eco160767, w_eco160768, w_eco160769, w_eco160770, w_eco160771, w_eco160772, w_eco160773, w_eco160774, w_eco160775, w_eco160776, w_eco160777, w_eco160778, w_eco160779, w_eco160780, w_eco160781, w_eco160782, w_eco160783, w_eco160784, w_eco160785, w_eco160786, w_eco160787, w_eco160788, w_eco160789, w_eco160790, w_eco160791, w_eco160792, w_eco160793, w_eco160794, w_eco160795, w_eco160796, w_eco160797, w_eco160798, w_eco160799, w_eco160800, w_eco160801, w_eco160802, w_eco160803, w_eco160804, w_eco160805, w_eco160806, w_eco160807, w_eco160808, w_eco160809, w_eco160810, w_eco160811, w_eco160812, w_eco160813, w_eco160814, w_eco160815, w_eco160816, w_eco160817, w_eco160818, w_eco160819, w_eco160820, w_eco160821, w_eco160822, w_eco160823, w_eco160824, w_eco160825, w_eco160826, w_eco160827, w_eco160828, w_eco160829, w_eco160830, w_eco160831, w_eco160832, w_eco160833, w_eco160834, w_eco160835, w_eco160836, w_eco160837, w_eco160838, w_eco160839, w_eco160840, w_eco160841, w_eco160842, w_eco160843, w_eco160844, w_eco160845, w_eco160846, w_eco160847, w_eco160848, w_eco160849, w_eco160850, w_eco160851, w_eco160852, w_eco160853, w_eco160854, w_eco160855, w_eco160856, w_eco160857, w_eco160858, w_eco160859, w_eco160860, w_eco160861, w_eco160862, w_eco160863, w_eco160864, w_eco160865, w_eco160866, w_eco160867, w_eco160868, w_eco160869, w_eco160870, w_eco160871, w_eco160872, w_eco160873, w_eco160874, w_eco160875, w_eco160876, w_eco160877, w_eco160878, w_eco160879, w_eco160880, w_eco160881, w_eco160882, w_eco160883, w_eco160884, w_eco160885, w_eco160886, w_eco160887, w_eco160888, w_eco160889, w_eco160890, w_eco160891, w_eco160892, w_eco160893, w_eco160894, w_eco160895, w_eco160896, w_eco160897, w_eco160898, w_eco160899, w_eco160900, w_eco160901, w_eco160902, w_eco160903, w_eco160904, w_eco160905, w_eco160906, w_eco160907, w_eco160908, w_eco160909, w_eco160910, w_eco160911, w_eco160912, w_eco160913, w_eco160914, w_eco160915, w_eco160916, w_eco160917, w_eco160918, w_eco160919, w_eco160920, w_eco160921, w_eco160922, w_eco160923, w_eco160924, w_eco160925, w_eco160926, w_eco160927, w_eco160928, w_eco160929, w_eco160930, w_eco160931, w_eco160932, w_eco160933, w_eco160934, w_eco160935, w_eco160936, w_eco160937, w_eco160938, w_eco160939, w_eco160940, w_eco160941, w_eco160942, w_eco160943, w_eco160944, w_eco160945, w_eco160946, w_eco160947, w_eco160948, w_eco160949, w_eco160950, w_eco160951, w_eco160952, w_eco160953, w_eco160954, w_eco160955, w_eco160956, w_eco160957, w_eco160958, w_eco160959, w_eco160960, w_eco160961, w_eco160962, w_eco160963, w_eco160964, w_eco160965, w_eco160966, w_eco160967, w_eco160968, w_eco160969, w_eco160970, w_eco160971, w_eco160972, w_eco160973, w_eco160974, w_eco160975, w_eco160976, w_eco160977, w_eco160978, w_eco160979, w_eco160980, w_eco160981, w_eco160982, w_eco160983, w_eco160984, w_eco160985, w_eco160986, w_eco160987, w_eco160988, w_eco160989, w_eco160990, w_eco160991, w_eco160992, w_eco160993, w_eco160994, w_eco160995, w_eco160996, w_eco160997, w_eco160998, w_eco160999, w_eco161000, w_eco161001, w_eco161002, w_eco161003, w_eco161004, w_eco161005, w_eco161006, w_eco161007, w_eco161008, w_eco161009, w_eco161010, w_eco161011, w_eco161012, w_eco161013, w_eco161014, w_eco161015, w_eco161016, w_eco161017, w_eco161018, w_eco161019, w_eco161020, w_eco161021, w_eco161022, w_eco161023, w_eco161024, w_eco161025, w_eco161026, w_eco161027, w_eco161028, w_eco161029, w_eco161030, w_eco161031, w_eco161032, w_eco161033, w_eco161034, w_eco161035, w_eco161036, w_eco161037, w_eco161038, w_eco161039, w_eco161040, w_eco161041, w_eco161042, w_eco161043, w_eco161044, w_eco161045, w_eco161046, w_eco161047, w_eco161048, w_eco161049, w_eco161050, w_eco161051, w_eco161052, w_eco161053, w_eco161054, w_eco161055, w_eco161056, w_eco161057, w_eco161058, w_eco161059, w_eco161060, w_eco161061, w_eco161062, w_eco161063, w_eco161064, w_eco161065, w_eco161066, w_eco161067, w_eco161068, w_eco161069, w_eco161070, w_eco161071, w_eco161072, w_eco161073, w_eco161074, w_eco161075, w_eco161076, w_eco161077, w_eco161078, w_eco161079, w_eco161080, w_eco161081, w_eco161082, w_eco161083, w_eco161084, w_eco161085, w_eco161086, w_eco161087, w_eco161088, w_eco161089, w_eco161090, w_eco161091, w_eco161092, w_eco161093, w_eco161094, w_eco161095, w_eco161096, w_eco161097, w_eco161098, w_eco161099, w_eco161100, w_eco161101, w_eco161102, w_eco161103, w_eco161104, w_eco161105, w_eco161106, w_eco161107, w_eco161108, w_eco161109, w_eco161110, w_eco161111, w_eco161112, w_eco161113, w_eco161114, w_eco161115, w_eco161116, w_eco161117, w_eco161118, w_eco161119, w_eco161120, w_eco161121, w_eco161122, w_eco161123, w_eco161124, w_eco161125, w_eco161126, w_eco161127, w_eco161128, w_eco161129, w_eco161130, w_eco161131, w_eco161132, w_eco161133, w_eco161134, w_eco161135, w_eco161136, w_eco161137, w_eco161138, w_eco161139, w_eco161140, w_eco161141, w_eco161142, w_eco161143, w_eco161144, w_eco161145, w_eco161146, w_eco161147, w_eco161148, w_eco161149, w_eco161150, w_eco161151, w_eco161152, w_eco161153, w_eco161154, w_eco161155, w_eco161156, w_eco161157, w_eco161158, w_eco161159, w_eco161160, w_eco161161, w_eco161162, w_eco161163, w_eco161164, w_eco161165, w_eco161166, w_eco161167, w_eco161168, w_eco161169, w_eco161170, w_eco161171, w_eco161172, w_eco161173, w_eco161174, w_eco161175, w_eco161176, w_eco161177, w_eco161178, w_eco161179, w_eco161180, w_eco161181, w_eco161182, w_eco161183, w_eco161184, w_eco161185, w_eco161186, w_eco161187, w_eco161188, w_eco161189, w_eco161190, w_eco161191, w_eco161192, w_eco161193, w_eco161194, w_eco161195, w_eco161196, w_eco161197, w_eco161198, w_eco161199, w_eco161200, w_eco161201, w_eco161202, w_eco161203, w_eco161204, w_eco161205, w_eco161206, w_eco161207, w_eco161208, w_eco161209, w_eco161210, w_eco161211, w_eco161212, w_eco161213, w_eco161214, w_eco161215, w_eco161216, w_eco161217, w_eco161218, w_eco161219, w_eco161220, w_eco161221, w_eco161222, w_eco161223, w_eco161224, w_eco161225, w_eco161226, w_eco161227, w_eco161228, w_eco161229, w_eco161230, w_eco161231, w_eco161232, w_eco161233, w_eco161234, w_eco161235, w_eco161236, w_eco161237, w_eco161238, w_eco161239, w_eco161240, w_eco161241, w_eco161242, w_eco161243, w_eco161244, w_eco161245, w_eco161246, w_eco161247, w_eco161248, w_eco161249, w_eco161250, w_eco161251, w_eco161252, w_eco161253, w_eco161254, w_eco161255, w_eco161256, w_eco161257, w_eco161258, w_eco161259, w_eco161260, w_eco161261, w_eco161262, w_eco161263, w_eco161264, w_eco161265, w_eco161266, w_eco161267, w_eco161268, w_eco161269, w_eco161270, w_eco161271, w_eco161272, w_eco161273, w_eco161274, w_eco161275, w_eco161276, w_eco161277, w_eco161278, w_eco161279, w_eco161280, w_eco161281, w_eco161282, w_eco161283, w_eco161284, w_eco161285, w_eco161286, w_eco161287, w_eco161288, w_eco161289, w_eco161290, w_eco161291, w_eco161292, w_eco161293, w_eco161294, w_eco161295, w_eco161296, w_eco161297, w_eco161298, w_eco161299, w_eco161300, w_eco161301, w_eco161302, w_eco161303, w_eco161304, w_eco161305, w_eco161306, w_eco161307, w_eco161308, w_eco161309, w_eco161310, w_eco161311, w_eco161312, w_eco161313, w_eco161314, w_eco161315, w_eco161316, w_eco161317, w_eco161318, w_eco161319, w_eco161320, w_eco161321, w_eco161322, w_eco161323, w_eco161324, w_eco161325, w_eco161326, w_eco161327, w_eco161328, w_eco161329, w_eco161330, w_eco161331, w_eco161332, w_eco161333, w_eco161334, w_eco161335, w_eco161336, w_eco161337, w_eco161338, w_eco161339, w_eco161340, w_eco161341, w_eco161342, w_eco161343, w_eco161344, w_eco161345, w_eco161346, w_eco161347, w_eco161348, w_eco161349, w_eco161350, w_eco161351, w_eco161352, w_eco161353, w_eco161354, w_eco161355, w_eco161356, w_eco161357, w_eco161358, w_eco161359, w_eco161360, w_eco161361, w_eco161362, w_eco161363, w_eco161364, w_eco161365, w_eco161366, w_eco161367, w_eco161368, w_eco161369, w_eco161370, w_eco161371, w_eco161372, w_eco161373, w_eco161374, w_eco161375, w_eco161376, w_eco161377, w_eco161378, w_eco161379, w_eco161380, w_eco161381, w_eco161382, w_eco161383, w_eco161384, w_eco161385, w_eco161386, w_eco161387, w_eco161388, w_eco161389, w_eco161390, w_eco161391, w_eco161392, w_eco161393, w_eco161394, w_eco161395, w_eco161396, w_eco161397, w_eco161398, w_eco161399, w_eco161400, w_eco161401, w_eco161402, w_eco161403, w_eco161404, w_eco161405, w_eco161406, w_eco161407, w_eco161408, w_eco161409, w_eco161410, w_eco161411, w_eco161412, w_eco161413, w_eco161414, w_eco161415, w_eco161416, w_eco161417, w_eco161418, w_eco161419, w_eco161420, w_eco161421, w_eco161422, w_eco161423, w_eco161424, w_eco161425, w_eco161426, w_eco161427, w_eco161428, w_eco161429, w_eco161430, w_eco161431, w_eco161432, w_eco161433, w_eco161434, w_eco161435, w_eco161436, w_eco161437, w_eco161438, w_eco161439, w_eco161440, w_eco161441, w_eco161442, w_eco161443, w_eco161444, w_eco161445, w_eco161446, w_eco161447, w_eco161448, w_eco161449, w_eco161450, w_eco161451, w_eco161452, w_eco161453, w_eco161454, w_eco161455, w_eco161456, w_eco161457, w_eco161458, w_eco161459, w_eco161460, w_eco161461, w_eco161462, w_eco161463, w_eco161464, w_eco161465, w_eco161466, w_eco161467, w_eco161468, w_eco161469, w_eco161470, w_eco161471, w_eco161472, w_eco161473, w_eco161474, w_eco161475, w_eco161476, w_eco161477, w_eco161478, w_eco161479, w_eco161480, w_eco161481, w_eco161482, w_eco161483, w_eco161484, w_eco161485, w_eco161486, w_eco161487, w_eco161488, w_eco161489, w_eco161490, w_eco161491, w_eco161492, w_eco161493, w_eco161494, w_eco161495, w_eco161496, w_eco161497, w_eco161498, w_eco161499, w_eco161500, w_eco161501, w_eco161502, w_eco161503, w_eco161504, w_eco161505, w_eco161506, w_eco161507, w_eco161508, w_eco161509, w_eco161510, w_eco161511, w_eco161512, w_eco161513, w_eco161514, w_eco161515, w_eco161516, w_eco161517, w_eco161518, w_eco161519, w_eco161520, w_eco161521, w_eco161522, w_eco161523, w_eco161524, w_eco161525, w_eco161526, w_eco161527, w_eco161528, w_eco161529, w_eco161530, w_eco161531, w_eco161532, w_eco161533, w_eco161534, w_eco161535, w_eco161536, w_eco161537, w_eco161538, w_eco161539, w_eco161540, w_eco161541, w_eco161542, w_eco161543, w_eco161544, w_eco161545, w_eco161546, w_eco161547, w_eco161548, w_eco161549, w_eco161550, w_eco161551, w_eco161552, w_eco161553, w_eco161554, w_eco161555, w_eco161556, w_eco161557, w_eco161558, w_eco161559, w_eco161560, w_eco161561, w_eco161562, w_eco161563, w_eco161564, w_eco161565, w_eco161566, w_eco161567, w_eco161568, w_eco161569, w_eco161570, w_eco161571, w_eco161572, w_eco161573, w_eco161574, w_eco161575, w_eco161576, w_eco161577, w_eco161578, w_eco161579, w_eco161580, w_eco161581, w_eco161582, w_eco161583, w_eco161584, w_eco161585, w_eco161586, w_eco161587, w_eco161588, w_eco161589, w_eco161590, w_eco161591, w_eco161592, w_eco161593, w_eco161594, w_eco161595, w_eco161596, w_eco161597, w_eco161598, w_eco161599, w_eco161600, w_eco161601, w_eco161602, w_eco161603, w_eco161604, w_eco161605, w_eco161606, w_eco161607, w_eco161608, w_eco161609, w_eco161610, w_eco161611, w_eco161612, w_eco161613, w_eco161614, w_eco161615, w_eco161616, w_eco161617, w_eco161618, w_eco161619, w_eco161620, w_eco161621, w_eco161622, w_eco161623, w_eco161624, w_eco161625, w_eco161626, w_eco161627, w_eco161628, w_eco161629, w_eco161630, w_eco161631, w_eco161632, w_eco161633, w_eco161634, w_eco161635, w_eco161636, w_eco161637, w_eco161638, w_eco161639, w_eco161640, w_eco161641, w_eco161642, w_eco161643, w_eco161644, w_eco161645, w_eco161646, w_eco161647, w_eco161648, w_eco161649, w_eco161650, w_eco161651, w_eco161652, w_eco161653, w_eco161654, w_eco161655, w_eco161656, w_eco161657, w_eco161658, w_eco161659, w_eco161660, w_eco161661, w_eco161662, w_eco161663, w_eco161664, w_eco161665, w_eco161666, w_eco161667, w_eco161668, w_eco161669, w_eco161670, w_eco161671, w_eco161672, w_eco161673, w_eco161674, w_eco161675, w_eco161676, w_eco161677, w_eco161678, w_eco161679, w_eco161680, w_eco161681, w_eco161682, w_eco161683, w_eco161684, w_eco161685, w_eco161686, w_eco161687, w_eco161688, w_eco161689, w_eco161690, w_eco161691, w_eco161692, w_eco161693, w_eco161694, w_eco161695, w_eco161696, w_eco161697, w_eco161698, w_eco161699, w_eco161700, w_eco161701, w_eco161702, w_eco161703, w_eco161704, w_eco161705, w_eco161706, w_eco161707, w_eco161708, w_eco161709, w_eco161710, w_eco161711, w_eco161712, w_eco161713, w_eco161714, w_eco161715, w_eco161716, w_eco161717, w_eco161718, w_eco161719, w_eco161720, w_eco161721, w_eco161722, w_eco161723, w_eco161724, w_eco161725, w_eco161726, w_eco161727, w_eco161728, w_eco161729, w_eco161730, w_eco161731, w_eco161732, w_eco161733, w_eco161734, w_eco161735, w_eco161736, w_eco161737, w_eco161738, w_eco161739, w_eco161740, w_eco161741, w_eco161742, w_eco161743, w_eco161744, w_eco161745, w_eco161746, w_eco161747, w_eco161748, w_eco161749, w_eco161750, w_eco161751, w_eco161752, w_eco161753, w_eco161754, w_eco161755, w_eco161756, w_eco161757, w_eco161758, w_eco161759, w_eco161760, w_eco161761, w_eco161762, w_eco161763, w_eco161764, w_eco161765, w_eco161766, w_eco161767, w_eco161768, w_eco161769, w_eco161770, w_eco161771, w_eco161772, w_eco161773, w_eco161774, w_eco161775, w_eco161776, w_eco161777, w_eco161778, w_eco161779, w_eco161780, w_eco161781, w_eco161782, w_eco161783, w_eco161784, w_eco161785, w_eco161786, w_eco161787, w_eco161788, w_eco161789, w_eco161790, w_eco161791, w_eco161792, w_eco161793, w_eco161794, w_eco161795, w_eco161796, w_eco161797, w_eco161798, w_eco161799, w_eco161800, w_eco161801, w_eco161802, w_eco161803, w_eco161804, w_eco161805, w_eco161806, w_eco161807, w_eco161808, w_eco161809, w_eco161810, w_eco161811, w_eco161812, w_eco161813, w_eco161814, w_eco161815, w_eco161816, w_eco161817, w_eco161818, w_eco161819, w_eco161820, w_eco161821, w_eco161822, w_eco161823, w_eco161824, w_eco161825, w_eco161826, w_eco161827, w_eco161828, w_eco161829, w_eco161830, w_eco161831, w_eco161832, w_eco161833, w_eco161834, w_eco161835, w_eco161836, w_eco161837, w_eco161838, w_eco161839, w_eco161840, w_eco161841, w_eco161842, w_eco161843, w_eco161844, w_eco161845, w_eco161846, w_eco161847, w_eco161848, w_eco161849, w_eco161850, w_eco161851, w_eco161852, w_eco161853, w_eco161854, w_eco161855, w_eco161856, w_eco161857, w_eco161858, w_eco161859, w_eco161860, w_eco161861, w_eco161862, w_eco161863, w_eco161864, w_eco161865, w_eco161866, w_eco161867, w_eco161868, w_eco161869, w_eco161870, w_eco161871, w_eco161872, w_eco161873, w_eco161874, w_eco161875, w_eco161876, w_eco161877, w_eco161878, w_eco161879, w_eco161880, w_eco161881, w_eco161882, w_eco161883, w_eco161884, w_eco161885, w_eco161886, w_eco161887, w_eco161888, w_eco161889, w_eco161890, w_eco161891, w_eco161892, w_eco161893, w_eco161894, w_eco161895, w_eco161896, w_eco161897, w_eco161898, w_eco161899, w_eco161900, w_eco161901, w_eco161902, w_eco161903, w_eco161904, w_eco161905, w_eco161906, w_eco161907, w_eco161908, w_eco161909, w_eco161910, w_eco161911, w_eco161912, w_eco161913, w_eco161914, w_eco161915, w_eco161916, w_eco161917, w_eco161918, w_eco161919, w_eco161920, w_eco161921, w_eco161922, w_eco161923, w_eco161924, w_eco161925, w_eco161926, w_eco161927, w_eco161928, w_eco161929, w_eco161930, w_eco161931, w_eco161932, w_eco161933, w_eco161934, w_eco161935, w_eco161936, w_eco161937, w_eco161938, w_eco161939, w_eco161940, w_eco161941, w_eco161942, w_eco161943, w_eco161944, w_eco161945, w_eco161946, w_eco161947, w_eco161948, w_eco161949, w_eco161950, w_eco161951, w_eco161952, w_eco161953, w_eco161954, w_eco161955, w_eco161956, w_eco161957, w_eco161958, w_eco161959, w_eco161960, w_eco161961, w_eco161962, w_eco161963, w_eco161964, w_eco161965, w_eco161966, w_eco161967, w_eco161968, w_eco161969, w_eco161970, w_eco161971, w_eco161972, w_eco161973, w_eco161974, w_eco161975, w_eco161976, w_eco161977, w_eco161978, w_eco161979, w_eco161980, w_eco161981, w_eco161982, w_eco161983, w_eco161984, w_eco161985, w_eco161986, w_eco161987, w_eco161988, w_eco161989, w_eco161990, w_eco161991, w_eco161992, w_eco161993, w_eco161994, w_eco161995, w_eco161996, w_eco161997, w_eco161998, w_eco161999, w_eco162000, w_eco162001, w_eco162002, w_eco162003, w_eco162004, w_eco162005, w_eco162006, w_eco162007, w_eco162008, w_eco162009, w_eco162010, w_eco162011, w_eco162012, w_eco162013, w_eco162014, w_eco162015, w_eco162016, w_eco162017, w_eco162018, w_eco162019, w_eco162020, w_eco162021, w_eco162022, w_eco162023, w_eco162024, w_eco162025, w_eco162026, w_eco162027, w_eco162028, w_eco162029, w_eco162030, w_eco162031, w_eco162032, w_eco162033, w_eco162034, w_eco162035, w_eco162036, w_eco162037, w_eco162038, w_eco162039, w_eco162040, w_eco162041, w_eco162042, w_eco162043, w_eco162044, w_eco162045, w_eco162046, w_eco162047, w_eco162048, w_eco162049, w_eco162050, w_eco162051, w_eco162052, w_eco162053, w_eco162054, w_eco162055, w_eco162056, w_eco162057, w_eco162058, w_eco162059, w_eco162060, w_eco162061, w_eco162062, w_eco162063, w_eco162064, w_eco162065, w_eco162066, w_eco162067, w_eco162068, w_eco162069, w_eco162070, w_eco162071, w_eco162072, w_eco162073, w_eco162074, w_eco162075, w_eco162076, w_eco162077, w_eco162078, w_eco162079, w_eco162080, w_eco162081, w_eco162082, w_eco162083, w_eco162084, w_eco162085, w_eco162086, w_eco162087, w_eco162088, w_eco162089, w_eco162090, w_eco162091, w_eco162092, w_eco162093, w_eco162094, w_eco162095, w_eco162096, w_eco162097, w_eco162098, w_eco162099, w_eco162100, w_eco162101, w_eco162102, w_eco162103, w_eco162104, w_eco162105, w_eco162106, w_eco162107, w_eco162108, w_eco162109, w_eco162110, w_eco162111, w_eco162112, w_eco162113, w_eco162114, w_eco162115, w_eco162116, w_eco162117, w_eco162118, w_eco162119, w_eco162120, w_eco162121, w_eco162122, w_eco162123, w_eco162124, w_eco162125, w_eco162126, w_eco162127, w_eco162128, w_eco162129, w_eco162130, w_eco162131, w_eco162132, w_eco162133, w_eco162134, w_eco162135, w_eco162136, w_eco162137, w_eco162138, w_eco162139, w_eco162140, w_eco162141, w_eco162142, w_eco162143, w_eco162144, w_eco162145, w_eco162146, w_eco162147, w_eco162148, w_eco162149, w_eco162150, w_eco162151, w_eco162152, w_eco162153, w_eco162154, w_eco162155, w_eco162156, w_eco162157, w_eco162158, w_eco162159, w_eco162160, w_eco162161, w_eco162162, w_eco162163, w_eco162164, w_eco162165, w_eco162166, w_eco162167, w_eco162168, w_eco162169, w_eco162170, w_eco162171, w_eco162172, w_eco162173, w_eco162174, w_eco162175, w_eco162176, w_eco162177, w_eco162178, w_eco162179, w_eco162180, w_eco162181, w_eco162182, w_eco162183, w_eco162184, w_eco162185, w_eco162186, w_eco162187, w_eco162188, w_eco162189, w_eco162190, w_eco162191, w_eco162192, w_eco162193, w_eco162194, w_eco162195, w_eco162196, w_eco162197, w_eco162198, w_eco162199, w_eco162200, w_eco162201, w_eco162202, w_eco162203, w_eco162204, w_eco162205, w_eco162206, w_eco162207, w_eco162208, w_eco162209, w_eco162210, w_eco162211, w_eco162212, w_eco162213, w_eco162214, w_eco162215, w_eco162216, w_eco162217, w_eco162218, w_eco162219, w_eco162220, w_eco162221, w_eco162222, w_eco162223, w_eco162224, w_eco162225, w_eco162226, w_eco162227, w_eco162228, w_eco162229, w_eco162230, w_eco162231, w_eco162232, w_eco162233, w_eco162234, w_eco162235, w_eco162236, w_eco162237, w_eco162238, w_eco162239, w_eco162240, w_eco162241, w_eco162242, w_eco162243, w_eco162244, w_eco162245, w_eco162246, w_eco162247, w_eco162248, w_eco162249, w_eco162250, w_eco162251, w_eco162252, w_eco162253, w_eco162254, w_eco162255, w_eco162256, w_eco162257, w_eco162258, w_eco162259, w_eco162260, w_eco162261, w_eco162262, w_eco162263, w_eco162264, w_eco162265, w_eco162266, w_eco162267, w_eco162268, w_eco162269, w_eco162270, w_eco162271, w_eco162272, w_eco162273, w_eco162274, w_eco162275, w_eco162276, w_eco162277, w_eco162278, w_eco162279, w_eco162280, w_eco162281, w_eco162282, w_eco162283, w_eco162284, w_eco162285, w_eco162286, w_eco162287, w_eco162288, w_eco162289, w_eco162290, w_eco162291, w_eco162292, w_eco162293, w_eco162294, w_eco162295, w_eco162296, w_eco162297, w_eco162298, w_eco162299, w_eco162300, w_eco162301, w_eco162302, w_eco162303, w_eco162304, w_eco162305, w_eco162306, w_eco162307, w_eco162308, w_eco162309, w_eco162310, w_eco162311, w_eco162312, w_eco162313, w_eco162314, w_eco162315, w_eco162316, w_eco162317, w_eco162318, w_eco162319, w_eco162320, w_eco162321, w_eco162322, w_eco162323, w_eco162324, w_eco162325, w_eco162326, w_eco162327, w_eco162328, w_eco162329, w_eco162330, w_eco162331, w_eco162332, w_eco162333, w_eco162334, w_eco162335, w_eco162336, w_eco162337, w_eco162338, w_eco162339, w_eco162340, w_eco162341, w_eco162342, w_eco162343, w_eco162344, w_eco162345, w_eco162346, w_eco162347, w_eco162348, w_eco162349, w_eco162350, w_eco162351, w_eco162352, w_eco162353, w_eco162354, w_eco162355, w_eco162356, w_eco162357, w_eco162358, w_eco162359, w_eco162360, w_eco162361, w_eco162362, w_eco162363, w_eco162364, w_eco162365, w_eco162366, w_eco162367, w_eco162368, w_eco162369, w_eco162370, w_eco162371, w_eco162372, w_eco162373, w_eco162374, w_eco162375, w_eco162376, w_eco162377, w_eco162378, w_eco162379, w_eco162380, w_eco162381, w_eco162382, w_eco162383, w_eco162384, w_eco162385, w_eco162386, w_eco162387, w_eco162388, w_eco162389, w_eco162390, w_eco162391, w_eco162392, w_eco162393, w_eco162394, w_eco162395, w_eco162396, w_eco162397, w_eco162398, w_eco162399, w_eco162400, w_eco162401, w_eco162402, w_eco162403, w_eco162404, w_eco162405, w_eco162406, w_eco162407, w_eco162408, w_eco162409, w_eco162410, w_eco162411, w_eco162412, w_eco162413, w_eco162414, w_eco162415, w_eco162416, w_eco162417, w_eco162418, w_eco162419, w_eco162420, w_eco162421, w_eco162422, w_eco162423, w_eco162424, w_eco162425, w_eco162426, w_eco162427, w_eco162428, w_eco162429, w_eco162430, w_eco162431, w_eco162432, w_eco162433, w_eco162434, w_eco162435, w_eco162436, w_eco162437, w_eco162438, w_eco162439, w_eco162440, w_eco162441, w_eco162442, w_eco162443, w_eco162444, w_eco162445, w_eco162446, w_eco162447, w_eco162448, w_eco162449, w_eco162450, w_eco162451, w_eco162452, w_eco162453, w_eco162454, w_eco162455, w_eco162456, w_eco162457, w_eco162458, w_eco162459, w_eco162460, w_eco162461, w_eco162462, w_eco162463, w_eco162464, w_eco162465, w_eco162466, w_eco162467, w_eco162468, w_eco162469, w_eco162470, w_eco162471, w_eco162472, w_eco162473, w_eco162474, w_eco162475, w_eco162476, w_eco162477, w_eco162478, w_eco162479, w_eco162480, w_eco162481, w_eco162482, w_eco162483, w_eco162484, w_eco162485, w_eco162486, w_eco162487, w_eco162488, w_eco162489, w_eco162490, w_eco162491, w_eco162492, w_eco162493, w_eco162494, w_eco162495, w_eco162496, w_eco162497, w_eco162498, w_eco162499, w_eco162500, w_eco162501, w_eco162502, w_eco162503, w_eco162504, w_eco162505, w_eco162506, w_eco162507, w_eco162508, w_eco162509, w_eco162510, w_eco162511, w_eco162512, w_eco162513, w_eco162514, w_eco162515, w_eco162516, w_eco162517, w_eco162518, w_eco162519, w_eco162520, w_eco162521, w_eco162522, w_eco162523, w_eco162524, w_eco162525, w_eco162526, w_eco162527, w_eco162528, w_eco162529, w_eco162530, w_eco162531, w_eco162532, w_eco162533, w_eco162534, w_eco162535, w_eco162536, w_eco162537, w_eco162538, w_eco162539, w_eco162540, w_eco162541, w_eco162542, w_eco162543, w_eco162544, w_eco162545, w_eco162546, w_eco162547, w_eco162548, w_eco162549, w_eco162550, w_eco162551, w_eco162552, w_eco162553, w_eco162554, w_eco162555, w_eco162556, w_eco162557, w_eco162558, w_eco162559, w_eco162560, w_eco162561, w_eco162562, w_eco162563, w_eco162564, w_eco162565, w_eco162566, w_eco162567, w_eco162568, w_eco162569, w_eco162570, w_eco162571, w_eco162572, w_eco162573, w_eco162574, w_eco162575, w_eco162576, w_eco162577, w_eco162578, w_eco162579, w_eco162580, w_eco162581, w_eco162582, w_eco162583, w_eco162584, w_eco162585, w_eco162586, w_eco162587, w_eco162588, w_eco162589, w_eco162590, w_eco162591, w_eco162592, w_eco162593, w_eco162594, w_eco162595, w_eco162596, w_eco162597, w_eco162598, w_eco162599, w_eco162600, w_eco162601, w_eco162602, w_eco162603, w_eco162604, w_eco162605, w_eco162606, w_eco162607, w_eco162608, w_eco162609, w_eco162610, w_eco162611, w_eco162612, w_eco162613, w_eco162614, w_eco162615, w_eco162616, w_eco162617, w_eco162618, w_eco162619, w_eco162620, w_eco162621, w_eco162622, w_eco162623, w_eco162624, w_eco162625, w_eco162626, w_eco162627, w_eco162628, w_eco162629, w_eco162630, w_eco162631, w_eco162632, w_eco162633, w_eco162634, w_eco162635, w_eco162636, w_eco162637, w_eco162638, w_eco162639, w_eco162640, w_eco162641, w_eco162642, w_eco162643, w_eco162644, w_eco162645, w_eco162646, w_eco162647, w_eco162648, w_eco162649, w_eco162650, w_eco162651, w_eco162652, w_eco162653, w_eco162654, w_eco162655, w_eco162656, w_eco162657, w_eco162658, w_eco162659, w_eco162660, w_eco162661, w_eco162662, w_eco162663, w_eco162664, w_eco162665, w_eco162666, w_eco162667, w_eco162668, w_eco162669, w_eco162670, w_eco162671, w_eco162672, w_eco162673, w_eco162674, w_eco162675, w_eco162676, w_eco162677, w_eco162678, w_eco162679, w_eco162680, w_eco162681, w_eco162682, w_eco162683, w_eco162684, w_eco162685, w_eco162686, w_eco162687, w_eco162688, w_eco162689, w_eco162690, w_eco162691, w_eco162692, w_eco162693, w_eco162694, w_eco162695, w_eco162696, w_eco162697, w_eco162698, w_eco162699, w_eco162700, w_eco162701, w_eco162702, w_eco162703, w_eco162704, w_eco162705, w_eco162706, w_eco162707, w_eco162708, w_eco162709, w_eco162710, w_eco162711, w_eco162712, w_eco162713, w_eco162714, w_eco162715, w_eco162716, w_eco162717, w_eco162718, w_eco162719, w_eco162720, w_eco162721, w_eco162722, w_eco162723, w_eco162724, w_eco162725, w_eco162726, w_eco162727, w_eco162728, w_eco162729, w_eco162730, w_eco162731, w_eco162732, w_eco162733, w_eco162734, w_eco162735, w_eco162736, w_eco162737, w_eco162738, w_eco162739, w_eco162740, w_eco162741, w_eco162742, w_eco162743, w_eco162744, w_eco162745, w_eco162746, w_eco162747, w_eco162748, w_eco162749, w_eco162750, w_eco162751, w_eco162752, w_eco162753, w_eco162754, w_eco162755, w_eco162756, w_eco162757, w_eco162758, w_eco162759, w_eco162760, w_eco162761, w_eco162762, w_eco162763, w_eco162764, w_eco162765, w_eco162766, w_eco162767, w_eco162768, w_eco162769, w_eco162770, w_eco162771, w_eco162772, w_eco162773, w_eco162774, w_eco162775, w_eco162776, w_eco162777, w_eco162778, w_eco162779, w_eco162780, w_eco162781, w_eco162782, w_eco162783, w_eco162784, w_eco162785, w_eco162786, w_eco162787, w_eco162788, w_eco162789, w_eco162790, w_eco162791, w_eco162792, w_eco162793, w_eco162794, w_eco162795, w_eco162796, w_eco162797, w_eco162798, w_eco162799, w_eco162800, w_eco162801, w_eco162802, w_eco162803, w_eco162804, w_eco162805, w_eco162806, w_eco162807, w_eco162808, w_eco162809, w_eco162810, w_eco162811, w_eco162812, w_eco162813, w_eco162814, w_eco162815, w_eco162816, w_eco162817, w_eco162818, w_eco162819, w_eco162820, w_eco162821, w_eco162822, w_eco162823, w_eco162824, w_eco162825, w_eco162826, w_eco162827, w_eco162828, w_eco162829, w_eco162830, w_eco162831, w_eco162832, w_eco162833, w_eco162834, w_eco162835, w_eco162836, w_eco162837, w_eco162838, w_eco162839, w_eco162840, w_eco162841, w_eco162842, w_eco162843, w_eco162844, w_eco162845, w_eco162846, w_eco162847, w_eco162848, w_eco162849, w_eco162850, w_eco162851, w_eco162852, w_eco162853, w_eco162854, w_eco162855, w_eco162856, w_eco162857, w_eco162858, w_eco162859, w_eco162860, w_eco162861, w_eco162862, w_eco162863, w_eco162864, w_eco162865, w_eco162866, w_eco162867, w_eco162868, w_eco162869, w_eco162870, w_eco162871, w_eco162872, w_eco162873, w_eco162874, w_eco162875, w_eco162876, w_eco162877, w_eco162878, w_eco162879, w_eco162880, w_eco162881, w_eco162882, w_eco162883, w_eco162884, w_eco162885, w_eco162886, w_eco162887, w_eco162888, w_eco162889, w_eco162890, w_eco162891, w_eco162892, w_eco162893, w_eco162894, w_eco162895, w_eco162896, w_eco162897, w_eco162898, w_eco162899, w_eco162900, w_eco162901, w_eco162902, w_eco162903, w_eco162904, w_eco162905, w_eco162906, w_eco162907, w_eco162908, w_eco162909, w_eco162910, w_eco162911, w_eco162912, w_eco162913, w_eco162914, w_eco162915, w_eco162916, w_eco162917, w_eco162918, w_eco162919, w_eco162920, w_eco162921, w_eco162922, w_eco162923, w_eco162924, w_eco162925, w_eco162926, w_eco162927, w_eco162928, w_eco162929, w_eco162930, w_eco162931, w_eco162932, w_eco162933, w_eco162934, w_eco162935, w_eco162936, w_eco162937, w_eco162938, w_eco162939, w_eco162940, w_eco162941, w_eco162942, w_eco162943, w_eco162944, w_eco162945, w_eco162946, w_eco162947, w_eco162948, w_eco162949, w_eco162950, w_eco162951, w_eco162952, w_eco162953, w_eco162954, w_eco162955, w_eco162956, w_eco162957, w_eco162958, w_eco162959, w_eco162960, w_eco162961, w_eco162962, w_eco162963, w_eco162964, w_eco162965, w_eco162966, w_eco162967, w_eco162968, w_eco162969, w_eco162970, w_eco162971, w_eco162972, w_eco162973, w_eco162974, w_eco162975, w_eco162976, w_eco162977, w_eco162978, w_eco162979, w_eco162980, w_eco162981, w_eco162982, w_eco162983, w_eco162984, w_eco162985, w_eco162986, w_eco162987, w_eco162988, w_eco162989, w_eco162990, w_eco162991, w_eco162992, w_eco162993, w_eco162994, w_eco162995, w_eco162996, w_eco162997, w_eco162998, w_eco162999, w_eco163000, w_eco163001, w_eco163002, w_eco163003, w_eco163004, w_eco163005, w_eco163006, w_eco163007, w_eco163008, w_eco163009, w_eco163010, w_eco163011, w_eco163012, w_eco163013, w_eco163014, w_eco163015, w_eco163016, w_eco163017, w_eco163018, w_eco163019, w_eco163020, w_eco163021, w_eco163022, w_eco163023, w_eco163024, w_eco163025, w_eco163026, w_eco163027, w_eco163028, w_eco163029, w_eco163030, w_eco163031, w_eco163032, w_eco163033, w_eco163034, w_eco163035, w_eco163036, w_eco163037, w_eco163038, w_eco163039, w_eco163040, w_eco163041, w_eco163042, w_eco163043, w_eco163044, w_eco163045, w_eco163046, w_eco163047, w_eco163048, w_eco163049, w_eco163050, w_eco163051, w_eco163052, w_eco163053, w_eco163054, w_eco163055, w_eco163056, w_eco163057, w_eco163058, w_eco163059, w_eco163060, w_eco163061, w_eco163062, w_eco163063, w_eco163064, w_eco163065, w_eco163066, w_eco163067, w_eco163068, w_eco163069, w_eco163070, w_eco163071, w_eco163072, w_eco163073, w_eco163074, w_eco163075, w_eco163076, w_eco163077, w_eco163078, w_eco163079, w_eco163080, w_eco163081, w_eco163082, w_eco163083, w_eco163084, w_eco163085, w_eco163086, w_eco163087, w_eco163088, w_eco163089, w_eco163090, w_eco163091, w_eco163092, w_eco163093, w_eco163094, w_eco163095, w_eco163096, w_eco163097, w_eco163098, w_eco163099, w_eco163100, w_eco163101, w_eco163102, w_eco163103, w_eco163104, w_eco163105, w_eco163106, w_eco163107, w_eco163108, w_eco163109, w_eco163110, w_eco163111, w_eco163112, w_eco163113, w_eco163114, w_eco163115, w_eco163116, w_eco163117, w_eco163118, w_eco163119, w_eco163120, w_eco163121, w_eco163122, w_eco163123, w_eco163124, w_eco163125, w_eco163126, w_eco163127, w_eco163128, w_eco163129, w_eco163130, w_eco163131, w_eco163132, w_eco163133, w_eco163134, w_eco163135, w_eco163136, w_eco163137, w_eco163138, w_eco163139, w_eco163140, w_eco163141, w_eco163142, w_eco163143, w_eco163144, w_eco163145, w_eco163146, w_eco163147, w_eco163148, w_eco163149, w_eco163150, w_eco163151, w_eco163152, w_eco163153, w_eco163154, w_eco163155, w_eco163156, w_eco163157, w_eco163158, w_eco163159, w_eco163160, w_eco163161, w_eco163162, w_eco163163, w_eco163164, w_eco163165, w_eco163166, w_eco163167, w_eco163168, w_eco163169, w_eco163170, w_eco163171, w_eco163172, w_eco163173, w_eco163174, w_eco163175, w_eco163176, w_eco163177, w_eco163178, w_eco163179, w_eco163180, w_eco163181, w_eco163182, w_eco163183, w_eco163184, w_eco163185, w_eco163186, w_eco163187, w_eco163188, w_eco163189, w_eco163190, w_eco163191, w_eco163192, w_eco163193, w_eco163194, w_eco163195, w_eco163196, w_eco163197, w_eco163198, w_eco163199, w_eco163200, w_eco163201, w_eco163202, w_eco163203, w_eco163204, w_eco163205, w_eco163206, w_eco163207, w_eco163208, w_eco163209, w_eco163210, w_eco163211, w_eco163212, w_eco163213, w_eco163214, w_eco163215, w_eco163216, w_eco163217, w_eco163218, w_eco163219, w_eco163220, w_eco163221, w_eco163222, w_eco163223, w_eco163224, w_eco163225, w_eco163226, w_eco163227, w_eco163228, w_eco163229, w_eco163230, w_eco163231, w_eco163232, w_eco163233, w_eco163234, w_eco163235, w_eco163236, w_eco163237, w_eco163238, w_eco163239, w_eco163240, w_eco163241, w_eco163242, w_eco163243, w_eco163244, w_eco163245, w_eco163246, w_eco163247, w_eco163248, w_eco163249, w_eco163250, w_eco163251, w_eco163252, w_eco163253, w_eco163254, w_eco163255, w_eco163256, w_eco163257, w_eco163258, w_eco163259, w_eco163260, w_eco163261, w_eco163262, w_eco163263, w_eco163264, w_eco163265, w_eco163266, w_eco163267, w_eco163268, w_eco163269, w_eco163270, w_eco163271, w_eco163272, w_eco163273, w_eco163274, w_eco163275, w_eco163276, w_eco163277, w_eco163278, w_eco163279, w_eco163280, w_eco163281, w_eco163282, w_eco163283, w_eco163284, w_eco163285, w_eco163286, w_eco163287, w_eco163288, w_eco163289, w_eco163290, w_eco163291, w_eco163292, w_eco163293, w_eco163294, w_eco163295, w_eco163296, w_eco163297, w_eco163298, w_eco163299, w_eco163300, w_eco163301, w_eco163302, w_eco163303, w_eco163304, w_eco163305, w_eco163306, w_eco163307, w_eco163308, w_eco163309, w_eco163310, w_eco163311, w_eco163312, w_eco163313, w_eco163314, w_eco163315, w_eco163316, w_eco163317, w_eco163318, w_eco163319, w_eco163320, w_eco163321, w_eco163322, w_eco163323, w_eco163324, w_eco163325, w_eco163326, w_eco163327, w_eco163328, w_eco163329, w_eco163330, w_eco163331, w_eco163332, w_eco163333, w_eco163334, w_eco163335, w_eco163336, w_eco163337, w_eco163338, w_eco163339, w_eco163340, w_eco163341, w_eco163342, w_eco163343, w_eco163344, w_eco163345, w_eco163346, w_eco163347, w_eco163348, w_eco163349, w_eco163350, w_eco163351, w_eco163352, w_eco163353, w_eco163354, w_eco163355, w_eco163356, w_eco163357, w_eco163358, w_eco163359, w_eco163360, w_eco163361, w_eco163362, w_eco163363, w_eco163364, w_eco163365, w_eco163366, w_eco163367, w_eco163368, w_eco163369, w_eco163370, w_eco163371, w_eco163372, w_eco163373, w_eco163374, w_eco163375, w_eco163376, w_eco163377, w_eco163378, w_eco163379, w_eco163380, w_eco163381, w_eco163382, w_eco163383, w_eco163384, w_eco163385, w_eco163386, w_eco163387, w_eco163388, w_eco163389, w_eco163390, w_eco163391, w_eco163392, w_eco163393, w_eco163394, w_eco163395, w_eco163396, w_eco163397, w_eco163398, w_eco163399, w_eco163400, w_eco163401, w_eco163402, w_eco163403, w_eco163404, w_eco163405, w_eco163406, w_eco163407, w_eco163408, w_eco163409, w_eco163410, w_eco163411, w_eco163412, w_eco163413, w_eco163414, w_eco163415, w_eco163416, w_eco163417, w_eco163418, w_eco163419, w_eco163420, w_eco163421, w_eco163422, w_eco163423, w_eco163424, w_eco163425, w_eco163426, w_eco163427, w_eco163428, w_eco163429, w_eco163430, w_eco163431, w_eco163432, w_eco163433, w_eco163434, w_eco163435, w_eco163436, w_eco163437, w_eco163438, w_eco163439, w_eco163440, w_eco163441, w_eco163442, w_eco163443, w_eco163444, w_eco163445, w_eco163446, w_eco163447, w_eco163448, w_eco163449, w_eco163450, w_eco163451, w_eco163452, w_eco163453, w_eco163454, w_eco163455, w_eco163456, w_eco163457, w_eco163458, w_eco163459, w_eco163460, w_eco163461, w_eco163462, w_eco163463, w_eco163464, w_eco163465, w_eco163466, w_eco163467, w_eco163468, w_eco163469, w_eco163470, w_eco163471, w_eco163472, w_eco163473, w_eco163474, w_eco163475, w_eco163476, w_eco163477, w_eco163478, w_eco163479, w_eco163480, w_eco163481, w_eco163482, w_eco163483, w_eco163484, w_eco163485, w_eco163486, w_eco163487, w_eco163488, w_eco163489, w_eco163490, w_eco163491, w_eco163492, w_eco163493, w_eco163494, w_eco163495, w_eco163496, w_eco163497, w_eco163498, w_eco163499, w_eco163500, w_eco163501, w_eco163502, w_eco163503, w_eco163504, w_eco163505, w_eco163506, w_eco163507, w_eco163508, w_eco163509, w_eco163510, w_eco163511, w_eco163512, w_eco163513, w_eco163514, w_eco163515, w_eco163516, w_eco163517, w_eco163518, w_eco163519, w_eco163520, w_eco163521, w_eco163522, w_eco163523, w_eco163524, w_eco163525, w_eco163526, w_eco163527, w_eco163528, w_eco163529, w_eco163530, w_eco163531, w_eco163532, w_eco163533, w_eco163534, w_eco163535, w_eco163536, w_eco163537, w_eco163538, w_eco163539, w_eco163540, w_eco163541, w_eco163542, w_eco163543, w_eco163544, w_eco163545, w_eco163546, w_eco163547, w_eco163548, w_eco163549, w_eco163550, w_eco163551, w_eco163552, w_eco163553, w_eco163554, w_eco163555, w_eco163556, w_eco163557, w_eco163558, w_eco163559, w_eco163560, w_eco163561, w_eco163562, w_eco163563, w_eco163564, w_eco163565, w_eco163566, w_eco163567, w_eco163568, w_eco163569, w_eco163570, w_eco163571, w_eco163572, w_eco163573, w_eco163574, w_eco163575, w_eco163576, w_eco163577, w_eco163578, w_eco163579, w_eco163580, w_eco163581, w_eco163582, w_eco163583, w_eco163584, w_eco163585, w_eco163586, w_eco163587, w_eco163588, w_eco163589, w_eco163590, w_eco163591, w_eco163592, w_eco163593, w_eco163594, w_eco163595, w_eco163596, w_eco163597, w_eco163598, w_eco163599, w_eco163600, w_eco163601, w_eco163602, w_eco163603, w_eco163604, w_eco163605, w_eco163606, w_eco163607, w_eco163608, w_eco163609, w_eco163610, w_eco163611, w_eco163612, w_eco163613, w_eco163614, w_eco163615, w_eco163616, w_eco163617, w_eco163618, w_eco163619, w_eco163620, w_eco163621, w_eco163622, w_eco163623, w_eco163624, w_eco163625, w_eco163626, w_eco163627, w_eco163628, w_eco163629, w_eco163630, w_eco163631, w_eco163632, w_eco163633, w_eco163634, w_eco163635, w_eco163636, w_eco163637, w_eco163638, w_eco163639, w_eco163640, w_eco163641, w_eco163642, w_eco163643, w_eco163644, w_eco163645, w_eco163646, w_eco163647, w_eco163648, w_eco163649, w_eco163650, w_eco163651, w_eco163652, w_eco163653, w_eco163654, w_eco163655, w_eco163656, w_eco163657, w_eco163658, w_eco163659, w_eco163660, w_eco163661, w_eco163662, w_eco163663, w_eco163664, w_eco163665, w_eco163666, w_eco163667, w_eco163668, w_eco163669, w_eco163670, w_eco163671, w_eco163672, w_eco163673, w_eco163674, w_eco163675, w_eco163676, w_eco163677, w_eco163678, w_eco163679, w_eco163680, w_eco163681, w_eco163682, w_eco163683, w_eco163684, w_eco163685, w_eco163686, w_eco163687, w_eco163688, w_eco163689, w_eco163690, w_eco163691, w_eco163692, w_eco163693, w_eco163694, w_eco163695, w_eco163696, w_eco163697, w_eco163698, w_eco163699, w_eco163700, w_eco163701, w_eco163702, w_eco163703, w_eco163704, w_eco163705, w_eco163706, w_eco163707, w_eco163708, w_eco163709, w_eco163710, w_eco163711, w_eco163712, w_eco163713, w_eco163714, w_eco163715, w_eco163716, w_eco163717, w_eco163718, w_eco163719, w_eco163720, w_eco163721, w_eco163722, w_eco163723, w_eco163724, w_eco163725, w_eco163726, w_eco163727, w_eco163728, w_eco163729, w_eco163730, w_eco163731, w_eco163732, w_eco163733, w_eco163734, w_eco163735, w_eco163736, w_eco163737, w_eco163738, w_eco163739, w_eco163740, w_eco163741, w_eco163742, w_eco163743, w_eco163744, w_eco163745, w_eco163746, w_eco163747, w_eco163748, w_eco163749, w_eco163750, w_eco163751, w_eco163752, w_eco163753, w_eco163754, w_eco163755, w_eco163756, w_eco163757, w_eco163758, w_eco163759, w_eco163760, w_eco163761, w_eco163762, w_eco163763, w_eco163764, w_eco163765, w_eco163766, w_eco163767, w_eco163768, w_eco163769, w_eco163770, w_eco163771, w_eco163772, w_eco163773, w_eco163774, w_eco163775, w_eco163776, w_eco163777, w_eco163778, w_eco163779, w_eco163780, w_eco163781, w_eco163782, w_eco163783, w_eco163784, w_eco163785, w_eco163786, w_eco163787, w_eco163788, w_eco163789, w_eco163790, w_eco163791, w_eco163792, w_eco163793, w_eco163794, w_eco163795, w_eco163796, w_eco163797, w_eco163798, w_eco163799, w_eco163800, w_eco163801, w_eco163802, w_eco163803, w_eco163804, w_eco163805, w_eco163806, w_eco163807, w_eco163808, w_eco163809, w_eco163810, w_eco163811, w_eco163812, w_eco163813, w_eco163814, w_eco163815, w_eco163816, w_eco163817, w_eco163818, w_eco163819, w_eco163820, w_eco163821, w_eco163822, w_eco163823, w_eco163824, w_eco163825, w_eco163826, w_eco163827, w_eco163828, w_eco163829, w_eco163830, w_eco163831, w_eco163832, w_eco163833, w_eco163834, w_eco163835, w_eco163836, w_eco163837, w_eco163838, w_eco163839, w_eco163840, w_eco163841, w_eco163842, w_eco163843, w_eco163844, w_eco163845, w_eco163846, w_eco163847, w_eco163848, w_eco163849, w_eco163850, w_eco163851, w_eco163852, w_eco163853, w_eco163854, w_eco163855, w_eco163856, w_eco163857, w_eco163858, w_eco163859, w_eco163860, w_eco163861, w_eco163862, w_eco163863, w_eco163864, w_eco163865, w_eco163866, w_eco163867, w_eco163868, w_eco163869, w_eco163870, w_eco163871, w_eco163872, w_eco163873, w_eco163874, w_eco163875, w_eco163876, w_eco163877, w_eco163878, w_eco163879, w_eco163880, w_eco163881, w_eco163882, w_eco163883, w_eco163884, w_eco163885, w_eco163886, w_eco163887, w_eco163888, w_eco163889, w_eco163890, w_eco163891, w_eco163892, w_eco163893, w_eco163894, w_eco163895, w_eco163896, w_eco163897, w_eco163898, w_eco163899, w_eco163900, w_eco163901, w_eco163902, w_eco163903, w_eco163904, w_eco163905, w_eco163906, w_eco163907, w_eco163908, w_eco163909, w_eco163910, w_eco163911, w_eco163912, w_eco163913, w_eco163914, w_eco163915, w_eco163916, w_eco163917, w_eco163918, w_eco163919, w_eco163920, w_eco163921, w_eco163922, w_eco163923, w_eco163924, w_eco163925, w_eco163926, w_eco163927, w_eco163928, w_eco163929, w_eco163930, w_eco163931, w_eco163932, w_eco163933, w_eco163934, w_eco163935, w_eco163936, w_eco163937, w_eco163938, w_eco163939, w_eco163940, w_eco163941, w_eco163942, w_eco163943, w_eco163944, w_eco163945, w_eco163946, w_eco163947, w_eco163948, w_eco163949, w_eco163950, w_eco163951, w_eco163952, w_eco163953, w_eco163954, w_eco163955, w_eco163956, w_eco163957, w_eco163958, w_eco163959, w_eco163960, w_eco163961, w_eco163962, w_eco163963, w_eco163964, w_eco163965, w_eco163966, w_eco163967, w_eco163968, w_eco163969, w_eco163970, w_eco163971, w_eco163972, w_eco163973, w_eco163974, w_eco163975, w_eco163976, w_eco163977, w_eco163978, w_eco163979, w_eco163980, w_eco163981, w_eco163982, w_eco163983, w_eco163984, w_eco163985, w_eco163986, w_eco163987, w_eco163988, w_eco163989, w_eco163990, w_eco163991, w_eco163992, w_eco163993, w_eco163994, w_eco163995, w_eco163996, w_eco163997, w_eco163998, w_eco163999, w_eco164000, w_eco164001, w_eco164002, w_eco164003, w_eco164004, w_eco164005, w_eco164006, w_eco164007, w_eco164008, w_eco164009, w_eco164010, w_eco164011, w_eco164012, w_eco164013, w_eco164014, w_eco164015, w_eco164016, w_eco164017, w_eco164018, w_eco164019, w_eco164020, w_eco164021, w_eco164022, w_eco164023, w_eco164024, w_eco164025, w_eco164026, w_eco164027, w_eco164028, w_eco164029, w_eco164030, w_eco164031, w_eco164032, w_eco164033, w_eco164034, w_eco164035, w_eco164036, w_eco164037, w_eco164038, w_eco164039, w_eco164040, w_eco164041, w_eco164042, w_eco164043, w_eco164044, w_eco164045, w_eco164046, w_eco164047, w_eco164048, w_eco164049, w_eco164050, w_eco164051, w_eco164052, w_eco164053, w_eco164054, w_eco164055, w_eco164056, w_eco164057, w_eco164058, w_eco164059, w_eco164060, w_eco164061, w_eco164062, w_eco164063, w_eco164064, w_eco164065, w_eco164066, w_eco164067, w_eco164068, w_eco164069, w_eco164070, w_eco164071, w_eco164072, w_eco164073, w_eco164074, w_eco164075, w_eco164076, w_eco164077, w_eco164078, w_eco164079, w_eco164080, w_eco164081, w_eco164082, w_eco164083, w_eco164084, w_eco164085, w_eco164086, w_eco164087, w_eco164088, w_eco164089, w_eco164090, w_eco164091, w_eco164092, w_eco164093, w_eco164094, w_eco164095, w_eco164096, w_eco164097, w_eco164098, w_eco164099, w_eco164100, w_eco164101, w_eco164102, w_eco164103, w_eco164104, w_eco164105, w_eco164106, w_eco164107, w_eco164108, w_eco164109, w_eco164110, w_eco164111, w_eco164112, w_eco164113, w_eco164114, w_eco164115, w_eco164116, w_eco164117, w_eco164118, w_eco164119, w_eco164120, w_eco164121, w_eco164122, w_eco164123, w_eco164124, w_eco164125, w_eco164126, w_eco164127, w_eco164128, w_eco164129, w_eco164130, w_eco164131, w_eco164132, w_eco164133, w_eco164134, w_eco164135, w_eco164136, w_eco164137, w_eco164138, w_eco164139, w_eco164140, w_eco164141, w_eco164142, w_eco164143, w_eco164144, w_eco164145, w_eco164146, w_eco164147, w_eco164148, w_eco164149, w_eco164150, w_eco164151, w_eco164152, w_eco164153, w_eco164154, w_eco164155, w_eco164156, w_eco164157, w_eco164158, w_eco164159, w_eco164160, w_eco164161, w_eco164162, w_eco164163, w_eco164164, w_eco164165, w_eco164166, w_eco164167, w_eco164168, w_eco164169, w_eco164170, w_eco164171, w_eco164172, w_eco164173, w_eco164174, w_eco164175, w_eco164176, w_eco164177, w_eco164178, w_eco164179, w_eco164180, w_eco164181, w_eco164182, w_eco164183, w_eco164184, w_eco164185, w_eco164186, w_eco164187, w_eco164188, w_eco164189, w_eco164190, w_eco164191, w_eco164192, w_eco164193, w_eco164194, w_eco164195, w_eco164196, w_eco164197, w_eco164198, w_eco164199, w_eco164200, w_eco164201, w_eco164202, w_eco164203, w_eco164204, w_eco164205, w_eco164206, w_eco164207, w_eco164208, w_eco164209, w_eco164210, w_eco164211, w_eco164212, w_eco164213, w_eco164214, w_eco164215, w_eco164216, w_eco164217, w_eco164218, w_eco164219, w_eco164220, w_eco164221, w_eco164222, w_eco164223, w_eco164224, w_eco164225, w_eco164226, w_eco164227, w_eco164228, w_eco164229, w_eco164230, w_eco164231, w_eco164232, w_eco164233, w_eco164234, w_eco164235, w_eco164236, w_eco164237, w_eco164238, w_eco164239, w_eco164240, w_eco164241, w_eco164242, w_eco164243, w_eco164244, w_eco164245, w_eco164246, w_eco164247, w_eco164248, w_eco164249, w_eco164250, w_eco164251, w_eco164252, w_eco164253, w_eco164254, w_eco164255, w_eco164256, w_eco164257, w_eco164258, w_eco164259, w_eco164260, w_eco164261, w_eco164262, w_eco164263, w_eco164264, w_eco164265, w_eco164266, w_eco164267, w_eco164268, w_eco164269, w_eco164270, w_eco164271, w_eco164272, w_eco164273, w_eco164274, w_eco164275, w_eco164276, w_eco164277, w_eco164278, w_eco164279, w_eco164280, w_eco164281, w_eco164282, w_eco164283, w_eco164284, w_eco164285, w_eco164286, w_eco164287, w_eco164288, w_eco164289, w_eco164290, w_eco164291, w_eco164292, w_eco164293, w_eco164294, w_eco164295, w_eco164296, w_eco164297, w_eco164298, w_eco164299, w_eco164300, w_eco164301, w_eco164302, w_eco164303, w_eco164304, w_eco164305, w_eco164306, w_eco164307, w_eco164308, w_eco164309, w_eco164310, w_eco164311, w_eco164312, w_eco164313, w_eco164314, w_eco164315, w_eco164316, w_eco164317, w_eco164318, w_eco164319, w_eco164320, w_eco164321, w_eco164322, w_eco164323, w_eco164324, w_eco164325, w_eco164326, w_eco164327, w_eco164328, w_eco164329, w_eco164330, w_eco164331, w_eco164332, w_eco164333, w_eco164334, w_eco164335, w_eco164336, w_eco164337, w_eco164338, w_eco164339, w_eco164340, w_eco164341, w_eco164342, w_eco164343, w_eco164344, w_eco164345, w_eco164346, w_eco164347, w_eco164348, w_eco164349, w_eco164350, w_eco164351, w_eco164352, w_eco164353, w_eco164354, w_eco164355, w_eco164356, w_eco164357, w_eco164358, w_eco164359, w_eco164360, w_eco164361, w_eco164362, w_eco164363, w_eco164364, w_eco164365, w_eco164366, w_eco164367, w_eco164368, w_eco164369, w_eco164370, w_eco164371, w_eco164372, w_eco164373, w_eco164374, w_eco164375, w_eco164376, w_eco164377, w_eco164378, w_eco164379, w_eco164380, w_eco164381, w_eco164382, w_eco164383, w_eco164384, w_eco164385, w_eco164386, w_eco164387, w_eco164388, w_eco164389, w_eco164390, w_eco164391, w_eco164392, w_eco164393, w_eco164394, w_eco164395, w_eco164396, w_eco164397, w_eco164398, w_eco164399, w_eco164400, w_eco164401, w_eco164402, w_eco164403, w_eco164404, w_eco164405, w_eco164406, w_eco164407, w_eco164408, w_eco164409, w_eco164410, w_eco164411, w_eco164412, w_eco164413, w_eco164414, w_eco164415, w_eco164416, w_eco164417, w_eco164418, w_eco164419, w_eco164420, w_eco164421, w_eco164422, w_eco164423, w_eco164424, w_eco164425, w_eco164426, w_eco164427, w_eco164428, w_eco164429, w_eco164430, w_eco164431, w_eco164432, w_eco164433, w_eco164434, w_eco164435, w_eco164436, w_eco164437, w_eco164438, w_eco164439, w_eco164440, w_eco164441, w_eco164442, w_eco164443, w_eco164444, w_eco164445, w_eco164446, w_eco164447, w_eco164448, w_eco164449, w_eco164450, w_eco164451, w_eco164452, w_eco164453, w_eco164454, w_eco164455, w_eco164456, w_eco164457, w_eco164458, w_eco164459, w_eco164460, w_eco164461, w_eco164462, w_eco164463, w_eco164464, w_eco164465, w_eco164466, w_eco164467, w_eco164468, w_eco164469, w_eco164470, w_eco164471, w_eco164472, w_eco164473, w_eco164474, w_eco164475, w_eco164476, w_eco164477, w_eco164478, w_eco164479, w_eco164480, w_eco164481, w_eco164482, w_eco164483, w_eco164484, w_eco164485, w_eco164486, w_eco164487, w_eco164488, w_eco164489, w_eco164490, w_eco164491, w_eco164492, w_eco164493, w_eco164494, w_eco164495, w_eco164496, w_eco164497, w_eco164498, w_eco164499, w_eco164500, w_eco164501, w_eco164502, w_eco164503, w_eco164504, w_eco164505, w_eco164506, w_eco164507, w_eco164508, w_eco164509, w_eco164510, w_eco164511, w_eco164512, w_eco164513, w_eco164514, w_eco164515, w_eco164516, w_eco164517, w_eco164518, w_eco164519, w_eco164520, w_eco164521, w_eco164522, w_eco164523, w_eco164524, w_eco164525, w_eco164526, w_eco164527, w_eco164528, w_eco164529, w_eco164530, w_eco164531, w_eco164532, w_eco164533, w_eco164534, w_eco164535, w_eco164536, w_eco164537, w_eco164538, w_eco164539, w_eco164540, w_eco164541, w_eco164542, w_eco164543, w_eco164544, w_eco164545, w_eco164546, w_eco164547, w_eco164548, w_eco164549, w_eco164550, w_eco164551, w_eco164552, w_eco164553, w_eco164554, w_eco164555, w_eco164556, w_eco164557, w_eco164558, w_eco164559, w_eco164560, w_eco164561, w_eco164562, w_eco164563, w_eco164564, w_eco164565, w_eco164566, w_eco164567, w_eco164568, w_eco164569, w_eco164570, w_eco164571, w_eco164572, w_eco164573, w_eco164574, w_eco164575, w_eco164576, w_eco164577, w_eco164578, w_eco164579, w_eco164580, w_eco164581, w_eco164582, w_eco164583, w_eco164584, w_eco164585, w_eco164586, w_eco164587, w_eco164588, w_eco164589, w_eco164590, w_eco164591, w_eco164592, w_eco164593, w_eco164594, w_eco164595, w_eco164596, w_eco164597, w_eco164598, w_eco164599, w_eco164600, w_eco164601, w_eco164602, w_eco164603, w_eco164604, w_eco164605, w_eco164606, w_eco164607, w_eco164608, w_eco164609, w_eco164610, w_eco164611, w_eco164612, w_eco164613, w_eco164614, w_eco164615, w_eco164616, w_eco164617, w_eco164618, w_eco164619, w_eco164620, w_eco164621, w_eco164622, w_eco164623, w_eco164624, w_eco164625, w_eco164626, w_eco164627, w_eco164628, w_eco164629, w_eco164630, w_eco164631, w_eco164632, w_eco164633, w_eco164634, w_eco164635, w_eco164636, w_eco164637, w_eco164638, w_eco164639, w_eco164640, w_eco164641, w_eco164642, w_eco164643, w_eco164644, w_eco164645, w_eco164646, w_eco164647, w_eco164648, w_eco164649, w_eco164650, w_eco164651, w_eco164652, w_eco164653, w_eco164654, w_eco164655, w_eco164656, w_eco164657, w_eco164658, w_eco164659, w_eco164660, w_eco164661, w_eco164662, w_eco164663, w_eco164664, w_eco164665, w_eco164666, w_eco164667, w_eco164668, w_eco164669, w_eco164670, w_eco164671, w_eco164672, w_eco164673, w_eco164674, w_eco164675, w_eco164676, w_eco164677, w_eco164678, w_eco164679, w_eco164680, w_eco164681, w_eco164682, w_eco164683, w_eco164684, w_eco164685, w_eco164686, w_eco164687, w_eco164688, w_eco164689, w_eco164690, w_eco164691, w_eco164692, w_eco164693, w_eco164694, w_eco164695, w_eco164696, w_eco164697, w_eco164698, w_eco164699, w_eco164700, w_eco164701, w_eco164702, w_eco164703, w_eco164704, w_eco164705, w_eco164706, w_eco164707, w_eco164708, w_eco164709, w_eco164710, w_eco164711, w_eco164712, w_eco164713, w_eco164714, w_eco164715, w_eco164716, w_eco164717, w_eco164718, w_eco164719, w_eco164720, w_eco164721, w_eco164722, w_eco164723, w_eco164724, w_eco164725, w_eco164726, w_eco164727, w_eco164728, w_eco164729, w_eco164730, w_eco164731, w_eco164732, w_eco164733, w_eco164734, w_eco164735, w_eco164736, w_eco164737, w_eco164738, w_eco164739, w_eco164740, w_eco164741, w_eco164742, w_eco164743, w_eco164744, w_eco164745, w_eco164746, w_eco164747, w_eco164748, w_eco164749, w_eco164750, w_eco164751, w_eco164752, w_eco164753, w_eco164754, w_eco164755, w_eco164756, w_eco164757, w_eco164758, w_eco164759, w_eco164760, w_eco164761, w_eco164762, w_eco164763, w_eco164764, w_eco164765, w_eco164766, w_eco164767, w_eco164768, w_eco164769, w_eco164770, w_eco164771, w_eco164772, w_eco164773, w_eco164774, w_eco164775, w_eco164776, w_eco164777, w_eco164778, w_eco164779, w_eco164780, w_eco164781, w_eco164782, w_eco164783, w_eco164784, w_eco164785, w_eco164786, w_eco164787, w_eco164788, w_eco164789, w_eco164790, w_eco164791, w_eco164792, w_eco164793, w_eco164794, w_eco164795, w_eco164796, w_eco164797, w_eco164798, w_eco164799, w_eco164800, w_eco164801, w_eco164802, w_eco164803, w_eco164804, w_eco164805, w_eco164806, w_eco164807, w_eco164808, w_eco164809, w_eco164810, w_eco164811, w_eco164812, w_eco164813, w_eco164814, w_eco164815, w_eco164816, w_eco164817, w_eco164818, w_eco164819, w_eco164820, w_eco164821, w_eco164822, w_eco164823, w_eco164824, w_eco164825, w_eco164826, w_eco164827, w_eco164828, w_eco164829, w_eco164830, w_eco164831, w_eco164832, w_eco164833, w_eco164834, 