module test_8(a_gtet_b,a,b);
	input [7:0]a, b;
	output a_gtet_b;
	wire [7:0]a, b;
	wire a_gtet_b, n_8, n_13, n_43, n_52, n_59, n_64, n_67, n_149, n_156, n_158, n_171, n_403, n_407, n_410, n_415, n_425, n_432, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196;

	not g468(n_442, a[2]);
	not g469(n_443, a[1]);
	not g470(n_444, b[2]);
	not g471(n_445, b[5]);
	not g472(n_446, a[5]);
	not g473(n_447, b[7]);
	not g474(n_448, a[7]);
	not g475(n_449, a[3]);
	not g476(n_450, b[4]);
	not g477(n_451, a[4]);
	not g478(n_452, b[6]);
	not g479(n_453, a[6]);
	not g480(n_454, b[1]);
	not g481(n_455, a[0]);
	nand g482(n_8, n_449, b[3]);
	nand g47(n_52, n_8, a[2]);
	not g483(n_456, n_8);
	nand g484(n_13, a[7], n_447);
	not g485(n_457, n_13);
	nor g486(n_458, a[6], n_452);
	not g487(n_459, n_458);
	nor g488(n_407, n_442, b[2]);
	not g489(n_460, n_407);
	nor g490(n_43, n_449, b[3]);
	nor g133(n_158, n_43, a[1]);
	not g491(n_461, n_43);
	not g492(n_462, n_158);
	nor g493(n_463, n_43, n_454);
	not g494(n_464, n_463);
	nand g495(n_465, n_462, n_464);
	nand g496(n_466, n_460, n_465, b[0]);
	nor g497(n_403, a[2], n_444);
	not g498(n_467, n_403);
	nand g499(n_410, n_467, n_8, n_454);
	not g500(n_468, n_410);
	nand g501(n_469, n_460, n_461, n_443);
	nor g502(n_470, n_468, n_469);
	not g503(n_471, n_470);
	nor g504(n_472, n_456, n_461);
	not g505(n_473, n_472);
	nor g506(n_474, n_456, b[2]);
	not g507(n_475, n_474);
	nand g508(n_476, n_52, n_473, n_475);
	nor g509(n_477, n_468, n_476);
	not g510(n_478, n_477);
	nand g511(n_59, n_466, n_471, n_478);
	not g512(n_479, n_59);
	nor g513(n_480, n_59, n_451);
	not g514(n_481, n_480);
	nor g515(n_482, n_479, a[4]);
	not g516(n_483, n_482);
	nand g517(n_484, n_483, n_450);
	nand g518(n_64, n_481, n_484);
	nand g519(n_485, n_13, n_459, n_64);
	nand g520(n_67, n_448, b[7]);
	not g521(n_486, n_67);
	nor g522(n_487, n_453, b[6]);
	not g523(n_488, n_487);
	nand g524(n_489, n_67, n_488, n_446);
	nor g525(n_415, n_486, a[6]);
	not g526(n_490, n_415);
	nand g527(n_425, n_13, n_490);
	not g528(n_491, n_425);
	nor g529(n_492, n_13, n_491);
	not g530(n_493, n_492);
	nor g531(n_494, n_491, n_452);
	not g532(n_495, n_494);
	nand g533(n_496, n_489, n_493, n_495);
	nand g58(n_149, n_485, n_496);
	nor g534(n_497, a[5], n_445);
	not g535(n_498, n_497);
	nand g536(n_156, n_467, n_498);
	nor g537(n_499, n_156, n_453, n_455);
	not g538(n_500, n_499);
	nor g539(n_501, n_156, n_455, b[6]);
	not g540(n_502, n_501);
	nand g541(n_503, n_500, n_502);
	not g542(n_504, n_503);
	nor g543(n_505, a[4], n_450);
	not g544(n_506, n_505);
	nand g545(n_171, n_8, n_506);
	nor g546(n_507, n_457, n_171, n_443);
	not g547(n_508, n_507);
	nor g548(n_509, n_457, n_171, b[1]);
	not g549(n_510, n_509);
	nand g550(n_511, n_508, n_510);
	not g551(n_512, n_511);
	nor g552(n_513, n_504, n_512);
	not g553(n_514, n_513);
	nor g554(n_515, n_486, n_452, n_445);
	not g555(n_516, n_515);
	nor g556(n_517, n_490, n_445);
	not g557(n_518, n_517);
	nand g558(n_432, n_516, n_518);
	not g559(n_519, n_432);
	nor g560(n_520, n_519, a[5]);
	not g561(n_521, n_520);
	nor g562(n_522, n_519, n_64);
	not g563(n_523, n_522);
	nand g564(n_524, n_149, n_521, n_523);
	nand g565(sub_wire0, n_514, n_524);
	and _ECO_0(w_eco0, b[5], b[4], !a[4], !b[6], !a[6]);
	and _ECO_1(w_eco1, b[5], !a[5], b[4], !a[4], !b[6]);
	and _ECO_2(w_eco2, b[5], b[4], !a[4], !b[6], !a[0]);
	and _ECO_3(w_eco3, b[5], a[5], b[6], !a[6], a[0]);
	and _ECO_4(w_eco4, b[5], b[4], !a[4], !a[6], a[0]);
	and _ECO_5(w_eco5, !b[5], !a[5], !b[6], a[6], !a[0]);
	and _ECO_6(w_eco6, a[5], !b[4], a[4], b[6], !a[6], a[0]);
	and _ECO_7(w_eco7, !b[5], !b[4], a[4], b[6], !a[6], a[0]);
	and _ECO_8(w_eco8, a[2], b[2], b[5], a[3], b[4], !b[6], !a[6]);
	and _ECO_9(w_eco9, a[2], b[2], b[5], !a[5], a[3], b[4], !b[6]);
	and _ECO_10(w_eco10, a[5], !b[7], a[7], !b[6], !a[6]);
	and _ECO_11(w_eco11, !b[5], !a[5], b[7], !a[7], !b[6], !a[6]);
	and _ECO_12(w_eco12, !b[5], !b[7], a[7], !b[6], !a[6]);
	and _ECO_13(w_eco13, !a[2], b[2], b[5], b[4], !a[4], !b[6]);
	and _ECO_14(w_eco14, !a[2], b[2], !b[5], !a[5], !b[6], a[6]);
	and _ECO_15(w_eco15, a[2], b[2], b[5], !a[5], a[3], !a[4], !b[6]);
	and _ECO_16(w_eco16, a[2], b[2], b[5], a[3], b[4], !b[6], !a[0]);
	and _ECO_17(w_eco17, a[2], b[2], b[5], a[3], b[4], !a[6], a[0]);
	and _ECO_18(w_eco18, a[2], b[2], b[5], !a[5], b[4], !b[6], !b[3]);
	and _ECO_19(w_eco19, !a[2], !a[1], b[2], b[5], !a[3], b[4], !b[6]);
	and _ECO_20(w_eco20, !a[2], !a[1], b[5], !a[5], !a[3], b[4], !b[6]);
	and _ECO_21(w_eco21, b[5], !a[5], b[7], !a[7], b[4], !a[4], a[0]);
	and _ECO_22(w_eco22, a[5], !b[7], a[7], !b[6], !a[0]);
	and _ECO_23(w_eco23, a[2], !a[1], !b[2], !b[5], a[3], a[4], b[6], !a[6], a[0]);
	and _ECO_24(w_eco24, !b[5], !a[5], b[7], !a[7], !a[6], a[0]);
	and _ECO_25(w_eco25, b[5], !a[5], !b[7], a[7], !b[4], a[4], b[6], a[6], a[0]);
	and _ECO_26(w_eco26, !a[2], b[2], a[5], !b[7], a[7], !b[4], a[4], a[0]);
	and _ECO_27(w_eco27, a[2], b[2], b[5], a[3], !a[4], !b[6], !a[6]);
	and _ECO_28(w_eco28, a[2], b[2], b[5], a[3], !a[4], !a[6], a[0]);
	and _ECO_29(w_eco29, a[2], b[2], b[5], !a[5], !a[4], !b[6], !b[3]);
	and _ECO_30(w_eco30, !a[1], b[2], b[5], !a[5], !a[3], !a[4], !b[6]);
	and _ECO_31(w_eco31, !a[2], !a[1], b[5], !a[5], !a[3], !a[4], !b[6]);
	and _ECO_32(w_eco32, a[1], b[5], !a[5], b[4], !b[6], !b[0]);
	and _ECO_33(w_eco33, !a[1], b[2], b[5], !a[5], b[4], !b[6], b[3]);
	and _ECO_34(w_eco34, !a[2], !a[1], b[5], !a[5], b[4], !b[6], b[3]);
	and _ECO_35(w_eco35, a[2], b[2], b[5], b[4], !b[6], !a[6], !b[3]);
	and _ECO_36(w_eco36, a[2], b[2], b[5], b[4], !a[6], a[0], !b[3]);
	and _ECO_37(w_eco37, !a[1], b[2], b[5], !a[3], b[4], !a[6], a[0]);
	and _ECO_38(w_eco38, !a[2], !a[1], b[5], !a[3], b[4], !b[6], !a[6]);
	and _ECO_39(w_eco39, !a[2], !a[1], b[5], !a[3], b[4], !a[6], a[0]);
	and _ECO_40(w_eco40, !a[2], b[2], b[5], b[7], !a[7], b[4], !a[4], a[0]);
	and _ECO_41(w_eco41, !a[2], b[2], a[5], !b[7], a[7], !b[6]);
	and _ECO_42(w_eco42, !a[2], b[2], !b[5], !a[5], b[7], !a[7], a[0]);
	and _ECO_43(w_eco43, !a[2], b[2], !b[7], a[7], !b[4], a[4], b[6], a[6], a[0]);
	and _ECO_44(w_eco44, a[2], b[2], b[5], a[3], !a[4], !b[6], !a[0]);
	and _ECO_45(w_eco45, a[1], b[5], !a[5], !a[4], !b[6], !b[0]);
	and _ECO_46(w_eco46, a[2], !a[1], !b[2], a[5], a[3], !b[4], b[6], !a[6], a[0]);
	and _ECO_47(w_eco47, !a[1], b[2], b[5], !a[5], !a[4], !b[6], b[3]);
	and _ECO_48(w_eco48, !a[2], !a[1], b[5], !a[5], !a[4], !b[6], b[3]);
	and _ECO_49(w_eco49, a[2], b[2], b[5], !a[4], !b[6], !a[6], !b[3]);
	and _ECO_50(w_eco50, a[2], b[2], b[5], !a[4], !a[6], a[0], !b[3]);
	and _ECO_51(w_eco51, !a[2], !a[1], b[2], b[5], !a[3], !a[4], !b[6]);
	and _ECO_52(w_eco52, !a[1], b[2], b[5], !a[3], !a[4], !a[6], a[0]);
	and _ECO_53(w_eco53, !a[2], !a[1], b[5], !a[3], !a[4], !b[6], !a[6]);
	and _ECO_54(w_eco54, !a[2], !a[1], b[5], !a[3], !a[4], !a[6], a[0]);
	and _ECO_55(w_eco55, a[2], b[2], b[5], !a[5], b[7], !a[7], a[3], b[4], a[0]);
	and _ECO_56(w_eco56, a[1], b[5], b[4], !b[6], !a[6], !b[0]);
	and _ECO_57(w_eco57, a[1], b[5], b[4], !a[6], a[0], !b[0]);
	and _ECO_58(w_eco58, a[2], !b[2], a[5], a[4], b[6], !a[6], a[0], b[0]);
	and _ECO_59(w_eco59, !a[2], !a[1], b[2], b[5], b[4], !b[6], b[3]);
	and _ECO_60(w_eco60, !a[1], b[2], b[5], b[4], !a[6], a[0], b[3]);
	and _ECO_61(w_eco61, !a[2], !a[1], b[5], b[4], !b[6], !a[6], b[3]);
	and _ECO_62(w_eco62, !a[2], !a[1], b[5], b[4], !a[6], a[0], b[3]);
	and _ECO_63(w_eco63, b[2], b[5], !a[5], b[4], !b[6], b[1]);
	and _ECO_64(w_eco64, !a[1], !b[2], a[5], a[3], a[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_65(w_eco65, !a[1], b[2], b[5], b[4], !b[6], !a[0], b[3]);
	and _ECO_66(w_eco66, a[2], b[2], b[5], b[4], !b[6], !a[0], !b[3]);
	and _ECO_67(w_eco67, !a[2], !a[1], b[2], b[5], b[7], !a[7], !a[3], b[4], a[0]);
	and _ECO_68(w_eco68, !a[2], b[5], !a[5], !a[3], b[4], !b[6], b[1]);
	and _ECO_69(w_eco69, !a[2], !a[1], b[5], !a[3], b[4], !b[6], !a[0]);
	and _ECO_70(w_eco70, a[2], b[2], b[5], !a[5], b[7], !a[7], a[3], !a[4], a[0]);
	and _ECO_71(w_eco71, a[1], b[5], !a[4], !b[6], !a[6], !b[0]);
	and _ECO_72(w_eco72, a[1], b[5], !a[4], !a[6], a[0], !b[0]);
	and _ECO_73(w_eco73, a[2], !b[2], a[5], !b[4], b[6], !a[6], a[0], b[0]);
	and _ECO_74(w_eco74, a[2], !a[1], !b[2], !b[5], a[3], !b[4], b[6], !a[6], a[0]);
	and _ECO_75(w_eco75, !a[2], !a[1], b[2], b[5], !a[4], !b[6], b[3]);
	and _ECO_76(w_eco76, !a[1], b[2], b[5], !a[4], !a[6], a[0], b[3]);
	and _ECO_77(w_eco77, !a[2], !a[1], b[5], !a[4], !b[6], !a[6], b[3]);
	and _ECO_78(w_eco78, !a[2], !a[1], b[5], !a[4], !a[6], a[0], b[3]);
	and _ECO_79(w_eco79, b[2], b[5], !a[5], !a[4], !b[6], b[1]);
	and _ECO_80(w_eco80, !a[1], !b[2], a[5], a[3], !b[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_81(w_eco81, !a[1], b[2], b[5], !a[4], !b[6], !a[0], b[3]);
	and _ECO_82(w_eco82, a[2], b[2], b[5], !a[4], !b[6], !a[0], !b[3]);
	and _ECO_83(w_eco83, !a[2], !a[1], b[2], b[5], b[7], !a[7], !a[3], !a[4], a[0]);
	and _ECO_84(w_eco84, !a[2], b[5], !a[5], !a[3], !a[4], !b[6], b[1]);
	and _ECO_85(w_eco85, !a[2], !a[1], b[5], !a[3], !a[4], !b[6], !a[0]);
	and _ECO_86(w_eco86, a[1], b[5], b[4], !b[6], !a[0], !b[0]);
	and _ECO_87(w_eco87, a[2], !b[2], !b[5], a[4], b[6], !a[6], a[0], b[0]);
	and _ECO_88(w_eco88, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], a[4], b[6], a[6], a[0]);
	and _ECO_89(w_eco89, !a[2], !a[1], b[2], b[5], b[7], !a[7], b[4], a[0], b[3]);
	and _ECO_90(w_eco90, !a[2], b[5], !a[5], b[4], !b[6], b[1], b[3]);
	and _ECO_91(w_eco91, !a[2], !a[1], b[5], b[4], !b[6], !a[0], b[3]);
	and _ECO_92(w_eco92, !a[2], b[2], b[5], b[4], !b[6], b[1]);
	and _ECO_93(w_eco93, b[2], b[5], b[4], !a[6], b[1], a[0]);
	and _ECO_94(w_eco94, b[2], b[5], !a[5], b[4], !b[6], !b[0]);
	and _ECO_95(w_eco95, !b[2], a[5], a[3], a[4], b[6], !a[6], a[0], !b[3], b[0]);
	and _ECO_96(w_eco96, !a[1], !b[2], !b[5], a[3], a[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_97(w_eco97, b[5], !a[5], !a[3], b[4], !b[6], !b[1], b[3], !b[0]);
	and _ECO_98(w_eco98, a[2], b[2], b[5], !a[5], b[7], !a[7], b[4], a[0], !b[3]);
	and _ECO_99(w_eco99, a[2], !a[1], !b[2], a[5], a[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_100(w_eco100, !a[2], b[2], b[5], b[7], !a[7], b[4], b[1], a[0]);
	and _ECO_101(w_eco101, !a[2], a[1], a[5], a[4], b[6], !a[6], !b[1], a[0], b[0]);
	and _ECO_102(w_eco102, !a[2], b[5], !a[3], b[4], !b[6], !a[6], b[1]);
	and _ECO_103(w_eco103, !a[2], b[5], !a[3], b[4], !a[6], b[1], a[0]);
	and _ECO_104(w_eco104, !a[2], !a[1], b[5], !a[5], b[7], !a[7], !a[3], b[4], a[0]);
	and _ECO_105(w_eco105, a[1], b[5], !a[4], !b[6], !a[0], !b[0]);
	and _ECO_106(w_eco106, a[2], !b[2], !b[5], !b[4], b[6], !a[6], a[0], b[0]);
	and _ECO_107(w_eco107, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], !b[4], b[6], a[6], a[0]);
	and _ECO_108(w_eco108, !a[2], !a[1], b[2], b[5], b[7], !a[7], !a[4], a[0], b[3]);
	and _ECO_109(w_eco109, !a[2], b[5], !a[5], !a[4], !b[6], b[1], b[3]);
	and _ECO_110(w_eco110, !a[2], !a[1], b[5], !a[4], !b[6], !a[0], b[3]);
	and _ECO_111(w_eco111, !a[2], b[2], b[5], !a[4], !b[6], b[1]);
	and _ECO_112(w_eco112, b[2], b[5], !a[4], !a[6], b[1], a[0]);
	and _ECO_113(w_eco113, b[2], b[5], !a[5], !a[4], !b[6], !b[0]);
	and _ECO_114(w_eco114, !b[2], a[5], a[3], !b[4], b[6], !a[6], a[0], !b[3], b[0]);
	and _ECO_115(w_eco115, !a[1], !b[2], !b[5], a[3], !b[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_116(w_eco116, b[5], !a[5], !a[3], !a[4], !b[6], !b[1], b[3], !b[0]);
	and _ECO_117(w_eco117, a[2], b[2], b[5], !a[5], b[7], !a[7], !a[4], a[0], !b[3]);
	and _ECO_118(w_eco118, a[2], !a[1], !b[2], a[5], !b[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_119(w_eco119, !a[2], b[2], b[5], b[7], !a[7], !a[4], b[1], a[0]);
	and _ECO_120(w_eco120, !a[2], a[1], a[5], !b[4], b[6], !a[6], !b[1], a[0], b[0]);
	and _ECO_121(w_eco121, !a[2], b[5], !a[3], !a[4], !b[6], !a[6], b[1]);
	and _ECO_122(w_eco122, !a[2], b[5], !a[3], !a[4], !a[6], b[1], a[0]);
	and _ECO_123(w_eco123, !a[2], !a[1], b[5], !a[5], b[7], !a[7], !a[3], !a[4], a[0]);
	and _ECO_124(w_eco124, a[2], !b[2], b[5], !a[5], !b[7], a[7], a[4], b[6], a[6], a[0], b[0]);
	and _ECO_125(w_eco125, a[1], b[5], !a[5], b[7], !a[7], b[4], a[0], !b[0]);
	and _ECO_126(w_eco126, !a[2], b[5], b[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_127(w_eco127, !a[2], b[5], b[4], !a[6], b[1], a[0], b[3]);
	and _ECO_128(w_eco128, !a[2], !a[1], b[5], !a[5], b[7], !a[7], b[4], a[0], b[3]);
	and _ECO_129(w_eco129, !a[2], b[2], b[5], b[4], !b[6], !b[0]);
	and _ECO_130(w_eco130, b[2], b[5], b[4], !a[6], a[0], !b[0]);
	and _ECO_131(w_eco131, !a[2], a[5], a[3], a[4], b[6], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_132(w_eco132, !b[2], !b[5], a[3], a[4], b[6], !a[6], a[0], !b[3], b[0]);
	and _ECO_133(w_eco133, !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], a[4], b[6], a[6], a[0], !b[3]);
	and _ECO_134(w_eco134, b[2], b[5], b[4], !b[6], b[1], !a[0]);
	and _ECO_135(w_eco135, a[1], a[5], !a[3], a[4], b[6], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_136(w_eco136, !a[1], b[2], b[5], !a[5], b[7], !a[7], b[4], a[0], b[3]);
	and _ECO_137(w_eco137, b[5], !a[3], b[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_138(w_eco138, b[5], !a[3], b[4], !a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_139(w_eco139, a[2], !a[1], !b[2], a[5], a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_140(w_eco140, a[2], !a[1], !b[2], !b[5], a[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_141(w_eco141, !a[2], a[1], b[2], !b[7], a[7], a[4], b[6], a[6], !b[1], a[0], b[0]);
	and _ECO_142(w_eco142, !a[2], a[1], !b[5], a[4], b[6], !a[6], !b[1], a[0], b[0]);
	and _ECO_143(w_eco143, !a[2], b[5], !a[3], b[4], !b[6], b[1], !a[0]);
	and _ECO_144(w_eco144, a[2], !b[2], b[5], !a[5], !b[7], a[7], !b[4], b[6], a[6], a[0], b[0]);
	and _ECO_145(w_eco145, a[1], b[5], !a[5], b[7], !a[7], !a[4], a[0], !b[0]);
	and _ECO_146(w_eco146, !a[2], b[5], !a[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_147(w_eco147, !a[2], b[5], !a[4], !a[6], b[1], a[0], b[3]);
	and _ECO_148(w_eco148, !a[2], !a[1], b[5], !a[5], b[7], !a[7], !a[4], a[0], b[3]);
	and _ECO_149(w_eco149, !a[2], b[2], b[5], !a[4], !b[6], !b[0]);
	and _ECO_150(w_eco150, b[2], b[5], !a[4], !a[6], a[0], !b[0]);
	and _ECO_151(w_eco151, !a[2], a[5], a[3], !b[4], b[6], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_152(w_eco152, !b[2], !b[5], a[3], !b[4], b[6], !a[6], a[0], !b[3], b[0]);
	and _ECO_153(w_eco153, !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], !b[4], b[6], a[6], a[0], !b[3]);
	and _ECO_154(w_eco154, b[2], b[5], !a[4], !b[6], b[1], !a[0]);
	and _ECO_155(w_eco155, a[1], a[5], !a[3], !b[4], b[6], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_156(w_eco156, !a[1], b[2], b[5], !a[5], b[7], !a[7], !a[4], a[0], b[3]);
	and _ECO_157(w_eco157, b[5], !a[3], !a[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_158(w_eco158, b[5], !a[3], !a[4], !a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_159(w_eco159, a[2], !a[1], !b[2], a[5], !b[4], b[6], !a[6], b[1], a[0]);
	and _ECO_160(w_eco160, a[2], !a[1], !b[2], !b[5], !b[4], b[6], !a[6], a[0], !b[3]);
	and _ECO_161(w_eco161, !a[2], a[1], b[2], !b[7], a[7], !b[4], b[6], a[6], !b[1], a[0], b[0]);
	and _ECO_162(w_eco162, !a[2], a[1], !b[5], !b[4], b[6], !a[6], !b[1], a[0], b[0]);
	and _ECO_163(w_eco163, !a[2], b[5], !a[3], !a[4], !b[6], b[1], !a[0]);
	and _ECO_164(w_eco164, !a[2], b[5], b[4], !b[6], b[1], !a[0], b[3]);
	and _ECO_165(w_eco165, !a[2], b[2], !b[7], a[7], a[3], a[4], b[6], a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_166(w_eco166, !a[2], b[2], b[5], b[7], !a[7], b[4], a[0], !b[0]);
	and _ECO_167(w_eco167, !a[2], !b[5], a[3], a[4], b[6], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_168(w_eco168, !b[2], b[5], !a[5], !b[7], a[7], a[3], a[4], b[6], a[6], a[0], !b[3], b[0]);
	and _ECO_169(w_eco169, a[1], !b[5], !a[3], a[4], b[6], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_170(w_eco170, b[5], !a[3], b[4], !b[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_171(w_eco171, a[2], !a[1], !b[2], !b[5], a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_172(w_eco172, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[4], b[6], a[6], a[0], !b[3]);
	and _ECO_173(w_eco173, !a[2], b[5], !a[5], b[7], !a[7], !a[3], b[4], b[1], a[0]);
	and _ECO_174(w_eco174, a[1], !b[2], b[5], !a[5], !b[7], a[7], a[4], b[6], a[6], !b[1], a[0], b[0]);
	and _ECO_175(w_eco175, !a[2], b[5], !a[4], !b[6], b[1], !a[0], b[3]);
	and _ECO_176(w_eco176, !a[2], b[2], !b[7], a[7], a[3], !b[4], b[6], a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_177(w_eco177, !a[2], b[2], b[5], b[7], !a[7], !a[4], a[0], !b[0]);
	and _ECO_178(w_eco178, !a[2], !b[5], a[3], !b[4], b[6], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_179(w_eco179, !b[2], b[5], !a[5], !b[7], a[7], a[3], !b[4], b[6], a[6], a[0], !b[3], b[0]);
	and _ECO_180(w_eco180, a[1], !b[5], !a[3], !b[4], b[6], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_181(w_eco181, b[5], !a[3], !a[4], !b[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_182(w_eco182, a[2], !a[1], !b[2], !b[5], !b[4], b[6], !a[6], b[1], a[0]);
	and _ECO_183(w_eco183, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], !b[4], b[6], a[6], a[0], !b[3]);
	and _ECO_184(w_eco184, !a[2], b[5], !a[5], b[7], !a[7], !a[3], !a[4], b[1], a[0]);
	and _ECO_185(w_eco185, a[1], !b[2], b[5], !a[5], !b[7], a[7], !b[4], b[6], a[6], !b[1], a[0], b[0]);
	and _ECO_186(w_eco186, !a[2], b[5], !a[5], b[7], !a[7], b[4], b[1], a[0], b[3]);
	and _ECO_187(w_eco187, b[2], b[5], !a[5], b[7], !a[7], b[4], b[1], a[0]);
	and _ECO_188(w_eco188, a[1], b[5], !a[5], !b[7], a[7], !a[3], a[4], b[6], a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_189(w_eco189, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[4], b[6], a[6], b[1], a[0]);
	and _ECO_190(w_eco190, b[5], !a[5], b[7], !a[7], !a[3], b[4], !b[1], a[0], b[3], !b[0]);
	and _ECO_191(w_eco191, !a[2], b[5], !a[5], b[7], !a[7], !a[4], b[1], a[0], b[3]);
	and _ECO_192(w_eco192, b[2], b[5], !a[5], b[7], !a[7], !a[4], b[1], a[0]);
	and _ECO_193(w_eco193, a[1], b[5], !a[5], !b[7], a[7], !a[3], !b[4], b[6], a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_194(w_eco194, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], !b[4], b[6], a[6], b[1], a[0]);
	and _ECO_195(w_eco195, b[5], !a[5], b[7], !a[7], !a[3], !a[4], !b[1], a[0], b[3], !b[0]);
	or _ECO_196(w_eco196, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195);
	xor _ECO_out0(a_gtet_b, sub_wire0, w_eco196);

endmodule