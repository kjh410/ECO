module top(z,a,shiftCnt);
	input [31:0]a;
	input [4:0]shiftCnt;
	output [31:0]z;
	wire m21_4_mux_24_18_g32_inv_sel0, m21_4_mux_24_18_g32_w_0, m21_4_mux_24_18_g32_w_1, m21_4_mux_24_18_g31_inv_sel0, m21_4_mux_24_18_g31_w_0, m21_4_mux_24_18_g31_w_1, m21_4_mux_24_18_g30_inv_sel0, m21_4_mux_24_18_g30_w_0, m21_4_mux_24_18_g30_w_1, m21_4_mux_24_18_g29_inv_sel0, m21_4_mux_24_18_g29_w_0, m21_4_mux_24_18_g29_w_1, m21_4_mux_24_18_g28_inv_sel0, m21_4_mux_24_18_g28_w_0, m21_4_mux_24_18_g28_w_1, m21_4_mux_24_18_g27_inv_sel0, m21_4_mux_24_18_g27_w_0, m21_4_mux_24_18_g27_w_1, m21_4_mux_24_18_g26_inv_sel0, m21_4_mux_24_18_g26_w_0, m21_4_mux_24_18_g26_w_1, m21_4_mux_24_18_g25_inv_sel0, m21_4_mux_24_18_g25_w_0, m21_4_mux_24_18_g25_w_1, m21_4_mux_24_18_g24_inv_sel0, m21_4_mux_24_18_g24_w_0, m21_4_mux_24_18_g24_w_1, m21_4_mux_24_18_g23_inv_sel0, m21_4_mux_24_18_g23_w_0, m21_4_mux_24_18_g23_w_1, m21_4_mux_24_18_g22_inv_sel0, m21_4_mux_24_18_g22_w_0, m21_4_mux_24_18_g22_w_1, m21_4_mux_24_18_g21_inv_sel0, m21_4_mux_24_18_g21_w_0, m21_4_mux_24_18_g21_w_1, m21_4_mux_24_18_g20_inv_sel0, m21_4_mux_24_18_g20_w_0, m21_4_mux_24_18_g20_w_1, m21_4_mux_24_18_g19_inv_sel0, m21_4_mux_24_18_g19_w_0, m21_4_mux_24_18_g19_w_1, m21_4_mux_24_18_g18_inv_sel0, m21_4_mux_24_18_g18_w_0, m21_4_mux_24_18_g18_w_1, m21_4_mux_24_18_g17_inv_sel0, m21_4_mux_24_18_g17_w_0, m21_4_mux_24_18_g17_w_1, m21_3_mux_24_18_g9_inv_sel0, m21_3_mux_24_18_g9_w_0, m21_3_mux_24_18_g9_w_1, m21_3_mux_24_18_g32_inv_sel0, m21_3_mux_24_18_g32_w_0, m21_3_mux_24_18_g32_w_1, m21_3_mux_24_18_g31_inv_sel0, m21_3_mux_24_18_g31_w_0, m21_3_mux_24_18_g31_w_1, m21_3_mux_24_18_g30_inv_sel0, m21_3_mux_24_18_g30_w_0, m21_3_mux_24_18_g30_w_1, m21_3_mux_24_18_g29_inv_sel0, m21_3_mux_24_18_g29_w_0, m21_3_mux_24_18_g29_w_1, m21_3_mux_24_18_g28_inv_sel0, m21_3_mux_24_18_g28_w_0, m21_3_mux_24_18_g28_w_1, m21_3_mux_24_18_g27_inv_sel0, m21_3_mux_24_18_g27_w_0, m21_3_mux_24_18_g27_w_1, m21_3_mux_24_18_g26_inv_sel0, m21_3_mux_24_18_g26_w_0, m21_3_mux_24_18_g26_w_1, m21_3_mux_24_18_g25_inv_sel0, m21_3_mux_24_18_g25_w_0, m21_3_mux_24_18_g25_w_1, m21_3_mux_24_18_g24_inv_sel0, m21_3_mux_24_18_g24_w_0, m21_3_mux_24_18_g24_w_1, m21_3_mux_24_18_g23_inv_sel0, m21_3_mux_24_18_g23_w_0, m21_3_mux_24_18_g23_w_1, m21_3_mux_24_18_g22_inv_sel0, m21_3_mux_24_18_g22_w_0, m21_3_mux_24_18_g22_w_1, m21_3_mux_24_18_g21_inv_sel0, m21_3_mux_24_18_g21_w_0, m21_3_mux_24_18_g21_w_1, m21_3_mux_24_18_g20_inv_sel0, m21_3_mux_24_18_g20_w_0, m21_3_mux_24_18_g20_w_1, m21_3_mux_24_18_g19_inv_sel0, m21_3_mux_24_18_g19_w_0, m21_3_mux_24_18_g19_w_1, m21_3_mux_24_18_g18_inv_sel0, m21_3_mux_24_18_g18_w_0, m21_3_mux_24_18_g18_w_1, m21_3_mux_24_18_g17_inv_sel0, m21_3_mux_24_18_g17_w_0, m21_3_mux_24_18_g17_w_1, m21_3_mux_24_18_g16_inv_sel0, m21_3_mux_24_18_g16_w_0, m21_3_mux_24_18_g16_w_1, m21_3_mux_24_18_g15_inv_sel0, m21_3_mux_24_18_g15_w_0, m21_3_mux_24_18_g15_w_1, m21_3_mux_24_18_g14_inv_sel0, m21_3_mux_24_18_g14_w_0, m21_3_mux_24_18_g14_w_1, m21_3_mux_24_18_g13_inv_sel0, m21_3_mux_24_18_g13_w_0, m21_3_mux_24_18_g13_w_1, m21_3_mux_24_18_g12_inv_sel0, m21_3_mux_24_18_g12_w_0, m21_3_mux_24_18_g12_w_1, m21_3_mux_24_18_g11_inv_sel0, m21_3_mux_24_18_g11_w_0, m21_3_mux_24_18_g11_w_1, m21_3_mux_24_18_g10_inv_sel0, m21_3_mux_24_18_g10_w_0, m21_3_mux_24_18_g10_w_1, m21_2_mux_24_18_g9_inv_sel0, m21_2_mux_24_18_g9_w_0, m21_2_mux_24_18_g9_w_1, m21_2_mux_24_18_g8_inv_sel0, m21_2_mux_24_18_g8_w_0, m21_2_mux_24_18_g8_w_1, m21_2_mux_24_18_g7_inv_sel0, m21_2_mux_24_18_g7_w_0, m21_2_mux_24_18_g7_w_1, m21_2_mux_24_18_g6_inv_sel0, m21_2_mux_24_18_g6_w_0, m21_2_mux_24_18_g6_w_1, m21_2_mux_24_18_g32_inv_sel0, m21_2_mux_24_18_g32_w_0, m21_2_mux_24_18_g32_w_1, m21_2_mux_24_18_g31_inv_sel0, m21_2_mux_24_18_g31_w_0, m21_2_mux_24_18_g31_w_1, m21_2_mux_24_18_g30_inv_sel0, m21_2_mux_24_18_g30_w_0, m21_2_mux_24_18_g30_w_1, m21_2_mux_24_18_g29_inv_sel0, m21_2_mux_24_18_g29_w_0, m21_2_mux_24_18_g29_w_1, m21_2_mux_24_18_g28_inv_sel0, m21_2_mux_24_18_g28_w_0, m21_2_mux_24_18_g28_w_1, m21_2_mux_24_18_g27_inv_sel0, m21_2_mux_24_18_g27_w_0, m21_2_mux_24_18_g27_w_1, m21_2_mux_24_18_g26_inv_sel0, m21_2_mux_24_18_g26_w_0, m21_2_mux_24_18_g26_w_1, m21_2_mux_24_18_g25_inv_sel0, m21_2_mux_24_18_g25_w_0, m21_2_mux_24_18_g25_w_1, m21_2_mux_24_18_g24_inv_sel0, m21_2_mux_24_18_g24_w_0, m21_2_mux_24_18_g24_w_1, m21_2_mux_24_18_g23_inv_sel0, m21_2_mux_24_18_g23_w_0, m21_2_mux_24_18_g23_w_1, m21_2_mux_24_18_g22_inv_sel0, m21_2_mux_24_18_g22_w_0, m21_2_mux_24_18_g22_w_1, m21_2_mux_24_18_g21_inv_sel0, m21_2_mux_24_18_g21_w_0, m21_2_mux_24_18_g21_w_1, m21_2_mux_24_18_g20_inv_sel0, m21_2_mux_24_18_g20_w_0, m21_2_mux_24_18_g20_w_1, m21_2_mux_24_18_g19_inv_sel0, m21_2_mux_24_18_g19_w_0, m21_2_mux_24_18_g19_w_1, m21_2_mux_24_18_g18_inv_sel0, m21_2_mux_24_18_g18_w_0, m21_2_mux_24_18_g18_w_1, m21_2_mux_24_18_g17_inv_sel0, m21_2_mux_24_18_g17_w_0, m21_2_mux_24_18_g17_w_1, m21_2_mux_24_18_g16_inv_sel0, m21_2_mux_24_18_g16_w_0, m21_2_mux_24_18_g16_w_1, m21_2_mux_24_18_g15_inv_sel0, m21_2_mux_24_18_g15_w_0, m21_2_mux_24_18_g15_w_1, m21_2_mux_24_18_g14_inv_sel0, m21_2_mux_24_18_g14_w_0, m21_2_mux_24_18_g14_w_1, m21_2_mux_24_18_g13_inv_sel0, m21_2_mux_24_18_g13_w_0, m21_2_mux_24_18_g13_w_1, m21_2_mux_24_18_g12_inv_sel0, m21_2_mux_24_18_g12_w_0, m21_2_mux_24_18_g12_w_1, m21_2_mux_24_18_g11_inv_sel0, m21_2_mux_24_18_g11_w_0, m21_2_mux_24_18_g11_w_1, m21_2_mux_24_18_g10_inv_sel0, m21_2_mux_24_18_g10_w_0, m21_2_mux_24_18_g10_w_1, m21_1_mux_24_18_g9_inv_sel0, m21_1_mux_24_18_g9_w_0, m21_1_mux_24_18_g9_w_1, m21_1_mux_24_18_g8_inv_sel0, m21_1_mux_24_18_g8_w_0, m21_1_mux_24_18_g8_w_1, m21_1_mux_24_18_g7_inv_sel0, m21_1_mux_24_18_g7_w_0, m21_1_mux_24_18_g7_w_1, m21_1_mux_24_18_g6_inv_sel0, m21_1_mux_24_18_g6_w_0, m21_1_mux_24_18_g6_w_1, m21_1_mux_24_18_g5_inv_sel0, m21_1_mux_24_18_g5_w_0, m21_1_mux_24_18_g5_w_1, m21_1_mux_24_18_g4_inv_sel0, m21_1_mux_24_18_g4_w_0, m21_1_mux_24_18_g4_w_1, m21_1_mux_24_18_g32_inv_sel0, m21_1_mux_24_18_g32_w_0, m21_1_mux_24_18_g32_w_1, m21_1_mux_24_18_g31_inv_sel0, m21_1_mux_24_18_g31_w_0, m21_1_mux_24_18_g31_w_1, m21_1_mux_24_18_g30_inv_sel0, m21_1_mux_24_18_g30_w_0, m21_1_mux_24_18_g30_w_1, m21_1_mux_24_18_g3_inv_sel0, m21_1_mux_24_18_g3_w_0, m21_1_mux_24_18_g3_w_1, m21_1_mux_24_18_g29_inv_sel0, m21_1_mux_24_18_g29_w_0, m21_1_mux_24_18_g29_w_1, m21_1_mux_24_18_g28_inv_sel0, m21_1_mux_24_18_g28_w_0, m21_1_mux_24_18_g28_w_1, m21_1_mux_24_18_g27_inv_sel0, m21_1_mux_24_18_g27_w_0, m21_1_mux_24_18_g27_w_1, m21_1_mux_24_18_g26_inv_sel0, m21_1_mux_24_18_g26_w_0, m21_1_mux_24_18_g26_w_1, m21_1_mux_24_18_g25_inv_sel0, m21_1_mux_24_18_g25_w_0, m21_1_mux_24_18_g25_w_1, m21_1_mux_24_18_g24_inv_sel0, m21_1_mux_24_18_g24_w_0, m21_1_mux_24_18_g24_w_1, m21_1_mux_24_18_g23_inv_sel0, m21_1_mux_24_18_g23_w_0, m21_1_mux_24_18_g23_w_1, m21_1_mux_24_18_g22_inv_sel0, m21_1_mux_24_18_g22_w_0, m21_1_mux_24_18_g22_w_1, m21_1_mux_24_18_g21_inv_sel0, m21_1_mux_24_18_g21_w_0, m21_1_mux_24_18_g21_w_1, m21_1_mux_24_18_g20_inv_sel0, m21_1_mux_24_18_g20_w_0, m21_1_mux_24_18_g20_w_1, m21_1_mux_24_18_g2_inv_sel0, m21_1_mux_24_18_g2_w_0, m21_1_mux_24_18_g2_w_1, m21_1_mux_24_18_g19_inv_sel0, m21_1_mux_24_18_g19_w_0, m21_1_mux_24_18_g19_w_1, m21_1_mux_24_18_g18_inv_sel0, m21_1_mux_24_18_g18_w_0, m21_1_mux_24_18_g18_w_1, m21_1_mux_24_18_g17_inv_sel0, m21_1_mux_24_18_g17_w_0, m21_1_mux_24_18_g17_w_1, m21_1_mux_24_18_g16_inv_sel0, m21_1_mux_24_18_g16_w_0, m21_1_mux_24_18_g16_w_1, m21_1_mux_24_18_g15_inv_sel0, m21_1_mux_24_18_g15_w_0, m21_1_mux_24_18_g15_w_1, m21_1_mux_24_18_g14_inv_sel0, m21_1_mux_24_18_g14_w_0, m21_1_mux_24_18_g14_w_1, m21_1_mux_24_18_g13_inv_sel0, m21_1_mux_24_18_g13_w_0, m21_1_mux_24_18_g13_w_1, m21_1_mux_24_18_g12_inv_sel0, m21_1_mux_24_18_g12_w_0, m21_1_mux_24_18_g12_w_1, m21_1_mux_24_18_g11_inv_sel0, m21_1_mux_24_18_g11_w_0, m21_1_mux_24_18_g11_w_1, m21_1_mux_24_18_g10_inv_sel0, m21_1_mux_24_18_g10_w_0, m21_1_mux_24_18_g10_w_1, m21_0_mux_24_18_g9_inv_sel0, m21_0_mux_24_18_g9_w_0, m21_0_mux_24_18_g9_w_1, m21_0_mux_24_18_g8_inv_sel0, m21_0_mux_24_18_g8_w_0, m21_0_mux_24_18_g8_w_1, m21_0_mux_24_18_g7_inv_sel0, m21_0_mux_24_18_g7_w_0, m21_0_mux_24_18_g7_w_1, m21_0_mux_24_18_g6_inv_sel0, m21_0_mux_24_18_g6_w_0, m21_0_mux_24_18_g6_w_1, m21_0_mux_24_18_g5_inv_sel0, m21_0_mux_24_18_g5_w_0, m21_0_mux_24_18_g5_w_1, m21_0_mux_24_18_g4_inv_sel0, m21_0_mux_24_18_g4_w_0, m21_0_mux_24_18_g4_w_1, m21_0_mux_24_18_g32_inv_sel0, m21_0_mux_24_18_g32_w_0, m21_0_mux_24_18_g32_w_1, m21_0_mux_24_18_g31_inv_sel0, m21_0_mux_24_18_g31_w_0, m21_0_mux_24_18_g31_w_1, m21_0_mux_24_18_g30_inv_sel0, m21_0_mux_24_18_g30_w_0, m21_0_mux_24_18_g30_w_1, m21_0_mux_24_18_g3_inv_sel0, m21_0_mux_24_18_g3_w_0, m21_0_mux_24_18_g3_w_1, m21_0_mux_24_18_g29_inv_sel0, m21_0_mux_24_18_g29_w_0, m21_0_mux_24_18_g29_w_1, m21_0_mux_24_18_g28_inv_sel0, m21_0_mux_24_18_g28_w_0, m21_0_mux_24_18_g28_w_1, m21_0_mux_24_18_g27_inv_sel0, m21_0_mux_24_18_g27_w_0, m21_0_mux_24_18_g27_w_1, m21_0_mux_24_18_g26_inv_sel0, m21_0_mux_24_18_g26_w_0, m21_0_mux_24_18_g26_w_1, m21_0_mux_24_18_g25_inv_sel0, m21_0_mux_24_18_g25_w_0, m21_0_mux_24_18_g25_w_1, m21_0_mux_24_18_g24_inv_sel0, m21_0_mux_24_18_g24_w_0, m21_0_mux_24_18_g24_w_1, m21_0_mux_24_18_g23_inv_sel0, m21_0_mux_24_18_g23_w_0, m21_0_mux_24_18_g23_w_1, m21_0_mux_24_18_g22_inv_sel0, m21_0_mux_24_18_g22_w_0, m21_0_mux_24_18_g22_w_1, m21_0_mux_24_18_g21_inv_sel0, m21_0_mux_24_18_g21_w_0, m21_0_mux_24_18_g21_w_1, m21_0_mux_24_18_g20_inv_sel0, m21_0_mux_24_18_g20_w_0, m21_0_mux_24_18_g20_w_1, m21_0_mux_24_18_g2_inv_sel0, m21_0_mux_24_18_g2_w_0, m21_0_mux_24_18_g2_w_1, m21_0_mux_24_18_g19_inv_sel0, m21_0_mux_24_18_g19_w_0, m21_0_mux_24_18_g19_w_1, m21_0_mux_24_18_g18_inv_sel0, m21_0_mux_24_18_g18_w_0, m21_0_mux_24_18_g18_w_1, m21_0_mux_24_18_g17_inv_sel0, m21_0_mux_24_18_g17_w_0, m21_0_mux_24_18_g17_w_1, m21_0_mux_24_18_g16_inv_sel0, m21_0_mux_24_18_g16_w_0, m21_0_mux_24_18_g16_w_1, m21_0_mux_24_18_g15_inv_sel0, m21_0_mux_24_18_g15_w_0, m21_0_mux_24_18_g15_w_1, m21_0_mux_24_18_g14_inv_sel0, m21_0_mux_24_18_g14_w_0, m21_0_mux_24_18_g14_w_1, m21_0_mux_24_18_g13_inv_sel0, m21_0_mux_24_18_g13_w_0, m21_0_mux_24_18_g13_w_1, m21_0_mux_24_18_g12_inv_sel0, m21_0_mux_24_18_g12_w_0, m21_0_mux_24_18_g12_w_1, m21_0_mux_24_18_g11_inv_sel0, m21_0_mux_24_18_g11_w_0, m21_0_mux_24_18_g11_w_1, m21_0_mux_24_18_g10_inv_sel0, m21_0_mux_24_18_g10_w_0, m21_0_mux_24_18_g10_w_1, n_247, n_246, n_243, n_242, n_239, n_238, n_235, n_234, n_231, n_230, n_227, n_226, n_223, n_222, n_219, n_218, n_215, n_214, n_211, n_210, n_207, n_206, n_203, n_202, n_199, n_198, n_195, n_194, n_191, n_190, n_187, n_186, n_185, n_184, n_183, n_182, n_179, n_178, n_175, n_174, n_171, n_170, n_167, n_166, n_163, n_162, n_159, n_158, n_155, n_154, n_153, n_152, n_151, n_150, n_147, n_146, n_143, n_142, n_139, n_138, n_135, n_134, n_133, n_132, m21_4_n_81, m21_4_n_80, m21_4_n_79, m21_4_n_78, m21_4_n_77, m21_4_n_76, m21_4_n_75, m21_4_n_74, m21_4_n_73, m21_4_n_72, m21_4_n_71, m21_4_n_70, m21_4_n_69, m21_4_n_68, m21_4_n_67, m21_4_n_66, m21_3_n_89, m21_3_n_88, m21_3_n_87, m21_3_n_86, m21_3_n_85, m21_3_n_84, m21_3_n_83, m21_3_n_82, m21_3_n_81, m21_3_n_80, m21_3_n_79, m21_3_n_78, m21_3_n_77, m21_3_n_76, m21_3_n_75, m21_3_n_74, m21_3_n_73, m21_3_n_72, m21_3_n_71, m21_3_n_70, m21_3_n_69, m21_3_n_68, m21_3_n_67, m21_3_n_66, m21_2_n_92, m21_2_n_91, m21_2_n_90, m21_2_n_89, m21_2_n_88, m21_2_n_87, m21_2_n_86, m21_2_n_85, m21_2_n_84, m21_2_n_83, m21_2_n_82, m21_2_n_81, m21_2_n_80, m21_2_n_79, m21_2_n_78, m21_2_n_77, m21_2_n_76, m21_2_n_75, m21_2_n_74, m21_2_n_73, m21_2_n_72, m21_2_n_71, m21_2_n_70, m21_2_n_69, m21_2_n_68, m21_2_n_67, m21_2_n_66, m21_1_n_96, m21_1_n_95, m21_1_n_94, m21_1_n_93, m21_1_n_92, m21_1_n_91, m21_1_n_90, m21_1_n_89, m21_1_n_88, m21_1_n_87, m21_1_n_86, m21_1_n_85, m21_1_n_84, m21_1_n_83, m21_1_n_82, m21_1_n_81, m21_1_n_80, m21_1_n_79, m21_1_n_78, m21_1_n_77, m21_1_n_76, m21_1_n_75, m21_1_n_74, m21_1_n_73, m21_1_n_72, m21_1_n_71, m21_1_n_70, m21_1_n_69, m21_1_n_68, m21_1_n_67, m21_1_n_66, m21_0_n_96, m21_0_n_95, m21_0_n_94, m21_0_n_93, m21_0_n_92, m21_0_n_91, m21_0_n_90, m21_0_n_89, m21_0_n_88, m21_0_n_87, m21_0_n_86, m21_0_n_85, m21_0_n_84, m21_0_n_83, m21_0_n_82, m21_0_n_81, m21_0_n_80, m21_0_n_79, m21_0_n_78, m21_0_n_77, m21_0_n_76, m21_0_n_75, m21_0_n_74, m21_0_n_73, m21_0_n_72, m21_0_n_71, m21_0_n_70, m21_0_n_69, m21_0_n_68, m21_0_n_67, m21_0_n_66;
	wire [31:0]d3, d2, d1, d0, notA, z;
	wire [4:0]shiftCnt;
	wire [31:0]a;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, sub_wire1, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, sub_wire2, w_eco9, sub_wire3, w_eco10, sub_wire4, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, sub_wire5, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, sub_wire6, w_eco21, sub_wire7, w_eco22, sub_wire8, w_eco23, w_eco24, w_eco25, w_eco26, sub_wire9, w_eco27, w_eco28, w_eco29, w_eco30, sub_wire10, w_eco31, w_eco32, w_eco33, sub_wire11, w_eco34, w_eco35, w_eco36, w_eco37, sub_wire12, w_eco38, w_eco39, w_eco40, sub_wire13, w_eco41, w_eco42, w_eco43, w_eco44, sub_wire14, w_eco45, w_eco46, w_eco47, w_eco48, sub_wire15, w_eco49, w_eco50, w_eco51, sub_wire16, w_eco52, w_eco53, w_eco54, sub_wire17, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, sub_wire18, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, sub_wire19, w_eco65, sub_wire20, w_eco66, sub_wire21, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, sub_wire22, w_eco72, w_eco73, w_eco74, sub_wire23, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, sub_wire24, w_eco80, sub_wire25, w_eco81, sub_wire26, w_eco82, w_eco83, w_eco84, sub_wire27, w_eco85, w_eco86, w_eco87, w_eco88, sub_wire28, w_eco89, w_eco90, w_eco91, w_eco92, sub_wire29, w_eco93, w_eco94, w_eco95, sub_wire30, w_eco96, w_eco97, w_eco98, sub_wire31, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103;

	and _ECO_1(w_eco1, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_2(w_eco2, !shiftCnt[3], shiftCnt[2]);
	or _ECO_3(w_eco3, w_eco0, w_eco1, w_eco2);
	xor _ECO_out0(z[31], sub_wire0, w_eco3);
	assign w_eco4 = !shiftCnt[1];
	assign w_eco5 = shiftCnt[4];
	assign w_eco6 = shiftCnt[2];
	assign w_eco7 = !shiftCnt[3];
	or _ECO_8(w_eco8, w_eco4, w_eco5, w_eco6, w_eco7);
	xor _ECO_out1(z[22], sub_wire1, w_eco8);
	assign w_eco9 = 1'b1;
	xor _ECO_out2(z[21], sub_wire2, w_eco9);
	assign w_eco10 = 1'b1;
	xor _ECO_out3(z[20], sub_wire3, w_eco10);
	assign w_eco11 = !shiftCnt[1];
	assign w_eco12 = shiftCnt[4];
	assign w_eco13 = !shiftCnt[2];
	assign w_eco14 = !shiftCnt[3];
	or _ECO_15(w_eco15, w_eco11, w_eco12, w_eco13, w_eco14);
	xor _ECO_out4(z[19], sub_wire4, w_eco15);
	assign w_eco16 = !shiftCnt[1];
	assign w_eco17 = shiftCnt[4];
	assign w_eco18 = !shiftCnt[2];
	assign w_eco19 = !shiftCnt[3];
	or _ECO_20(w_eco20, w_eco16, w_eco17, w_eco18, w_eco19);
	xor _ECO_out5(z[18], sub_wire5, w_eco20);
	assign w_eco21 = 1'b1;
	xor _ECO_out6(z[17], sub_wire6, w_eco21);
	assign w_eco22 = 1'b1;
	xor _ECO_out7(z[16], sub_wire7, w_eco22);
	assign w_eco23 = !shiftCnt[4];
	and _ECO_24(w_eco24, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_25(w_eco25, !shiftCnt[3], shiftCnt[2]);
	or _ECO_26(w_eco26, w_eco23, w_eco24, w_eco25);
	xor _ECO_out8(z[15], sub_wire8, w_eco26);
	assign w_eco27 = !shiftCnt[4];
	and _ECO_28(w_eco28, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_29(w_eco29, !shiftCnt[3], shiftCnt[2]);
	or _ECO_30(w_eco30, w_eco27, w_eco28, w_eco29);
	xor _ECO_out9(z[14], sub_wire9, w_eco30);
	assign w_eco31 = !shiftCnt[4];
	assign w_eco32 = !shiftCnt[3];
	or _ECO_33(w_eco33, w_eco31, w_eco32);
	xor _ECO_out10(z[13], sub_wire10, w_eco33);
	assign w_eco34 = shiftCnt[4];
	and _ECO_35(w_eco35, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_36(w_eco36, !shiftCnt[3], shiftCnt[2]);
	or _ECO_37(w_eco37, w_eco34, w_eco35, w_eco36);
	xor _ECO_out11(z[30], sub_wire11, w_eco37);
	assign w_eco38 = !shiftCnt[4];
	assign w_eco39 = !shiftCnt[3];
	or _ECO_40(w_eco40, w_eco38, w_eco39);
	xor _ECO_out12(z[12], sub_wire12, w_eco40);
	assign w_eco41 = !shiftCnt[4];
	and _ECO_42(w_eco42, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_43(w_eco43, !shiftCnt[3], !shiftCnt[2]);
	or _ECO_44(w_eco44, w_eco41, w_eco42, w_eco43);
	xor _ECO_out13(z[11], sub_wire13, w_eco44);
	assign w_eco45 = !shiftCnt[4];
	and _ECO_46(w_eco46, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_47(w_eco47, !shiftCnt[3], !shiftCnt[2]);
	or _ECO_48(w_eco48, w_eco45, w_eco46, w_eco47);
	xor _ECO_out14(z[10], sub_wire14, w_eco48);
	assign w_eco49 = !shiftCnt[4];
	assign w_eco50 = !shiftCnt[3];
	or _ECO_51(w_eco51, w_eco49, w_eco50);
	xor _ECO_out15(z[9], sub_wire15, w_eco51);
	assign w_eco52 = !shiftCnt[4];
	assign w_eco53 = !shiftCnt[3];
	or _ECO_54(w_eco54, w_eco52, w_eco53);
	xor _ECO_out16(z[8], sub_wire16, w_eco54);
	assign w_eco55 = !shiftCnt[1];
	assign w_eco56 = !shiftCnt[4];
	assign w_eco57 = shiftCnt[2];
	assign w_eco58 = !shiftCnt[3];
	or _ECO_59(w_eco59, w_eco55, w_eco56, w_eco57, w_eco58);
	xor _ECO_out17(z[7], sub_wire17, w_eco59);
	assign w_eco60 = !shiftCnt[1];
	assign w_eco61 = !shiftCnt[4];
	assign w_eco62 = shiftCnt[2];
	assign w_eco63 = !shiftCnt[3];
	or _ECO_64(w_eco64, w_eco60, w_eco61, w_eco62, w_eco63);
	xor _ECO_out18(z[6], sub_wire18, w_eco64);
	assign w_eco65 = 1'b1;
	xor _ECO_out19(z[5], sub_wire19, w_eco65);
	assign w_eco66 = 1'b1;
	xor _ECO_out20(z[4], sub_wire20, w_eco66);
	assign w_eco67 = !shiftCnt[1];
	assign w_eco68 = !shiftCnt[4];
	assign w_eco69 = !shiftCnt[2];
	assign w_eco70 = !shiftCnt[3];
	or _ECO_71(w_eco71, w_eco67, w_eco68, w_eco69, w_eco70);
	xor _ECO_out21(z[3], sub_wire21, w_eco71);
	assign w_eco72 = shiftCnt[4];
	assign w_eco73 = !shiftCnt[3];
	or _ECO_74(w_eco74, w_eco72, w_eco73);
	xor _ECO_out22(z[29], sub_wire22, w_eco74);
	assign w_eco75 = !shiftCnt[1];
	assign w_eco76 = !shiftCnt[4];
	assign w_eco77 = !shiftCnt[2];
	assign w_eco78 = !shiftCnt[3];
	or _ECO_79(w_eco79, w_eco75, w_eco76, w_eco77, w_eco78);
	xor _ECO_out23(z[2], sub_wire23, w_eco79);
	assign w_eco80 = 1'b1;
	xor _ECO_out24(z[1], sub_wire24, w_eco80);
	assign w_eco81 = 1'b1;
	xor _ECO_out25(z[0], sub_wire25, w_eco81);
	assign w_eco82 = shiftCnt[4];
	assign w_eco83 = !shiftCnt[3];
	or _ECO_84(w_eco84, w_eco82, w_eco83);
	xor _ECO_out26(z[28], sub_wire26, w_eco84);
	assign w_eco85 = shiftCnt[4];
	and _ECO_86(w_eco86, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_87(w_eco87, !shiftCnt[3], !shiftCnt[2]);
	or _ECO_88(w_eco88, w_eco85, w_eco86, w_eco87);
	xor _ECO_out27(z[27], sub_wire27, w_eco88);
	assign w_eco89 = shiftCnt[4];
	and _ECO_90(w_eco90, !shiftCnt[3], !shiftCnt[1]);
	and _ECO_91(w_eco91, !shiftCnt[3], !shiftCnt[2]);
	or _ECO_92(w_eco92, w_eco89, w_eco90, w_eco91);
	xor _ECO_out28(z[26], sub_wire28, w_eco92);
	assign w_eco93 = shiftCnt[4];
	assign w_eco94 = !shiftCnt[3];
	or _ECO_95(w_eco95, w_eco93, w_eco94);
	xor _ECO_out29(z[25], sub_wire29, w_eco95);
	assign w_eco96 = shiftCnt[4];
	assign w_eco97 = !shiftCnt[3];
	or _ECO_98(w_eco98, w_eco96, w_eco97);
	xor _ECO_out30(z[24], sub_wire30, w_eco98);
	assign w_eco99 = !shiftCnt[1];
	assign w_eco100 = shiftCnt[4];
	assign w_eco101 = shiftCnt[2];
	assign w_eco102 = !shiftCnt[3];
	or _ECO_103(w_eco103, w_eco99, w_eco100, w_eco101, w_eco102);
	xor _ECO_out31(z[23], sub_wire31, w_eco103);

endmodule