module top(prim_out,sel_prim);
	input [18:0]sel_prim;
	output [31:0]prim_out;
	wire [18:0]sel_prim;
	wire [31:0]prim_out;
	wire ctl_sel_prim_412_12_n_205, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_411, ctl_sel_prim_412_12_n_442, ctl_sel_prim_412_12_n_467, ctl_sel_prim_412_12_n_493, ctl_sel_prim_412_12_n_538, n_663, n_678, n_700, n_707, n_717, n_725, n_749, n_855, n_856, n_863, n_864, n_865, n_866, n_867, n_868, n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_883, n_884, n_886, n_889, n_890, n_893, n_894, n_895, n_898, n_901, n_905, n_912, n_913, n_918, n_919, n_1234, n_1256, n_1259, n_1260, n_1261, n_1262, n_1263, n_1264, n_1265, n_1266, n_1267, n_1268, n_1269, n_1270, n_1271, n_1272, n_1273, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280, n_1281, n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1288, n_1289, n_1290, n_1291, n_1292, n_1293, n_1294, n_1295, n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316, n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325, n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349, n_1350, n_1351;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, sub_wire1, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, sub_wire2, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, sub_wire3, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, sub_wire4, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, sub_wire5, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, sub_wire6, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, sub_wire7, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, sub_wire8, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, sub_wire9, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, sub_wire10, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, sub_wire11, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, sub_wire12, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, sub_wire13, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, sub_wire14, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, sub_wire15, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, sub_wire16, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, sub_wire17, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, sub_wire18, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, sub_wire19, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, sub_wire20, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, sub_wire21, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, sub_wire22, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634, sub_wire23, w_eco1635, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, sub_wire24, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, sub_wire25, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, sub_wire26, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914;

	assign prim_out[0] = 0;
	assign prim_out[2] = prim_out[5];
	assign prim_out[3] = 1;
	assign prim_out[4] = prim_out[5];
	assign sub_wire0 = prim_out[12];
	assign sub_wire2 = prim_out[11];
	assign sub_wire4 = prim_out[12];
	assign sub_wire5 = prim_out[25];
	assign sub_wire7 = prim_out[26];
	assign sub_wire9 = prim_out[27];
	assign sub_wire11 = prim_out[30];
	assign sub_wire13 = prim_out[31];
	not ctl_sel_prim_412_12_g171(sub_wire15, prim_out[5]);
	nor ctl_sel_prim_412_12_g150(ctl_sel_prim_412_12_n_493, n_1277, ctl_sel_prim_412_12_n_411, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_205);
	nand ctl_sel_prim_412_12_g177(ctl_sel_prim_412_12_n_538, n_1284, n_1291, n_883, n_884);
	nor ctl_sel_prim_412_12_g134(ctl_sel_prim_412_12_n_442, n_1309, ctl_sel_prim_412_12_n_411, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_205);
	nor ctl_sel_prim_412_12_g142(ctl_sel_prim_412_12_n_467, n_1310, ctl_sel_prim_412_12_n_411, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_205);
	nand g424(n_886, n_855, n_856, n_873, n_874);
	nand g427(n_889, n_867, n_868, n_869, n_875);
	nand g428(n_890, n_870, n_871, n_872, n_876);
	nand g429(n_678, prim_out[5], n_863);
	nand g431(n_893, n_855, n_864, n_873, n_874);
	nand g432(n_894, n_865, n_866, n_867, n_868);
	nand g433(n_895, n_869, n_871, n_872, n_875);
	nand g436(n_898, n_864, n_865, n_870, n_875);
	nand g439(n_901, n_863, n_866, n_869, n_870);
	nand g443(n_905, n_855, n_865, n_868, n_869);
	nand g450(n_912, n_863, n_864, n_865, n_866);
	nand g451(n_913, n_855, n_863, n_864, n_865);
	nand g456(n_918, n_855, n_856, n_865, n_874);
	nand g457(n_919, n_868, n_869, n_871, n_876);
	not g687(sub_wire16, n_678);
	not g688(sub_wire6, n_700);
	not g689(sub_wire17, n_707);
	not g691(sub_wire18, n_725);
	not g692(sub_wire12, n_663);
	not g694(sub_wire19, n_749);
	not g695(sub_wire20, n_717);
	not g961(n_1259, sel_prim[0]);
	not g962(n_1260, sel_prim[1]);
	not g963(n_1261, sel_prim[2]);
	not g964(n_1262, sel_prim[15]);
	not g965(n_1263, sel_prim[16]);
	not g966(n_1264, sel_prim[11]);
	not g967(n_1265, sel_prim[12]);
	not g968(n_1266, sel_prim[13]);
	not g969(n_1267, sel_prim[14]);
	not g970(n_1268, sel_prim[7]);
	not g971(n_1269, sel_prim[8]);
	not g972(n_1270, sel_prim[9]);
	not g973(n_1271, sel_prim[10]);
	not g974(n_1272, sel_prim[3]);
	not g975(n_1273, sel_prim[4]);
	not g976(n_1274, sel_prim[5]);
	not g977(n_1275, sel_prim[6]);
	not g978(n_1276, sel_prim[17]);
	nand g979(n_1277, sel_prim[18], n_1276, n_1263, n_1262);
	nand g980(ctl_sel_prim_412_12_n_411, n_1267, n_1266, n_1265, n_1264);
	nand g981(ctl_sel_prim_412_12_n_308, n_1271, n_1270, n_1269, n_1268);
	not g982(n_1278, ctl_sel_prim_412_12_n_308);
	nand g983(ctl_sel_prim_412_12_n_205, n_1275, n_1274, n_1273, n_1272);
	not g984(n_1279, ctl_sel_prim_412_12_n_205);
	nand g985(n_1234, n_1261, n_1260, n_1259);
	not g986(n_1280, n_1234);
	nand g987(prim_out[5], ctl_sel_prim_412_12_n_493, n_1280);
	nand g988(n_855, sel_prim[1], n_1259);
	not g989(n_1281, n_855);
	nand g990(n_856, sel_prim[2], n_1260, n_1259);
	not g991(n_1282, n_856);
	nand g992(n_873, n_1280, sel_prim[3]);
	not g993(n_1283, n_873);
	nor g994(n_1284, n_1281, n_1282, n_1283, sel_prim[0]);
	nand g995(n_874, n_1280, sel_prim[4], n_1272);
	not g996(n_1285, n_874);
	nand g997(n_865, n_1280, n_1279, sel_prim[7]);
	not g998(n_1286, n_865);
	nand g999(n_863, n_1280, sel_prim[5], n_1273, n_1272);
	not g1000(n_1287, n_863);
	nand g1001(n_1288, sel_prim[6], n_1274, n_1273, n_1272);
	not g1002(n_1289, n_1288);
	nand g1003(n_864, n_1280, n_1289);
	not g1004(n_1290, n_864);
	nor g1005(n_1291, n_1285, n_1286, n_1287, n_1290);
	nand g1006(n_875, n_1280, n_1278, n_1279, sel_prim[11]);
	not g1007(n_1292, n_875);
	nand g1008(n_1293, sel_prim[10], n_1270, n_1269, n_1268);
	not g1009(n_1294, n_1293);
	nand g1010(n_868, n_1280, n_1279, n_1294);
	not g1011(n_1295, n_868);
	nand g1012(n_866, n_1280, n_1279, sel_prim[8], n_1268);
	not g1013(n_1296, n_866);
	nor g1014(n_1297, ctl_sel_prim_412_12_n_205, n_1270, sel_prim[8], sel_prim[7]);
	nand g1015(n_867, n_1280, n_1297);
	not g1016(n_1298, n_867);
	nor g1017(n_883, n_1292, n_1295, n_1296, n_1298);
	nor g1018(n_1299, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_205, n_1265, sel_prim[11]);
	nand g1019(n_869, n_1280, n_1299);
	not g1020(n_1300, n_869);
	nand g1021(n_1301, sel_prim[14], n_1266, n_1265, n_1264);
	not g1022(n_1302, n_1301);
	nand g1023(n_871, n_1280, n_1278, n_1279, n_1302);
	not g1024(n_1303, n_871);
	nor g1025(n_1304, ctl_sel_prim_412_12_n_411, ctl_sel_prim_412_12_n_308, ctl_sel_prim_412_12_n_205, n_1262);
	nand g1026(n_872, n_1280, n_1304);
	not g1027(n_1305, n_872);
	nand g1028(n_1306, sel_prim[13], n_1265, n_1264);
	not g1029(n_1307, n_1306);
	nand g1030(n_870, n_1280, n_1278, n_1279, n_1307);
	not g1031(n_1308, n_870);
	nor g1032(n_884, n_1300, n_1303, n_1305, n_1308);
	nand g1033(n_1309, sel_prim[16], n_1262);
	nand g1034(n_1310, sel_prim[17], n_1263, n_1262);
	not g1035(n_1311, n_886);
	not g1036(n_1312, n_889);
	nand g1037(n_876, ctl_sel_prim_412_12_n_442, n_1280);
	not g1038(n_1313, n_876);
	not g1039(n_1314, n_890);
	not g1040(n_1315, n_893);
	not g1041(n_1316, n_894);
	not g1042(n_1317, n_895);
	not g1043(n_1318, n_898);
	not g1044(n_1319, n_901);
	not g1045(n_1320, n_905);
	not g1046(n_1321, n_912);
	not g1047(n_1322, n_913);
	not g1048(n_1323, n_918);
	not g1049(n_1324, n_919);
	nand g1050(n_877, ctl_sel_prim_412_12_n_467, n_1280);
	not g1051(n_1325, n_877);
	nand g1052(sub_wire14, n_1311, n_876, n_877, n_875);
	nand g1053(n_1326, n_1311, n_1318, n_876, n_872);
	not g1054(n_1327, n_1326);
	nand g1055(n_700, n_877, n_1327);
	nand g1056(n_707, n_1319, prim_out[5]);
	nand g1057(sub_wire21, n_1320, n_877, n_872);
	nand g1058(n_1328, n_869, n_863, n_866, n_1259);
	not g1059(n_1329, n_1328);
	nor g1060(n_1256, ctl_sel_prim_412_12_n_538, n_1313, n_1325, prim_out[1]);
	not g1061(n_1330, n_1256);
	nand g1062(n_725, n_870, prim_out[5], n_1329, n_1330);
	nand g1063(n_663, n_1323, n_1324);
	nand g1064(n_1331, n_855, n_865, n_868, n_1259);
	not g1065(n_1332, n_1331);
	nand g1066(n_1333, n_877, n_869, n_872, n_1330);
	not g1067(n_1334, n_1333);
	nand g1068(sub_wire22, n_1332, n_1334);
	nand g1069(n_1335, n_855, n_872, n_863, n_1259);
	not g1070(n_1336, n_1335);
	nand g1071(n_1337, n_876, n_877, prim_out[5], n_1330);
	not g1072(n_1338, n_1337);
	nand g1073(n_749, n_1336, n_1338);
	nand g1074(sub_wire23, n_1330, n_1259);
	not g1075(n_1339, prim_out[7]);
	nand g1076(sub_wire24, prim_out[5], n_1339);
	not g1077(n_1340, prim_out[14]);
	nand g1078(n_717, n_863, n_1340);
	nand g1079(n_1341, n_856, n_863, n_870, n_1259);
	not g1080(n_1342, n_1341);
	nand g1081(n_1343, n_856, n_873, n_874, n_1259);
	not g1082(n_1344, n_1343);
	nand g1083(n_1345, n_1315, n_1316, n_1317, n_876);
	not g1084(n_1346, n_1345);
	nand g1085(n_1347, n_1311, n_1312, n_1314, n_1321);
	not g1086(n_1348, n_1347);
	nand g1087(n_1349, n_1322, n_876, n_883, n_884);
	not g1088(n_1350, n_1349);
	nand g1089(sub_wire8, n_877, n_1346);
	nand g1090(sub_wire25, n_877, n_1348);
	not g1091(n_1351, prim_out[15]);
	nand g1092(sub_wire1, n_877, n_1350);
	nand g1093(sub_wire10, prim_out[5], n_1342, n_1330);
	nand g1094(sub_wire3, prim_out[5], n_1344, n_1330);
	nand g1095(sub_wire26, prim_out[5], n_1351);
	and _ECO_0(w_eco0, sel_prim[0], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1(w_eco1, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_2(w_eco2, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_3(w_eco3, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_4(w_eco4, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_5(w_eco5, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_6(w_eco6, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_7(w_eco7, !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_8(w_eco8, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_9(w_eco9, sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_10(w_eco10, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_11(w_eco11, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_12(w_eco12, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_13(w_eco13, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_14(w_eco14, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_15(w_eco15, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_16(w_eco16, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_17(w_eco17, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_18(w_eco18, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_19(w_eco19, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_20(w_eco20, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_21(w_eco21, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_22(w_eco22, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_23(w_eco23, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_24(w_eco24, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_25(w_eco25, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_26(w_eco26, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_27(w_eco27, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_28(w_eco28, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_29(w_eco29, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_30(w_eco30, sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_31(w_eco31, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_32(w_eco32, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_33(w_eco33, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_34(w_eco34, sel_prim[0], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_35(w_eco35, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_36(w_eco36, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_37(w_eco37, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_38(w_eco38, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_39(w_eco39, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_40(w_eco40, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_41(w_eco41, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_42(w_eco42, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_43(w_eco43, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_44(w_eco44, !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_45(w_eco45, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_46(w_eco46, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_47(w_eco47, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_48(w_eco48, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_49(w_eco49, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_50(w_eco50, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_51(w_eco51, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_52(w_eco52, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_53(w_eco53, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_54(w_eco54, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_55(w_eco55, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_56(w_eco56, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_57(w_eco57, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_58(w_eco58, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_59(w_eco59, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_60(w_eco60, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_61(w_eco61, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_62(w_eco62, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_63(w_eco63, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_64(w_eco64, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_65(w_eco65, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_66(w_eco66, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_67(w_eco67, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6]);
	and _ECO_68(w_eco68, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_69(w_eco69, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_70(w_eco70, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_71(w_eco71, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_72(w_eco72, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_73(w_eco73, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_74(w_eco74, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_75(w_eco75, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_76(w_eco76, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_77(w_eco77, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_78(w_eco78, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_79(w_eco79, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_80(w_eco80, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[5]);
	and _ECO_81(w_eco81, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_82(w_eco82, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_83(w_eco83, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_84(w_eco84, !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_85(w_eco85, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_86(w_eco86, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_87(w_eco87, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_88(w_eco88, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_89(w_eco89, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_90(w_eco90, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_91(w_eco91, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_92(w_eco92, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_93(w_eco93, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_94(w_eco94, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_95(w_eco95, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_96(w_eco96, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_97(w_eco97, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96);
	xor _ECO_out0(prim_out[8], sub_wire0, w_eco97);
	and _ECO_98(w_eco98, sel_prim[0], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_99(w_eco99, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_100(w_eco100, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_101(w_eco101, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_102(w_eco102, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_103(w_eco103, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_104(w_eco104, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_105(w_eco105, !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_106(w_eco106, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_107(w_eco107, sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_108(w_eco108, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_109(w_eco109, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_110(w_eco110, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_111(w_eco111, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_112(w_eco112, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_113(w_eco113, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_114(w_eco114, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_115(w_eco115, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_116(w_eco116, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_117(w_eco117, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_118(w_eco118, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_119(w_eco119, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_120(w_eco120, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_121(w_eco121, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_122(w_eco122, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_123(w_eco123, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_124(w_eco124, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_125(w_eco125, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_126(w_eco126, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_127(w_eco127, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_128(w_eco128, sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_129(w_eco129, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_130(w_eco130, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_131(w_eco131, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_132(w_eco132, sel_prim[0], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_133(w_eco133, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_134(w_eco134, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_135(w_eco135, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_136(w_eco136, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_137(w_eco137, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_138(w_eco138, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_139(w_eco139, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_140(w_eco140, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_141(w_eco141, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_142(w_eco142, !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_143(w_eco143, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_144(w_eco144, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_145(w_eco145, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_146(w_eco146, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_147(w_eco147, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_148(w_eco148, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_149(w_eco149, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_150(w_eco150, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_151(w_eco151, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_152(w_eco152, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_153(w_eco153, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_154(w_eco154, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_155(w_eco155, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_156(w_eco156, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_157(w_eco157, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_158(w_eco158, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_159(w_eco159, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_160(w_eco160, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_161(w_eco161, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_162(w_eco162, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_163(w_eco163, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_164(w_eco164, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_165(w_eco165, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6]);
	and _ECO_166(w_eco166, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_167(w_eco167, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_168(w_eco168, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_169(w_eco169, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_170(w_eco170, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_171(w_eco171, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_172(w_eco172, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_173(w_eco173, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_174(w_eco174, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_175(w_eco175, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_176(w_eco176, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_177(w_eco177, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_178(w_eco178, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[5]);
	and _ECO_179(w_eco179, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_180(w_eco180, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_181(w_eco181, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_182(w_eco182, !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_183(w_eco183, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_184(w_eco184, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_185(w_eco185, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_186(w_eco186, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_187(w_eco187, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_188(w_eco188, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_189(w_eco189, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_190(w_eco190, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_191(w_eco191, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_192(w_eco192, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_193(w_eco193, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_194(w_eco194, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_195(w_eco195, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194);
	xor _ECO_out1(prim_out[12], sub_wire1, w_eco195);
	and _ECO_196(w_eco196, sel_prim[0], sel_prim[11], !sel_prim[7]);
	and _ECO_197(w_eco197, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_198(w_eco198, sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_199(w_eco199, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_200(w_eco200, sel_prim[0], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_201(w_eco201, sel_prim[0], sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_202(w_eco202, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_203(w_eco203, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_204(w_eco204, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_205(w_eco205, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_206(w_eco206, sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_207(w_eco207, sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_208(w_eco208, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_209(w_eco209, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_210(w_eco210, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_211(w_eco211, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_212(w_eco212, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_213(w_eco213, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_214(w_eco214, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_215(w_eco215, sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_216(w_eco216, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_217(w_eco217, sel_prim[0], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_218(w_eco218, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_219(w_eco219, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_220(w_eco220, sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_221(w_eco221, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_222(w_eco222, sel_prim[0], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_223(w_eco223, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[18]);
	and _ECO_224(w_eco224, sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_225(w_eco225, sel_prim[0], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_226(w_eco226, sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_227(w_eco227, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_228(w_eco228, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_229(w_eco229, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_230(w_eco230, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], sel_prim[17]);
	and _ECO_231(w_eco231, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_232(w_eco232, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_233(w_eco233, !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_234(w_eco234, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_235(w_eco235, !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_236(w_eco236, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], !sel_prim[18]);
	and _ECO_237(w_eco237, sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_238(w_eco238, !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_239(w_eco239, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_240(w_eco240, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], sel_prim[17]);
	and _ECO_241(w_eco241, sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_242(w_eco242, sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	or _ECO_243(w_eco243, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242);
	xor _ECO_out2(prim_out[9], sub_wire2, w_eco243);
	and _ECO_244(w_eco244, sel_prim[0], sel_prim[11], !sel_prim[7]);
	and _ECO_245(w_eco245, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_246(w_eco246, sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_247(w_eco247, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_248(w_eco248, sel_prim[0], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_249(w_eco249, sel_prim[0], sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_250(w_eco250, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_251(w_eco251, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_252(w_eco252, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_253(w_eco253, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_254(w_eco254, sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_255(w_eco255, sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_256(w_eco256, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_257(w_eco257, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_258(w_eco258, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_259(w_eco259, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_260(w_eco260, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_261(w_eco261, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_262(w_eco262, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_263(w_eco263, sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_264(w_eco264, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_265(w_eco265, sel_prim[0], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_266(w_eco266, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_267(w_eco267, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_268(w_eco268, sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_269(w_eco269, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_270(w_eco270, sel_prim[0], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_271(w_eco271, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[18]);
	and _ECO_272(w_eco272, sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_273(w_eco273, sel_prim[0], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_274(w_eco274, sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_275(w_eco275, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_276(w_eco276, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_277(w_eco277, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_278(w_eco278, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], sel_prim[17]);
	and _ECO_279(w_eco279, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_280(w_eco280, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_281(w_eco281, !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_282(w_eco282, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_283(w_eco283, !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_284(w_eco284, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], !sel_prim[18]);
	and _ECO_285(w_eco285, sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_286(w_eco286, !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_287(w_eco287, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_288(w_eco288, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], sel_prim[17]);
	and _ECO_289(w_eco289, sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_290(w_eco290, sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	or _ECO_291(w_eco291, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290);
	xor _ECO_out3(prim_out[11], sub_wire3, w_eco291);
	and _ECO_292(w_eco292, sel_prim[0], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_293(w_eco293, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_294(w_eco294, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_295(w_eco295, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_296(w_eco296, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_297(w_eco297, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_298(w_eco298, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_299(w_eco299, !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_300(w_eco300, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_301(w_eco301, sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_302(w_eco302, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_303(w_eco303, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_304(w_eco304, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_305(w_eco305, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_306(w_eco306, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_307(w_eco307, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_308(w_eco308, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_309(w_eco309, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_310(w_eco310, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_311(w_eco311, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_312(w_eco312, sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_313(w_eco313, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_314(w_eco314, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_315(w_eco315, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_316(w_eco316, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_317(w_eco317, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_318(w_eco318, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_319(w_eco319, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_320(w_eco320, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_321(w_eco321, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_322(w_eco322, sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_323(w_eco323, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_324(w_eco324, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_325(w_eco325, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_326(w_eco326, sel_prim[0], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_327(w_eco327, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_328(w_eco328, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_329(w_eco329, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_330(w_eco330, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_331(w_eco331, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_332(w_eco332, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_333(w_eco333, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_334(w_eco334, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_335(w_eco335, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_336(w_eco336, !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_337(w_eco337, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_338(w_eco338, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_339(w_eco339, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_340(w_eco340, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_341(w_eco341, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_342(w_eco342, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_343(w_eco343, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_344(w_eco344, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_345(w_eco345, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_346(w_eco346, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_347(w_eco347, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_348(w_eco348, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_349(w_eco349, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_350(w_eco350, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_351(w_eco351, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_352(w_eco352, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_353(w_eco353, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_354(w_eco354, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_355(w_eco355, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_356(w_eco356, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_357(w_eco357, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_358(w_eco358, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_359(w_eco359, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6]);
	and _ECO_360(w_eco360, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_361(w_eco361, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_362(w_eco362, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_363(w_eco363, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_364(w_eco364, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[4]);
	and _ECO_365(w_eco365, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_366(w_eco366, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_367(w_eco367, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_368(w_eco368, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_369(w_eco369, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_370(w_eco370, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_371(w_eco371, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_372(w_eco372, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[5]);
	and _ECO_373(w_eco373, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_374(w_eco374, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_375(w_eco375, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_376(w_eco376, !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_377(w_eco377, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_378(w_eco378, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[5]);
	and _ECO_379(w_eco379, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_380(w_eco380, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_381(w_eco381, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[17]);
	and _ECO_382(w_eco382, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_383(w_eco383, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_384(w_eco384, !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_385(w_eco385, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[6]);
	and _ECO_386(w_eco386, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_387(w_eco387, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_388(w_eco388, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_389(w_eco389, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388);
	xor _ECO_out4(prim_out[10], sub_wire4, w_eco389);
	and _ECO_390(w_eco390, sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_391(w_eco391, sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_392(w_eco392, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_393(w_eco393, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_394(w_eco394, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_395(w_eco395, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_396(w_eco396, sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_397(w_eco397, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_398(w_eco398, !sel_prim[0], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_399(w_eco399, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_400(w_eco400, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[3]);
	and _ECO_401(w_eco401, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_402(w_eco402, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_403(w_eco403, sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_404(w_eco404, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_405(w_eco405, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_406(w_eco406, sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_407(w_eco407, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_408(w_eco408, sel_prim[0], !sel_prim[11], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_409(w_eco409, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], sel_prim[3]);
	and _ECO_410(w_eco410, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_411(w_eco411, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_412(w_eco412, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3]);
	and _ECO_413(w_eco413, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[3]);
	and _ECO_414(w_eco414, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_415(w_eco415, sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_416(w_eco416, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_417(w_eco417, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_418(w_eco418, sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_419(w_eco419, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_420(w_eco420, !sel_prim[0], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_421(w_eco421, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_422(w_eco422, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_423(w_eco423, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_424(w_eco424, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_425(w_eco425, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_426(w_eco426, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_427(w_eco427, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_428(w_eco428, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], sel_prim[3]);
	and _ECO_429(w_eco429, !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[17]);
	and _ECO_430(w_eco430, sel_prim[0], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3]);
	and _ECO_431(w_eco431, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[4]);
	and _ECO_432(w_eco432, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_433(w_eco433, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_434(w_eco434, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_435(w_eco435, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_436(w_eco436, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_437(w_eco437, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_438(w_eco438, sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_439(w_eco439, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_440(w_eco440, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_441(w_eco441, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_442(w_eco442, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_443(w_eco443, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_444(w_eco444, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_445(w_eco445, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14]);
	and _ECO_446(w_eco446, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[17]);
	and _ECO_447(w_eco447, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[4]);
	and _ECO_448(w_eco448, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_449(w_eco449, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[4], !sel_prim[17]);
	and _ECO_450(w_eco450, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14]);
	and _ECO_451(w_eco451, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_452(w_eco452, sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3]);
	and _ECO_453(w_eco453, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_454(w_eco454, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[4]);
	and _ECO_455(w_eco455, sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_456(w_eco456, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_457(w_eco457, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_458(w_eco458, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_459(w_eco459, sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_460(w_eco460, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[5], !sel_prim[6]);
	or _ECO_461(w_eco461, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460);
	xor _ECO_out5(prim_out[17], sub_wire5, w_eco461);
	and _ECO_462(w_eco462, sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_463(w_eco463, sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_464(w_eco464, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_465(w_eco465, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_466(w_eco466, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_467(w_eco467, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_468(w_eco468, sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_469(w_eco469, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_470(w_eco470, !sel_prim[0], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_471(w_eco471, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_472(w_eco472, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[3]);
	and _ECO_473(w_eco473, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_474(w_eco474, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_475(w_eco475, sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_476(w_eco476, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_477(w_eco477, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_478(w_eco478, sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_479(w_eco479, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_480(w_eco480, sel_prim[0], !sel_prim[11], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_481(w_eco481, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], sel_prim[3]);
	and _ECO_482(w_eco482, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_483(w_eco483, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_484(w_eco484, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3]);
	and _ECO_485(w_eco485, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[3]);
	and _ECO_486(w_eco486, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_487(w_eco487, sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_488(w_eco488, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_489(w_eco489, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_490(w_eco490, sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_491(w_eco491, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_492(w_eco492, !sel_prim[0], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_493(w_eco493, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_494(w_eco494, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_495(w_eco495, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_496(w_eco496, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_497(w_eco497, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_498(w_eco498, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_499(w_eco499, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_500(w_eco500, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], sel_prim[3]);
	and _ECO_501(w_eco501, !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[17]);
	and _ECO_502(w_eco502, sel_prim[0], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3]);
	and _ECO_503(w_eco503, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[4]);
	and _ECO_504(w_eco504, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_505(w_eco505, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_506(w_eco506, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_507(w_eco507, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_508(w_eco508, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_509(w_eco509, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_510(w_eco510, sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_511(w_eco511, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_512(w_eco512, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_513(w_eco513, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_514(w_eco514, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_515(w_eco515, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_516(w_eco516, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_517(w_eco517, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14]);
	and _ECO_518(w_eco518, !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[17]);
	and _ECO_519(w_eco519, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[4]);
	and _ECO_520(w_eco520, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_521(w_eco521, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[4], !sel_prim[17]);
	and _ECO_522(w_eco522, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14]);
	and _ECO_523(w_eco523, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_524(w_eco524, sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3]);
	and _ECO_525(w_eco525, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_526(w_eco526, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[4]);
	and _ECO_527(w_eco527, sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_528(w_eco528, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_529(w_eco529, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_530(w_eco530, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_531(w_eco531, sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_532(w_eco532, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[5], !sel_prim[6]);
	or _ECO_533(w_eco533, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532);
	xor _ECO_out6(prim_out[25], sub_wire6, w_eco533);
	and _ECO_534(w_eco534, !sel_prim[15], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_535(w_eco535, sel_prim[11], !sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_536(w_eco536, sel_prim[0], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_537(w_eco537, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_538(w_eco538, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_539(w_eco539, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_540(w_eco540, sel_prim[0], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_541(w_eco541, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_542(w_eco542, !sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_543(w_eco543, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_544(w_eco544, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[5]);
	and _ECO_545(w_eco545, !sel_prim[15], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_546(w_eco546, !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_547(w_eco547, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11]);
	and _ECO_548(w_eco548, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_549(w_eco549, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[3]);
	and _ECO_550(w_eco550, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8]);
	and _ECO_551(w_eco551, sel_prim[0], !sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_552(w_eco552, !sel_prim[0], sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_553(w_eco553, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_554(w_eco554, sel_prim[0], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_555(w_eco555, !sel_prim[1], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_556(w_eco556, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_557(w_eco557, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[3]);
	and _ECO_558(w_eco558, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_559(w_eco559, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_560(w_eco560, !sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_561(w_eco561, !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_562(w_eco562, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_563(w_eco563, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8]);
	and _ECO_564(w_eco564, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_565(w_eco565, !sel_prim[0], sel_prim[1], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_566(w_eco566, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[3], sel_prim[5]);
	and _ECO_567(w_eco567, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_568(w_eco568, !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_569(w_eco569, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_570(w_eco570, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_571(w_eco571, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[8]);
	and _ECO_572(w_eco572, sel_prim[0], !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_573(w_eco573, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_574(w_eco574, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_575(w_eco575, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[3]);
	and _ECO_576(w_eco576, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[13]);
	and _ECO_577(w_eco577, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[9], sel_prim[10]);
	and _ECO_578(w_eco578, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_579(w_eco579, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7]);
	and _ECO_580(w_eco580, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_581(w_eco581, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[18]);
	and _ECO_582(w_eco582, sel_prim[0], !sel_prim[11], !sel_prim[9], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_583(w_eco583, !sel_prim[0], sel_prim[2], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_584(w_eco584, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_585(w_eco585, !sel_prim[0], sel_prim[1], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_586(w_eco586, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_587(w_eco587, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_588(w_eco588, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_589(w_eco589, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_590(w_eco590, !sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_591(w_eco591, !sel_prim[1], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_592(w_eco592, !sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_593(w_eco593, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[6]);
	and _ECO_594(w_eco594, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_595(w_eco595, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_596(w_eco596, !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_597(w_eco597, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_598(w_eco598, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_599(w_eco599, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_600(w_eco600, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], sel_prim[3]);
	and _ECO_601(w_eco601, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[10]);
	and _ECO_602(w_eco602, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_603(w_eco603, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[17]);
	and _ECO_604(w_eco604, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[18]);
	and _ECO_605(w_eco605, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_606(w_eco606, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_607(w_eco607, !sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_608(w_eco608, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[5]);
	and _ECO_609(w_eco609, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5]);
	and _ECO_610(w_eco610, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_611(w_eco611, !sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_612(w_eco612, !sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_613(w_eco613, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[6]);
	and _ECO_614(w_eco614, sel_prim[0], !sel_prim[11], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_615(w_eco615, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_616(w_eco616, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_617(w_eco617, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_618(w_eco618, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_619(w_eco619, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_620(w_eco620, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_621(w_eco621, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_622(w_eco622, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_623(w_eco623, !sel_prim[1], !sel_prim[2], !sel_prim[12], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_624(w_eco624, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[4]);
	and _ECO_625(w_eco625, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[17]);
	and _ECO_626(w_eco626, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_627(w_eco627, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_628(w_eco628, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[9]);
	and _ECO_629(w_eco629, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4]);
	and _ECO_630(w_eco630, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[5]);
	and _ECO_631(w_eco631, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_632(w_eco632, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[5]);
	and _ECO_633(w_eco633, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_634(w_eco634, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_635(w_eco635, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_636(w_eco636, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_637(w_eco637, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5]);
	and _ECO_638(w_eco638, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	and _ECO_639(w_eco639, !sel_prim[11], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_640(w_eco640, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_641(w_eco641, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_642(w_eco642, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_643(w_eco643, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_644(w_eco644, !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_645(w_eco645, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_646(w_eco646, !sel_prim[1], !sel_prim[2], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_647(w_eco647, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[4]);
	and _ECO_648(w_eco648, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_649(w_eco649, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_650(w_eco650, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[5]);
	and _ECO_651(w_eco651, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_652(w_eco652, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_653(w_eco653, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_654(w_eco654, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], !sel_prim[4]);
	and _ECO_655(w_eco655, !sel_prim[15], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_656(w_eco656, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_657(w_eco657, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_658(w_eco658, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[9], sel_prim[10], !sel_prim[4]);
	and _ECO_659(w_eco659, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[5], sel_prim[6]);
	and _ECO_660(w_eco660, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_661(w_eco661, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[4]);
	and _ECO_662(w_eco662, !sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_663(w_eco663, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_664(w_eco664, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_665(w_eco665, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_666(w_eco666, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_667(w_eco667, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[3], !sel_prim[6]);
	and _ECO_668(w_eco668, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_669(w_eco669, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[10]);
	and _ECO_670(w_eco670, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_671(w_eco671, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_672(w_eco672, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_673(w_eco673, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[3], sel_prim[4]);
	and _ECO_674(w_eco674, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_675(w_eco675, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_676(w_eco676, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_677(w_eco677, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_678(w_eco678, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_679(w_eco679, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[7], !sel_prim[5]);
	and _ECO_680(w_eco680, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[5], sel_prim[6]);
	and _ECO_681(w_eco681, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[4], !sel_prim[5]);
	and _ECO_682(w_eco682, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_683(w_eco683, sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_684(w_eco684, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], !sel_prim[3], !sel_prim[4], !sel_prim[6], !sel_prim[17]);
	and _ECO_685(w_eco685, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[3], sel_prim[4]);
	and _ECO_686(w_eco686, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[9], sel_prim[10], !sel_prim[4]);
	and _ECO_687(w_eco687, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[10], !sel_prim[5]);
	and _ECO_688(w_eco688, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_689(w_eco689, !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_690(w_eco690, sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[9], !sel_prim[4], !sel_prim[5]);
	and _ECO_691(w_eco691, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[9], !sel_prim[4]);
	and _ECO_692(w_eco692, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[13], !sel_prim[3], !sel_prim[6]);
	and _ECO_693(w_eco693, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], !sel_prim[3], !sel_prim[4], !sel_prim[6], !sel_prim[17]);
	and _ECO_694(w_eco694, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[9], !sel_prim[5]);
	and _ECO_695(w_eco695, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_696(w_eco696, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_697(w_eco697, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[13], !sel_prim[3], !sel_prim[6]);
	and _ECO_698(w_eco698, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	or _ECO_699(w_eco699, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698);
	xor _ECO_out7(prim_out[18], sub_wire7, w_eco699);
	and _ECO_700(w_eco700, !sel_prim[15], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_701(w_eco701, sel_prim[11], !sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_702(w_eco702, sel_prim[0], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_703(w_eco703, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_704(w_eco704, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_705(w_eco705, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_706(w_eco706, sel_prim[0], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_707(w_eco707, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_708(w_eco708, !sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[3]);
	and _ECO_709(w_eco709, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_710(w_eco710, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[5]);
	and _ECO_711(w_eco711, !sel_prim[15], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_712(w_eco712, !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_713(w_eco713, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11]);
	and _ECO_714(w_eco714, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_715(w_eco715, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[3]);
	and _ECO_716(w_eco716, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8]);
	and _ECO_717(w_eco717, sel_prim[0], !sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_718(w_eco718, !sel_prim[0], sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_719(w_eco719, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_720(w_eco720, sel_prim[0], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_721(w_eco721, !sel_prim[1], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_722(w_eco722, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_723(w_eco723, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[3]);
	and _ECO_724(w_eco724, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_725(w_eco725, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_726(w_eco726, !sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_727(w_eco727, !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_728(w_eco728, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_729(w_eco729, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8]);
	and _ECO_730(w_eco730, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_731(w_eco731, !sel_prim[0], sel_prim[1], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_732(w_eco732, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[3], sel_prim[5]);
	and _ECO_733(w_eco733, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_734(w_eco734, !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_735(w_eco735, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_736(w_eco736, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_737(w_eco737, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[8]);
	and _ECO_738(w_eco738, sel_prim[0], !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_739(w_eco739, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_740(w_eco740, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_741(w_eco741, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[3]);
	and _ECO_742(w_eco742, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[13]);
	and _ECO_743(w_eco743, sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[9], sel_prim[10]);
	and _ECO_744(w_eco744, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_745(w_eco745, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7]);
	and _ECO_746(w_eco746, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_747(w_eco747, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[18]);
	and _ECO_748(w_eco748, sel_prim[0], !sel_prim[11], !sel_prim[9], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_749(w_eco749, !sel_prim[0], sel_prim[2], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_750(w_eco750, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_751(w_eco751, !sel_prim[0], sel_prim[1], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_752(w_eco752, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_753(w_eco753, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_754(w_eco754, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_755(w_eco755, !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_756(w_eco756, !sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_757(w_eco757, !sel_prim[1], sel_prim[11], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_758(w_eco758, !sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_759(w_eco759, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[6]);
	and _ECO_760(w_eco760, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_761(w_eco761, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_762(w_eco762, !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_763(w_eco763, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_764(w_eco764, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_765(w_eco765, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_766(w_eco766, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], sel_prim[3]);
	and _ECO_767(w_eco767, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[10]);
	and _ECO_768(w_eco768, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_769(w_eco769, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[17]);
	and _ECO_770(w_eco770, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[18]);
	and _ECO_771(w_eco771, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_772(w_eco772, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_773(w_eco773, !sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_774(w_eco774, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[5]);
	and _ECO_775(w_eco775, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5]);
	and _ECO_776(w_eco776, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_777(w_eco777, !sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_778(w_eco778, !sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_779(w_eco779, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[6]);
	and _ECO_780(w_eco780, sel_prim[0], !sel_prim[11], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_781(w_eco781, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_782(w_eco782, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_783(w_eco783, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_784(w_eco784, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_785(w_eco785, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_786(w_eco786, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_787(w_eco787, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_788(w_eco788, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_789(w_eco789, !sel_prim[1], !sel_prim[2], !sel_prim[12], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_790(w_eco790, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[4]);
	and _ECO_791(w_eco791, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[4], sel_prim[17]);
	and _ECO_792(w_eco792, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_793(w_eco793, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_794(w_eco794, sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[9]);
	and _ECO_795(w_eco795, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4]);
	and _ECO_796(w_eco796, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[3], sel_prim[5]);
	and _ECO_797(w_eco797, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_798(w_eco798, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[5]);
	and _ECO_799(w_eco799, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_800(w_eco800, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_801(w_eco801, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_802(w_eco802, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_803(w_eco803, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5]);
	and _ECO_804(w_eco804, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	and _ECO_805(w_eco805, !sel_prim[11], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_806(w_eco806, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_807(w_eco807, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_808(w_eco808, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_809(w_eco809, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_810(w_eco810, !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_811(w_eco811, !sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_812(w_eco812, !sel_prim[1], !sel_prim[2], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_813(w_eco813, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[4]);
	and _ECO_814(w_eco814, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_815(w_eco815, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_816(w_eco816, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[3], sel_prim[5]);
	and _ECO_817(w_eco817, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_818(w_eco818, sel_prim[0], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_819(w_eco819, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_820(w_eco820, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[8], !sel_prim[4]);
	and _ECO_821(w_eco821, !sel_prim[15], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_822(w_eco822, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_823(w_eco823, sel_prim[0], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_824(w_eco824, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[9], sel_prim[10], !sel_prim[4]);
	and _ECO_825(w_eco825, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[5], sel_prim[6]);
	and _ECO_826(w_eco826, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_827(w_eco827, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[4]);
	and _ECO_828(w_eco828, !sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_829(w_eco829, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_830(w_eco830, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_831(w_eco831, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_832(w_eco832, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_833(w_eco833, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[3], !sel_prim[6]);
	and _ECO_834(w_eco834, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_835(w_eco835, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[10]);
	and _ECO_836(w_eco836, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_837(w_eco837, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_838(w_eco838, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_839(w_eco839, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[3], sel_prim[4]);
	and _ECO_840(w_eco840, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_841(w_eco841, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[5]);
	and _ECO_842(w_eco842, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_843(w_eco843, !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_844(w_eco844, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_845(w_eco845, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[7], !sel_prim[5]);
	and _ECO_846(w_eco846, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[5], sel_prim[6]);
	and _ECO_847(w_eco847, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[4], !sel_prim[5]);
	and _ECO_848(w_eco848, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_849(w_eco849, sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_850(w_eco850, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[13], !sel_prim[3], !sel_prim[4], !sel_prim[6], !sel_prim[17]);
	and _ECO_851(w_eco851, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[3], sel_prim[4]);
	and _ECO_852(w_eco852, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[9], sel_prim[10], !sel_prim[4]);
	and _ECO_853(w_eco853, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[10], !sel_prim[5]);
	and _ECO_854(w_eco854, !sel_prim[1], !sel_prim[2], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_855(w_eco855, !sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_856(w_eco856, sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[8], sel_prim[9], !sel_prim[4], !sel_prim[5]);
	and _ECO_857(w_eco857, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[9], !sel_prim[4]);
	and _ECO_858(w_eco858, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[13], !sel_prim[3], !sel_prim[6]);
	and _ECO_859(w_eco859, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[13], !sel_prim[3], !sel_prim[4], !sel_prim[6], !sel_prim[17]);
	and _ECO_860(w_eco860, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[8], sel_prim[9], !sel_prim[5]);
	and _ECO_861(w_eco861, !sel_prim[1], !sel_prim[2], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_862(w_eco862, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_863(w_eco863, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[13], !sel_prim[3], !sel_prim[6]);
	and _ECO_864(w_eco864, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	or _ECO_865(w_eco865, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864);
	xor _ECO_out8(prim_out[26], sub_wire8, w_eco865);
	and _ECO_866(w_eco866, sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_867(w_eco867, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_868(w_eco868, sel_prim[11], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_869(w_eco869, sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_870(w_eco870, !sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[3]);
	and _ECO_871(w_eco871, sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_872(w_eco872, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_873(w_eco873, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[3]);
	and _ECO_874(w_eco874, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[7]);
	and _ECO_875(w_eco875, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_876(w_eco876, !sel_prim[0], sel_prim[2], sel_prim[12], sel_prim[8]);
	and _ECO_877(w_eco877, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12]);
	and _ECO_878(w_eco878, sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_879(w_eco879, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[4], sel_prim[5]);
	and _ECO_880(w_eco880, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[3]);
	and _ECO_881(w_eco881, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7]);
	and _ECO_882(w_eco882, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[10], sel_prim[4]);
	and _ECO_883(w_eco883, !sel_prim[0], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_884(w_eco884, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12]);
	and _ECO_885(w_eco885, !sel_prim[0], sel_prim[2], !sel_prim[13], sel_prim[8]);
	and _ECO_886(w_eco886, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[13]);
	and _ECO_887(w_eco887, sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_888(w_eco888, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_889(w_eco889, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[9], sel_prim[4]);
	and _ECO_890(w_eco890, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[10], sel_prim[4]);
	and _ECO_891(w_eco891, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_892(w_eco892, !sel_prim[0], !sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_893(w_eco893, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[13]);
	and _ECO_894(w_eco894, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[4]);
	and _ECO_895(w_eco895, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_896(w_eco896, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[7], sel_prim[3]);
	and _ECO_897(w_eco897, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_898(w_eco898, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[3]);
	and _ECO_899(w_eco899, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[9], sel_prim[4]);
	and _ECO_900(w_eco900, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_901(w_eco901, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_902(w_eco902, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_903(w_eco903, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[4], sel_prim[6]);
	and _ECO_904(w_eco904, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[10], !sel_prim[5], !sel_prim[6]);
	and _ECO_905(w_eco905, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[7], sel_prim[3]);
	and _ECO_906(w_eco906, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_907(w_eco907, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_908(w_eco908, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_909(w_eco909, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[4]);
	and _ECO_910(w_eco910, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[4], sel_prim[6]);
	and _ECO_911(w_eco911, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[9], !sel_prim[5], !sel_prim[6]);
	and _ECO_912(w_eco912, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_913(w_eco913, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_914(w_eco914, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[4], !sel_prim[5]);
	and _ECO_915(w_eco915, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_916(w_eco916, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_917(w_eco917, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_918(w_eco918, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917);
	xor _ECO_out9(prim_out[19], sub_wire9, w_eco918);
	and _ECO_919(w_eco919, sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_920(w_eco920, sel_prim[11], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_921(w_eco921, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[3]);
	and _ECO_922(w_eco922, sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_923(w_eco923, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_924(w_eco924, sel_prim[0], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_925(w_eco925, sel_prim[0], !sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_926(w_eco926, !sel_prim[0], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_927(w_eco927, !sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_928(w_eco928, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_929(w_eco929, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_930(w_eco930, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_931(w_eco931, sel_prim[0], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_932(w_eco932, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_933(w_eco933, !sel_prim[0], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_934(w_eco934, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[3]);
	and _ECO_935(w_eco935, sel_prim[1], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_936(w_eco936, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_937(w_eco937, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_938(w_eco938, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_939(w_eco939, !sel_prim[0], sel_prim[1], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_940(w_eco940, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_941(w_eco941, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_942(w_eco942, !sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_943(w_eco943, !sel_prim[0], !sel_prim[2], sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_944(w_eco944, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_945(w_eco945, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_946(w_eco946, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_947(w_eco947, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_948(w_eco948, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[3]);
	and _ECO_949(w_eco949, !sel_prim[0], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_950(w_eco950, !sel_prim[0], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_951(w_eco951, sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_952(w_eco952, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3]);
	and _ECO_953(w_eco953, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_954(w_eco954, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_955(w_eco955, !sel_prim[0], sel_prim[1], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_956(w_eco956, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_957(w_eco957, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_958(w_eco958, !sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_959(w_eco959, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[7], sel_prim[3]);
	and _ECO_960(w_eco960, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_961(w_eco961, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_962(w_eco962, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_963(w_eco963, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[4], sel_prim[5]);
	and _ECO_964(w_eco964, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_965(w_eco965, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[3]);
	and _ECO_966(w_eco966, !sel_prim[0], sel_prim[1], !sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[18]);
	and _ECO_967(w_eco967, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_968(w_eco968, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_969(w_eco969, !sel_prim[0], !sel_prim[1], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_970(w_eco970, !sel_prim[0], sel_prim[1], !sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_971(w_eco971, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_972(w_eco972, !sel_prim[0], sel_prim[1], !sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[17]);
	and _ECO_973(w_eco973, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_974(w_eco974, !sel_prim[0], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[18]);
	and _ECO_975(w_eco975, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_976(w_eco976, !sel_prim[1], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_977(w_eco977, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_978(w_eco978, !sel_prim[0], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], sel_prim[17]);
	and _ECO_979(w_eco979, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_980(w_eco980, !sel_prim[0], !sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[18]);
	and _ECO_981(w_eco981, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4]);
	and _ECO_982(w_eco982, !sel_prim[0], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_983(w_eco983, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_984(w_eco984, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_985(w_eco985, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_986(w_eco986, !sel_prim[0], !sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[17]);
	and _ECO_987(w_eco987, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_988(w_eco988, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_989(w_eco989, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_990(w_eco990, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[18]);
	and _ECO_991(w_eco991, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4]);
	and _ECO_992(w_eco992, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_993(w_eco993, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[17]);
	or _ECO_994(w_eco994, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993);
	xor _ECO_out10(prim_out[27], sub_wire10, w_eco994);
	and _ECO_995(w_eco995, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_996(w_eco996, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_997(w_eco997, sel_prim[0], sel_prim[7], sel_prim[3]);
	and _ECO_998(w_eco998, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_999(w_eco999, sel_prim[0], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_1000(w_eco1000, !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_1001(w_eco1001, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[3]);
	and _ECO_1002(w_eco1002, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1003(w_eco1003, !sel_prim[0], sel_prim[2], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1004(w_eco1004, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1005(w_eco1005, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_1006(w_eco1006, sel_prim[0], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1007(w_eco1007, !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_1008(w_eco1008, !sel_prim[1], sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[8], sel_prim[3]);
	and _ECO_1009(w_eco1009, !sel_prim[11], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_1010(w_eco1010, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[3]);
	and _ECO_1011(w_eco1011, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[3]);
	and _ECO_1012(w_eco1012, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4]);
	and _ECO_1013(w_eco1013, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1014(w_eco1014, sel_prim[1], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_1015(w_eco1015, !sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1016(w_eco1016, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_1017(w_eco1017, !sel_prim[1], !sel_prim[2], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1018(w_eco1018, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1019(w_eco1019, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1020(w_eco1020, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[7], !sel_prim[3]);
	and _ECO_1021(w_eco1021, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4]);
	and _ECO_1022(w_eco1022, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4]);
	and _ECO_1023(w_eco1023, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1024(w_eco1024, !sel_prim[0], sel_prim[2], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1025(w_eco1025, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_1026(w_eco1026, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1027(w_eco1027, !sel_prim[1], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_1028(w_eco1028, sel_prim[1], !sel_prim[11], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1029(w_eco1029, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1030(w_eco1030, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1031(w_eco1031, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4]);
	and _ECO_1032(w_eco1032, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1033(w_eco1033, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4]);
	and _ECO_1034(w_eco1034, !sel_prim[0], sel_prim[1], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1035(w_eco1035, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4]);
	and _ECO_1036(w_eco1036, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1037(w_eco1037, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[4]);
	and _ECO_1038(w_eco1038, !sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1039(w_eco1039, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1040(w_eco1040, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	or _ECO_1041(w_eco1041, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040);
	xor _ECO_out11(prim_out[22], sub_wire11, w_eco1041);
	and _ECO_1042(w_eco1042, !sel_prim[0], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_1043(w_eco1043, sel_prim[0], !sel_prim[3]);
	and _ECO_1044(w_eco1044, sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1045(w_eco1045, !sel_prim[0], !sel_prim[2], sel_prim[11], sel_prim[3]);
	and _ECO_1046(w_eco1046, !sel_prim[0], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1047(w_eco1047, !sel_prim[0], !sel_prim[2], !sel_prim[7], sel_prim[3]);
	and _ECO_1048(w_eco1048, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[4]);
	and _ECO_1049(w_eco1049, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1050(w_eco1050, !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4]);
	and _ECO_1051(w_eco1051, sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10]);
	and _ECO_1052(w_eco1052, !sel_prim[0], sel_prim[1], !sel_prim[7], sel_prim[3]);
	and _ECO_1053(w_eco1053, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1054(w_eco1054, !sel_prim[1], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1055(w_eco1055, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7], sel_prim[4]);
	and _ECO_1056(w_eco1056, sel_prim[2], sel_prim[11], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1057(w_eco1057, !sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3]);
	and _ECO_1058(w_eco1058, !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3]);
	and _ECO_1059(w_eco1059, !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5]);
	and _ECO_1060(w_eco1060, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[5], !sel_prim[6]);
	and _ECO_1061(w_eco1061, sel_prim[0], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_1062(w_eco1062, sel_prim[2], sel_prim[11], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1063(w_eco1063, sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10]);
	and _ECO_1064(w_eco1064, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[8], sel_prim[9], sel_prim[4]);
	and _ECO_1065(w_eco1065, !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[10], !sel_prim[3]);
	and _ECO_1066(w_eco1066, !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1067(w_eco1067, !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3]);
	and _ECO_1068(w_eco1068, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[5], !sel_prim[6]);
	and _ECO_1069(w_eco1069, !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1070(w_eco1070, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], sel_prim[3]);
	and _ECO_1071(w_eco1071, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], sel_prim[10]);
	and _ECO_1072(w_eco1072, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1073(w_eco1073, !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1074(w_eco1074, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8]);
	and _ECO_1075(w_eco1075, !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[9], !sel_prim[3]);
	and _ECO_1076(w_eco1076, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_1077(w_eco1077, !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[3]);
	and _ECO_1078(w_eco1078, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[4]);
	and _ECO_1079(w_eco1079, !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1080(w_eco1080, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[12], !sel_prim[14], sel_prim[3]);
	and _ECO_1081(w_eco1081, sel_prim[0], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], sel_prim[10]);
	and _ECO_1082(w_eco1082, !sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[3]);
	and _ECO_1083(w_eco1083, !sel_prim[1], !sel_prim[15], sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_1084(w_eco1084, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[4]);
	and _ECO_1085(w_eco1085, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[4]);
	and _ECO_1086(w_eco1086, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[9], sel_prim[10]);
	and _ECO_1087(w_eco1087, !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[9], !sel_prim[3]);
	and _ECO_1088(w_eco1088, !sel_prim[1], sel_prim[2], !sel_prim[15], sel_prim[16], sel_prim[12], !sel_prim[3], sel_prim[4]);
	or _ECO_1089(w_eco1089, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088);
	xor _ECO_out12(prim_out[30], sub_wire12, w_eco1089);
	and _ECO_1090(w_eco1090, sel_prim[0], !sel_prim[11], sel_prim[3]);
	and _ECO_1091(w_eco1091, sel_prim[2], !sel_prim[11], sel_prim[3]);
	and _ECO_1092(w_eco1092, sel_prim[0], !sel_prim[3], sel_prim[4]);
	and _ECO_1093(w_eco1093, !sel_prim[0], sel_prim[2], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1094(w_eco1094, sel_prim[1], !sel_prim[11], sel_prim[3]);
	and _ECO_1095(w_eco1095, !sel_prim[0], sel_prim[1], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1096(w_eco1096, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1097(w_eco1097, !sel_prim[1], !sel_prim[2], !sel_prim[3], sel_prim[4]);
	and _ECO_1098(w_eco1098, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1099(w_eco1099, sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1100(w_eco1100, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1101(w_eco1101, sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[4], sel_prim[17]);
	and _ECO_1102(w_eco1102, sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1103(w_eco1103, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1104(w_eco1104, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1105(w_eco1105, sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], sel_prim[17]);
	and _ECO_1106(w_eco1106, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1107(w_eco1107, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1108(w_eco1108, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1109(w_eco1109, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1110(w_eco1110, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1111(w_eco1111, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1112(w_eco1112, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1113(w_eco1113, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1114(w_eco1114, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	or _ECO_1115(w_eco1115, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114);
	xor _ECO_out13(prim_out[23], sub_wire13, w_eco1115);
	and _ECO_1116(w_eco1116, !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1117(w_eco1117, sel_prim[0], sel_prim[11]);
	and _ECO_1118(w_eco1118, !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1119(w_eco1119, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[3]);
	and _ECO_1120(w_eco1120, !sel_prim[15], sel_prim[11], !sel_prim[4]);
	and _ECO_1121(w_eco1121, !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1122(w_eco1122, !sel_prim[1], !sel_prim[2], sel_prim[11]);
	and _ECO_1123(w_eco1123, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[12]);
	and _ECO_1124(w_eco1124, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1125(w_eco1125, sel_prim[0], !sel_prim[3]);
	and _ECO_1126(w_eco1126, sel_prim[2], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1127(w_eco1127, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], sel_prim[3]);
	and _ECO_1128(w_eco1128, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[3]);
	and _ECO_1129(w_eco1129, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1130(w_eco1130, sel_prim[1], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1131(w_eco1131, sel_prim[1], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1132(w_eco1132, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13]);
	and _ECO_1133(w_eco1133, sel_prim[2], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1134(w_eco1134, !sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1135(w_eco1135, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1136(w_eco1136, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14]);
	and _ECO_1137(w_eco1137, sel_prim[1], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1138(w_eco1138, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1139(w_eco1139, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[3]);
	and _ECO_1140(w_eco1140, sel_prim[1], !sel_prim[15], !sel_prim[16], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[17]);
	and _ECO_1141(w_eco1141, sel_prim[1], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1142(w_eco1142, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_1143(w_eco1143, sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4]);
	and _ECO_1144(w_eco1144, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1145(w_eco1145, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1146(w_eco1146, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8]);
	and _ECO_1147(w_eco1147, !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1148(w_eco1148, sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4]);
	and _ECO_1149(w_eco1149, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4]);
	and _ECO_1150(w_eco1150, !sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[3], !sel_prim[4]);
	and _ECO_1151(w_eco1151, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1152(w_eco1152, sel_prim[1], !sel_prim[15], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[17]);
	and _ECO_1153(w_eco1153, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1154(w_eco1154, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], sel_prim[17]);
	and _ECO_1155(w_eco1155, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4]);
	and _ECO_1156(w_eco1156, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[7], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1157(w_eco1157, sel_prim[2], !sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1158(w_eco1158, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1159(w_eco1159, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[7], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1160(w_eco1160, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1161(w_eco1161, sel_prim[1], !sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1162(w_eco1162, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[17]);
	and _ECO_1163(w_eco1163, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], sel_prim[17]);
	and _ECO_1164(w_eco1164, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1165(w_eco1165, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4]);
	and _ECO_1166(w_eco1166, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[17]);
	and _ECO_1167(w_eco1167, !sel_prim[0], !sel_prim[15], sel_prim[16], !sel_prim[12], !sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4]);
	or _ECO_1168(w_eco1168, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167);
	xor _ECO_out14(prim_out[31], sub_wire14, w_eco1168);
	and _ECO_1169(w_eco1169, sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_1170(w_eco1170, sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1171(w_eco1171, !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1172(w_eco1172, sel_prim[0], sel_prim[11], sel_prim[8], !sel_prim[4]);
	and _ECO_1173(w_eco1173, !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_1174(w_eco1174, !sel_prim[0], sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[4]);
	and _ECO_1175(w_eco1175, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_1176(w_eco1176, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4]);
	and _ECO_1177(w_eco1177, sel_prim[11], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1178(w_eco1178, !sel_prim[0], sel_prim[1], sel_prim[11], sel_prim[7], sel_prim[4]);
	and _ECO_1179(w_eco1179, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1180(w_eco1180, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13]);
	and _ECO_1181(w_eco1181, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[8], !sel_prim[4]);
	and _ECO_1182(w_eco1182, sel_prim[0], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1183(w_eco1183, sel_prim[11], sel_prim[7], !sel_prim[4], !sel_prim[5]);
	and _ECO_1184(w_eco1184, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1185(w_eco1185, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1186(w_eco1186, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1187(w_eco1187, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[4]);
	and _ECO_1188(w_eco1188, sel_prim[0], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1189(w_eco1189, !sel_prim[11], !sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1190(w_eco1190, !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1191(w_eco1191, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1192(w_eco1192, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1193(w_eco1193, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1194(w_eco1194, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1195(w_eco1195, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1196(w_eco1196, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1197(w_eco1197, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_1198(w_eco1198, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1199(w_eco1199, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1200(w_eco1200, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1201(w_eco1201, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1202(w_eco1202, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1203(w_eco1203, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_1204(w_eco1204, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1205(w_eco1205, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1206(w_eco1206, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1207(w_eco1207, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1208(w_eco1208, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_1209(w_eco1209, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1210(w_eco1210, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[17], sel_prim[18]);
	and _ECO_1211(w_eco1211, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_1212(w_eco1212, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1213(w_eco1213, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1214(w_eco1214, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5], !sel_prim[17], sel_prim[18]);
	and _ECO_1215(w_eco1215, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5]);
	and _ECO_1216(w_eco1216, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4], !sel_prim[17], sel_prim[18]);
	and _ECO_1217(w_eco1217, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1218(w_eco1218, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[17], sel_prim[18]);
	and _ECO_1219(w_eco1219, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8]);
	and _ECO_1220(w_eco1220, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1221(w_eco1221, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5], !sel_prim[17], sel_prim[18]);
	and _ECO_1222(w_eco1222, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5]);
	and _ECO_1223(w_eco1223, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[17], sel_prim[18]);
	and _ECO_1224(w_eco1224, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1225(w_eco1225, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], sel_prim[18]);
	and _ECO_1226(w_eco1226, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1227(w_eco1227, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[17], sel_prim[18]);
	and _ECO_1228(w_eco1228, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1229(w_eco1229, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], sel_prim[18]);
	and _ECO_1230(w_eco1230, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_1231(w_eco1231, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230);
	xor _ECO_out15(prim_out[1], sub_wire15, w_eco1231);
	and _ECO_1232(w_eco1232, sel_prim[0], !sel_prim[3], !sel_prim[4]);
	and _ECO_1233(w_eco1233, !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1234(w_eco1234, !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1235(w_eco1235, sel_prim[0], sel_prim[11], sel_prim[3]);
	and _ECO_1236(w_eco1236, !sel_prim[1], !sel_prim[2], !sel_prim[3], !sel_prim[4]);
	and _ECO_1237(w_eco1237, !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1238(w_eco1238, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1239(w_eco1239, !sel_prim[0], !sel_prim[2], !sel_prim[7], sel_prim[3]);
	and _ECO_1240(w_eco1240, sel_prim[0], sel_prim[12], !sel_prim[7], !sel_prim[10], sel_prim[3]);
	and _ECO_1241(w_eco1241, sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1242(w_eco1242, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[13], sel_prim[3]);
	and _ECO_1243(w_eco1243, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[3]);
	and _ECO_1244(w_eco1244, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1245(w_eco1245, sel_prim[0], sel_prim[12], !sel_prim[7], sel_prim[9], sel_prim[3]);
	and _ECO_1246(w_eco1246, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[13], sel_prim[3]);
	and _ECO_1247(w_eco1247, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[14], sel_prim[3]);
	and _ECO_1248(w_eco1248, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1249(w_eco1249, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1250(w_eco1250, sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_1251(w_eco1251, !sel_prim[0], sel_prim[1], !sel_prim[7], sel_prim[3]);
	and _ECO_1252(w_eco1252, sel_prim[0], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[9], sel_prim[3]);
	and _ECO_1253(w_eco1253, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[14], sel_prim[3]);
	and _ECO_1254(w_eco1254, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1255(w_eco1255, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[3]);
	and _ECO_1256(w_eco1256, sel_prim[0], sel_prim[14], !sel_prim[7], !sel_prim[10], sel_prim[3]);
	and _ECO_1257(w_eco1257, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1258(w_eco1258, sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5]);
	and _ECO_1259(w_eco1259, sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1260(w_eco1260, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[3]);
	and _ECO_1261(w_eco1261, sel_prim[0], sel_prim[14], !sel_prim[7], sel_prim[9], sel_prim[3]);
	and _ECO_1262(w_eco1262, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[4], !sel_prim[17]);
	and _ECO_1263(w_eco1263, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1264(w_eco1264, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], sel_prim[4]);
	and _ECO_1265(w_eco1265, !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1266(w_eco1266, !sel_prim[16], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1267(w_eco1267, sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1268(w_eco1268, !sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1269(w_eco1269, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4], !sel_prim[17]);
	and _ECO_1270(w_eco1270, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], sel_prim[4]);
	and _ECO_1271(w_eco1271, !sel_prim[16], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1272(w_eco1272, !sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1273(w_eco1273, !sel_prim[15], !sel_prim[16], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1274(w_eco1274, !sel_prim[12], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1275(w_eco1275, !sel_prim[15], !sel_prim[16], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1276(w_eco1276, !sel_prim[15], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	or _ECO_1277(w_eco1277, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276);
	xor _ECO_out16(prim_out[28], sub_wire16, w_eco1277);
	and _ECO_1278(w_eco1278, sel_prim[0], sel_prim[11], sel_prim[8], sel_prim[3]);
	and _ECO_1279(w_eco1279, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1280(w_eco1280, sel_prim[0], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1281(w_eco1281, !sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1282(w_eco1282, !sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[3]);
	and _ECO_1283(w_eco1283, sel_prim[0], sel_prim[11], sel_prim[8], !sel_prim[4]);
	and _ECO_1284(w_eco1284, sel_prim[0], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1285(w_eco1285, sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[4]);
	and _ECO_1286(w_eco1286, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1287(w_eco1287, sel_prim[0], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_1288(w_eco1288, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_1289(w_eco1289, sel_prim[0], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4]);
	and _ECO_1290(w_eco1290, !sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1291(w_eco1291, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1292(w_eco1292, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1293(w_eco1293, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[4]);
	and _ECO_1294(w_eco1294, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1295(w_eco1295, sel_prim[0], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1296(w_eco1296, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1297(w_eco1297, sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1298(w_eco1298, sel_prim[0], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1299(w_eco1299, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1300(w_eco1300, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1301(w_eco1301, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[4], sel_prim[5]);
	and _ECO_1302(w_eco1302, sel_prim[1], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1303(w_eco1303, sel_prim[0], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1304(w_eco1304, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1305(w_eco1305, !sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1306(w_eco1306, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1307(w_eco1307, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1308(w_eco1308, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1309(w_eco1309, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1310(w_eco1310, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1311(w_eco1311, !sel_prim[0], sel_prim[15], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1312(w_eco1312, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1313(w_eco1313, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1314(w_eco1314, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1315(w_eco1315, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1316(w_eco1316, !sel_prim[0], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1317(w_eco1317, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5]);
	and _ECO_1318(w_eco1318, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1319(w_eco1319, !sel_prim[0], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1320(w_eco1320, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1321(w_eco1321, !sel_prim[0], sel_prim[15], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5]);
	and _ECO_1322(w_eco1322, !sel_prim[0], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1323(w_eco1323, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1324(w_eco1324, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1325(w_eco1325, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	and _ECO_1326(w_eco1326, !sel_prim[0], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], !sel_prim[18]);
	and _ECO_1327(w_eco1327, !sel_prim[0], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], !sel_prim[5], sel_prim[17]);
	or _ECO_1328(w_eco1328, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327);
	xor _ECO_out17(prim_out[24], sub_wire17, w_eco1328);
	and _ECO_1329(w_eco1329, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1330(w_eco1330, sel_prim[0], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1331(w_eco1331, sel_prim[0], !sel_prim[7], !sel_prim[8]);
	and _ECO_1332(w_eco1332, !sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1333(w_eco1333, sel_prim[0], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1334(w_eco1334, sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1335(w_eco1335, sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1336(w_eco1336, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1337(w_eco1337, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_1338(w_eco1338, sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1339(w_eco1339, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8]);
	and _ECO_1340(w_eco1340, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[3]);
	and _ECO_1341(w_eco1341, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1342(w_eco1342, sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], sel_prim[5]);
	and _ECO_1343(w_eco1343, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[4], sel_prim[5]);
	and _ECO_1344(w_eco1344, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[4], sel_prim[6]);
	and _ECO_1345(w_eco1345, !sel_prim[11], sel_prim[7], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1346(w_eco1346, !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[8], sel_prim[3]);
	and _ECO_1347(w_eco1347, sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1348(w_eco1348, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1349(w_eco1349, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[8]);
	and _ECO_1350(w_eco1350, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[5]);
	and _ECO_1351(w_eco1351, sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[6]);
	and _ECO_1352(w_eco1352, sel_prim[0], !sel_prim[11], sel_prim[7]);
	and _ECO_1353(w_eco1353, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1354(w_eco1354, sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1355(w_eco1355, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_1356(w_eco1356, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1357(w_eco1357, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[5]);
	and _ECO_1358(w_eco1358, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[10], !sel_prim[3], sel_prim[5]);
	and _ECO_1359(w_eco1359, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1360(w_eco1360, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_1361(w_eco1361, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[4], sel_prim[6]);
	and _ECO_1362(w_eco1362, sel_prim[2], !sel_prim[11], sel_prim[7], !sel_prim[4], !sel_prim[5]);
	and _ECO_1363(w_eco1363, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1364(w_eco1364, !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1365(w_eco1365, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[5]);
	and _ECO_1366(w_eco1366, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[5]);
	and _ECO_1367(w_eco1367, sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1368(w_eco1368, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[4], sel_prim[5]);
	and _ECO_1369(w_eco1369, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[5]);
	and _ECO_1370(w_eco1370, !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[5], sel_prim[6]);
	and _ECO_1371(w_eco1371, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_1372(w_eco1372, sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_1373(w_eco1373, sel_prim[1], !sel_prim[11], sel_prim[7], !sel_prim[4], !sel_prim[5]);
	and _ECO_1374(w_eco1374, !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1375(w_eco1375, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[5]);
	and _ECO_1376(w_eco1376, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[10], !sel_prim[3], sel_prim[5]);
	and _ECO_1377(w_eco1377, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[6]);
	and _ECO_1378(w_eco1378, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1379(w_eco1379, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[9], !sel_prim[3], sel_prim[5]);
	and _ECO_1380(w_eco1380, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1381(w_eco1381, !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5]);
	or _ECO_1382(w_eco1382, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381);
	xor _ECO_out18(prim_out[16], sub_wire18, w_eco1382);
	and _ECO_1383(w_eco1383, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7]);
	and _ECO_1384(w_eco1384, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1385(w_eco1385, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1386(w_eco1386, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1387(w_eco1387, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1388(w_eco1388, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1389(w_eco1389, !sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1390(w_eco1390, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1391(w_eco1391, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1392(w_eco1392, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1393(w_eco1393, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1394(w_eco1394, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1395(w_eco1395, !sel_prim[0], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1396(w_eco1396, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1397(w_eco1397, !sel_prim[0], !sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1398(w_eco1398, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1399(w_eco1399, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1400(w_eco1400, !sel_prim[0], !sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1401(w_eco1401, !sel_prim[0], !sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1402(w_eco1402, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1403(w_eco1403, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1404(w_eco1404, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], sel_prim[3]);
	and _ECO_1405(w_eco1405, !sel_prim[0], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], !sel_prim[18]);
	and _ECO_1406(w_eco1406, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1407(w_eco1407, !sel_prim[0], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1408(w_eco1408, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1409(w_eco1409, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1410(w_eco1410, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1411(w_eco1411, !sel_prim[0], !sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[6]);
	and _ECO_1412(w_eco1412, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1413(w_eco1413, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], !sel_prim[6]);
	and _ECO_1414(w_eco1414, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1415(w_eco1415, !sel_prim[0], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_1416(w_eco1416, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1417(w_eco1417, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1418(w_eco1418, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1419(w_eco1419, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_1420(w_eco1420, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_1421(w_eco1421, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1422(w_eco1422, !sel_prim[0], !sel_prim[15], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[18]);
	and _ECO_1423(w_eco1423, !sel_prim[0], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1424(w_eco1424, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1425(w_eco1425, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1426(w_eco1426, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1427(w_eco1427, !sel_prim[0], !sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5]);
	and _ECO_1428(w_eco1428, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1429(w_eco1429, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1430(w_eco1430, !sel_prim[0], !sel_prim[15], !sel_prim[16], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], sel_prim[17]);
	and _ECO_1431(w_eco1431, !sel_prim[0], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_1432(w_eco1432, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1433(w_eco1433, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_1434(w_eco1434, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5], !sel_prim[6], !sel_prim[18]);
	and _ECO_1435(w_eco1435, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1436(w_eco1436, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[4], sel_prim[6]);
	and _ECO_1437(w_eco1437, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[5], !sel_prim[6], sel_prim[17]);
	and _ECO_1438(w_eco1438, !sel_prim[0], !sel_prim[15], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_1439(w_eco1439, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_1440(w_eco1440, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[12], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1441(w_eco1441, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_1442(w_eco1442, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1443(w_eco1443, !sel_prim[0], !sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	or _ECO_1444(w_eco1444, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443);
	xor _ECO_out19(prim_out[13], sub_wire19, w_eco1444);
	and _ECO_1445(w_eco1445, !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1446(w_eco1446, !sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[3]);
	assign w_eco1447 = sel_prim[0];
	and _ECO_1448(w_eco1448, !sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[4]);
	and _ECO_1449(w_eco1449, !sel_prim[15], sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1450(w_eco1450, sel_prim[2], !sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1451(w_eco1451, !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1452(w_eco1452, !sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[5]);
	and _ECO_1453(w_eco1453, sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[5]);
	and _ECO_1454(w_eco1454, sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_1455(w_eco1455, sel_prim[11], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1456(w_eco1456, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1457(w_eco1457, sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1458(w_eco1458, !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1459(w_eco1459, sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1460(w_eco1460, sel_prim[2], !sel_prim[15], sel_prim[11], sel_prim[5]);
	and _ECO_1461(w_eco1461, sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[5]);
	and _ECO_1462(w_eco1462, !sel_prim[15], sel_prim[11], sel_prim[8], sel_prim[6]);
	and _ECO_1463(w_eco1463, sel_prim[2], sel_prim[11], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1464(w_eco1464, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1465(w_eco1465, sel_prim[1], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_1466(w_eco1466, !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1467(w_eco1467, sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], sel_prim[4]);
	and _ECO_1468(w_eco1468, sel_prim[11], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1469(w_eco1469, !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1470(w_eco1470, sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[4]);
	and _ECO_1471(w_eco1471, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[5]);
	and _ECO_1472(w_eco1472, !sel_prim[15], sel_prim[11], sel_prim[7], sel_prim[6]);
	and _ECO_1473(w_eco1473, sel_prim[2], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1474(w_eco1474, sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[3]);
	and _ECO_1475(w_eco1475, !sel_prim[15], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_1476(w_eco1476, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[5]);
	and _ECO_1477(w_eco1477, sel_prim[1], !sel_prim[15], sel_prim[11], sel_prim[5]);
	and _ECO_1478(w_eco1478, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[4]);
	and _ECO_1479(w_eco1479, !sel_prim[1], !sel_prim[2], sel_prim[11], sel_prim[7], sel_prim[6]);
	and _ECO_1480(w_eco1480, !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1481(w_eco1481, !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1482(w_eco1482, sel_prim[1], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1483(w_eco1483, sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[5], !sel_prim[6]);
	and _ECO_1484(w_eco1484, !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], sel_prim[3]);
	and _ECO_1485(w_eco1485, !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1486(w_eco1486, sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1487(w_eco1487, sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[4]);
	and _ECO_1488(w_eco1488, sel_prim[11], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1489(w_eco1489, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1490(w_eco1490, sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], sel_prim[5]);
	and _ECO_1491(w_eco1491, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[4]);
	and _ECO_1492(w_eco1492, sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3], sel_prim[5]);
	and _ECO_1493(w_eco1493, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], sel_prim[7], !sel_prim[4]);
	and _ECO_1494(w_eco1494, sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[5], !sel_prim[6]);
	and _ECO_1495(w_eco1495, sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[5], !sel_prim[6]);
	and _ECO_1496(w_eco1496, sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_1497(w_eco1497, !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1498(w_eco1498, sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], sel_prim[5]);
	and _ECO_1499(w_eco1499, sel_prim[1], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3], sel_prim[5]);
	and _ECO_1500(w_eco1500, sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[5]);
	and _ECO_1501(w_eco1501, sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1502(w_eco1502, sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[5], !sel_prim[6]);
	and _ECO_1503(w_eco1503, sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_1504(w_eco1504, !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1505(w_eco1505, sel_prim[2], !sel_prim[15], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[6], !sel_prim[17]);
	and _ECO_1506(w_eco1506, sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[6]);
	and _ECO_1507(w_eco1507, sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1508(w_eco1508, sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_1509(w_eco1509, sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[5]);
	and _ECO_1510(w_eco1510, sel_prim[1], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[5]);
	and _ECO_1511(w_eco1511, sel_prim[2], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[6]);
	and _ECO_1512(w_eco1512, sel_prim[1], !sel_prim[15], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[6], !sel_prim[17]);
	and _ECO_1513(w_eco1513, sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	and _ECO_1514(w_eco1514, sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[6]);
	and _ECO_1515(w_eco1515, sel_prim[2], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1516(w_eco1516, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1517(w_eco1517, sel_prim[1], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[6]);
	and _ECO_1518(w_eco1518, sel_prim[1], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[5]);
	and _ECO_1519(w_eco1519, sel_prim[1], !sel_prim[15], sel_prim[16], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[6]);
	and _ECO_1520(w_eco1520, sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[6]);
	and _ECO_1521(w_eco1521, sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[6], !sel_prim[17]);
	and _ECO_1522(w_eco1522, sel_prim[1], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1523(w_eco1523, !sel_prim[15], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1524(w_eco1524, sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[6]);
	and _ECO_1525(w_eco1525, sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[6], !sel_prim[17]);
	and _ECO_1526(w_eco1526, !sel_prim[15], sel_prim[16], !sel_prim[13], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1527(w_eco1527, sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[6]);
	and _ECO_1528(w_eco1528, sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1529(w_eco1529, sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	and _ECO_1530(w_eco1530, sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1531(w_eco1531, sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[3], !sel_prim[4], !sel_prim[5], !sel_prim[6]);
	or _ECO_1532(w_eco1532, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531);
	xor _ECO_out20(prim_out[20], sub_wire20, w_eco1532);
	and _ECO_1533(w_eco1533, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1534(w_eco1534, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1535(w_eco1535, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[3]);
	and _ECO_1536(w_eco1536, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[5]);
	and _ECO_1537(w_eco1537, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], sel_prim[3]);
	and _ECO_1538(w_eco1538, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[7]);
	and _ECO_1539(w_eco1539, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1540(w_eco1540, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[5]);
	and _ECO_1541(w_eco1541, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11]);
	and _ECO_1542(w_eco1542, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1543(w_eco1543, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[8], sel_prim[10]);
	and _ECO_1544(w_eco1544, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1545(w_eco1545, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1546(w_eco1546, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_1547(w_eco1547, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[4], sel_prim[5]);
	and _ECO_1548(w_eco1548, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[7]);
	and _ECO_1549(w_eco1549, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[8], !sel_prim[10]);
	and _ECO_1550(w_eco1550, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[8], sel_prim[9]);
	and _ECO_1551(w_eco1551, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1552(w_eco1552, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1553(w_eco1553, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1554(w_eco1554, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1555(w_eco1555, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[6]);
	and _ECO_1556(w_eco1556, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1557(w_eco1557, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1558(w_eco1558, !sel_prim[0], sel_prim[2], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1559(w_eco1559, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1560(w_eco1560, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14]);
	and _ECO_1561(w_eco1561, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1562(w_eco1562, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1563(w_eco1563, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1564(w_eco1564, !sel_prim[0], sel_prim[1], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], sel_prim[4]);
	and _ECO_1565(w_eco1565, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14]);
	and _ECO_1566(w_eco1566, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1567(w_eco1567, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[4], sel_prim[6]);
	and _ECO_1568(w_eco1568, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1569(w_eco1569, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1570(w_eco1570, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1571(w_eco1571, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1572(w_eco1572, !sel_prim[0], sel_prim[2], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1573(w_eco1573, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1574(w_eco1574, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[4], sel_prim[6]);
	and _ECO_1575(w_eco1575, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1576(w_eco1576, !sel_prim[0], sel_prim[2], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1577(w_eco1577, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1578(w_eco1578, !sel_prim[0], sel_prim[1], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1579(w_eco1579, !sel_prim[0], sel_prim[1], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1580(w_eco1580, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1581(w_eco1581, !sel_prim[0], sel_prim[2], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1582(w_eco1582, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1583(w_eco1583, !sel_prim[0], sel_prim[1], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_1584(w_eco1584, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583);
	xor _ECO_out21(prim_out[21], sub_wire21, w_eco1584);
	and _ECO_1585(w_eco1585, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1586(w_eco1586, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1587(w_eco1587, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], !sel_prim[8]);
	and _ECO_1588(w_eco1588, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1589(w_eco1589, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1590(w_eco1590, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1591(w_eco1591, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1592(w_eco1592, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[7]);
	and _ECO_1593(w_eco1593, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_1594(w_eco1594, !sel_prim[0], !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_1595(w_eco1595, !sel_prim[0], !sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8]);
	and _ECO_1596(w_eco1596, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[11], !sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1597(w_eco1597, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8]);
	and _ECO_1598(w_eco1598, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1599(w_eco1599, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1600(w_eco1600, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1601(w_eco1601, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7]);
	and _ECO_1602(w_eco1602, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8]);
	and _ECO_1603(w_eco1603, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[17]);
	and _ECO_1604(w_eco1604, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1605(w_eco1605, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8]);
	and _ECO_1606(w_eco1606, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1607(w_eco1607, !sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1608(w_eco1608, !sel_prim[0], !sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[5]);
	and _ECO_1609(w_eco1609, !sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1610(w_eco1610, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1611(w_eco1611, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7]);
	and _ECO_1612(w_eco1612, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1613(w_eco1613, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[7]);
	and _ECO_1614(w_eco1614, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1615(w_eco1615, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1616(w_eco1616, !sel_prim[0], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[9], sel_prim[10], sel_prim[3]);
	and _ECO_1617(w_eco1617, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1618(w_eco1618, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[9]);
	and _ECO_1619(w_eco1619, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1620(w_eco1620, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1621(w_eco1621, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1622(w_eco1622, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1623(w_eco1623, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1624(w_eco1624, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1625(w_eco1625, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1626(w_eco1626, !sel_prim[0], !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1627(w_eco1627, !sel_prim[0], sel_prim[15], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1628(w_eco1628, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[4], !sel_prim[5], sel_prim[6]);
	and _ECO_1629(w_eco1629, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1630(w_eco1630, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1631(w_eco1631, !sel_prim[0], !sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1632(w_eco1632, !sel_prim[0], !sel_prim[1], sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1633(w_eco1633, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_1634(w_eco1634, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633);
	xor _ECO_out22(prim_out[29], sub_wire22, w_eco1634);
	and _ECO_1635(w_eco1635, !sel_prim[0], sel_prim[11], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1636(w_eco1636, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7]);
	and _ECO_1637(w_eco1637, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[3]);
	and _ECO_1638(w_eco1638, !sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1639(w_eco1639, !sel_prim[0], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1640(w_eco1640, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1641(w_eco1641, !sel_prim[0], sel_prim[11], !sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1642(w_eco1642, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8]);
	and _ECO_1643(w_eco1643, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[7]);
	and _ECO_1644(w_eco1644, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1645(w_eco1645, !sel_prim[0], sel_prim[1], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3]);
	and _ECO_1646(w_eco1646, !sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1647(w_eco1647, sel_prim[0], !sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1648(w_eco1648, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1649(w_eco1649, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], sel_prim[4]);
	and _ECO_1650(w_eco1650, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_1651(w_eco1651, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1652(w_eco1652, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1653(w_eco1653, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3]);
	and _ECO_1654(w_eco1654, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1655(w_eco1655, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8]);
	and _ECO_1656(w_eco1656, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_1657(w_eco1657, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1658(w_eco1658, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1659(w_eco1659, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[3], sel_prim[4], sel_prim[18]);
	and _ECO_1660(w_eco1660, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[3]);
	and _ECO_1661(w_eco1661, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1662(w_eco1662, !sel_prim[0], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[5]);
	and _ECO_1663(w_eco1663, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1664(w_eco1664, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1665(w_eco1665, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[17]);
	and _ECO_1666(w_eco1666, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1667(w_eco1667, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[3]);
	and _ECO_1668(w_eco1668, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[3]);
	and _ECO_1669(w_eco1669, sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[12], !sel_prim[13], sel_prim[14], sel_prim[7], !sel_prim[3]);
	and _ECO_1670(w_eco1670, !sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1671(w_eco1671, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1672(w_eco1672, !sel_prim[0], sel_prim[2], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7]);
	and _ECO_1673(w_eco1673, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[17]);
	and _ECO_1674(w_eco1674, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3]);
	and _ECO_1675(w_eco1675, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], !sel_prim[7], !sel_prim[3]);
	and _ECO_1676(w_eco1676, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[12], sel_prim[14], sel_prim[7], !sel_prim[3]);
	and _ECO_1677(w_eco1677, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[8], !sel_prim[3], !sel_prim[5]);
	and _ECO_1678(w_eco1678, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1679(w_eco1679, !sel_prim[0], sel_prim[1], sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7]);
	and _ECO_1680(w_eco1680, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[10]);
	and _ECO_1681(w_eco1681, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[17]);
	and _ECO_1682(w_eco1682, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7], !sel_prim[3], !sel_prim[5]);
	and _ECO_1683(w_eco1683, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1684(w_eco1684, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1685(w_eco1685, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[7], !sel_prim[3]);
	and _ECO_1686(w_eco1686, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[17]);
	and _ECO_1687(w_eco1687, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[18]);
	and _ECO_1688(w_eco1688, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[7], !sel_prim[3]);
	and _ECO_1689(w_eco1689, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[18]);
	and _ECO_1690(w_eco1690, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[18]);
	and _ECO_1691(w_eco1691, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[7], !sel_prim[3], sel_prim[18]);
	or _ECO_1692(w_eco1692, w_eco1635, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691);
	xor _ECO_out23(prim_out[7], sub_wire23, w_eco1692);
	and _ECO_1693(w_eco1693, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1694(w_eco1694, !sel_prim[0], sel_prim[15], sel_prim[11], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1695(w_eco1695, !sel_prim[0], !sel_prim[15], sel_prim[11], !sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1696(w_eco1696, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[3]);
	and _ECO_1697(w_eco1697, !sel_prim[0], sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1698(w_eco1698, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[7]);
	and _ECO_1699(w_eco1699, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7]);
	and _ECO_1700(w_eco1700, !sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1701(w_eco1701, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[3]);
	and _ECO_1702(w_eco1702, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[4]);
	and _ECO_1703(w_eco1703, !sel_prim[0], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1704(w_eco1704, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[10], sel_prim[4]);
	and _ECO_1705(w_eco1705, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[12], sel_prim[7], sel_prim[4]);
	and _ECO_1706(w_eco1706, !sel_prim[0], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1707(w_eco1707, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1708(w_eco1708, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1709(w_eco1709, !sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1710(w_eco1710, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[5]);
	and _ECO_1711(w_eco1711, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3]);
	and _ECO_1712(w_eco1712, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1713(w_eco1713, !sel_prim[0], sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1714(w_eco1714, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1715(w_eco1715, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1716(w_eco1716, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[9], sel_prim[4]);
	and _ECO_1717(w_eco1717, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], sel_prim[7], sel_prim[4]);
	and _ECO_1718(w_eco1718, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1719(w_eco1719, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[4]);
	and _ECO_1720(w_eco1720, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[12], !sel_prim[8], sel_prim[10], sel_prim[4]);
	and _ECO_1721(w_eco1721, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1722(w_eco1722, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1723(w_eco1723, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1724(w_eco1724, !sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1725(w_eco1725, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[5], !sel_prim[6]);
	and _ECO_1726(w_eco1726, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8]);
	and _ECO_1727(w_eco1727, !sel_prim[0], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10], sel_prim[3]);
	and _ECO_1728(w_eco1728, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1729(w_eco1729, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[4]);
	and _ECO_1730(w_eco1730, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1731(w_eco1731, !sel_prim[0], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1732(w_eco1732, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1733(w_eco1733, !sel_prim[0], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1734(w_eco1734, !sel_prim[0], !sel_prim[1], sel_prim[2], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1735(w_eco1735, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[7]);
	and _ECO_1736(w_eco1736, !sel_prim[0], !sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[3], !sel_prim[5]);
	and _ECO_1737(w_eco1737, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[10], !sel_prim[5], !sel_prim[6]);
	and _ECO_1738(w_eco1738, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[5], !sel_prim[6]);
	and _ECO_1739(w_eco1739, !sel_prim[0], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1740(w_eco1740, !sel_prim[0], sel_prim[2], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1741(w_eco1741, !sel_prim[0], sel_prim[15], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1742(w_eco1742, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1743(w_eco1743, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1744(w_eco1744, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_1745(w_eco1745, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], !sel_prim[8], sel_prim[10], sel_prim[4]);
	and _ECO_1746(w_eco1746, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1747(w_eco1747, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[3], sel_prim[4]);
	and _ECO_1748(w_eco1748, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1749(w_eco1749, !sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1750(w_eco1750, !sel_prim[0], sel_prim[15], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1751(w_eco1751, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[9], !sel_prim[5], !sel_prim[6]);
	and _ECO_1752(w_eco1752, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[5], !sel_prim[6]);
	and _ECO_1753(w_eco1753, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1754(w_eco1754, !sel_prim[0], sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[5], !sel_prim[6]);
	and _ECO_1755(w_eco1755, !sel_prim[0], sel_prim[1], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1756(w_eco1756, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1757(w_eco1757, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[13], !sel_prim[7], sel_prim[3]);
	and _ECO_1758(w_eco1758, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1759(w_eco1759, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[10]);
	and _ECO_1760(w_eco1760, !sel_prim[0], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1761(w_eco1761, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_1762(w_eco1762, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_1763(w_eco1763, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[3], sel_prim[4], !sel_prim[17]);
	and _ECO_1764(w_eco1764, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[5], !sel_prim[6]);
	and _ECO_1765(w_eco1765, !sel_prim[0], sel_prim[2], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1766(w_eco1766, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1767(w_eco1767, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1768(w_eco1768, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1769(w_eco1769, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[8], sel_prim[10], sel_prim[3]);
	and _ECO_1770(w_eco1770, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], sel_prim[4]);
	and _ECO_1771(w_eco1771, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[3], sel_prim[4]);
	and _ECO_1772(w_eco1772, !sel_prim[0], sel_prim[1], !sel_prim[8], sel_prim[9], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1773(w_eco1773, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1774(w_eco1774, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1775(w_eco1775, !sel_prim[0], sel_prim[2], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1776(w_eco1776, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17]);
	and _ECO_1777(w_eco1777, !sel_prim[0], sel_prim[1], !sel_prim[15], sel_prim[16], !sel_prim[11], !sel_prim[13], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	or _ECO_1778(w_eco1778, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777);
	xor _ECO_out24(prim_out[14], sub_wire24, w_eco1778);
	and _ECO_1779(w_eco1779, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1780(w_eco1780, !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1781(w_eco1781, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1782(w_eco1782, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1783(w_eco1783, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1784(w_eco1784, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1785(w_eco1785, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1786(w_eco1786, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1787(w_eco1787, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1788(w_eco1788, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1789(w_eco1789, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1790(w_eco1790, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], sel_prim[3]);
	and _ECO_1791(w_eco1791, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1792(w_eco1792, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1793(w_eco1793, sel_prim[0], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1794(w_eco1794, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1795(w_eco1795, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1796(w_eco1796, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1797(w_eco1797, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1798(w_eco1798, sel_prim[0], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1799(w_eco1799, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1800(w_eco1800, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1801(w_eco1801, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1802(w_eco1802, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1803(w_eco1803, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1804(w_eco1804, !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1805(w_eco1805, !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1806(w_eco1806, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1807(w_eco1807, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[11], !sel_prim[13], !sel_prim[14], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	or _ECO_1808(w_eco1808, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807);
	xor _ECO_out25(prim_out[15], sub_wire25, w_eco1808);
	and _ECO_1809(w_eco1809, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1810(w_eco1810, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[8], sel_prim[3]);
	and _ECO_1811(w_eco1811, sel_prim[0], !sel_prim[11], sel_prim[7], sel_prim[3]);
	and _ECO_1812(w_eco1812, !sel_prim[0], sel_prim[15], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1813(w_eco1813, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], sel_prim[3]);
	and _ECO_1814(w_eco1814, sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[8], sel_prim[3]);
	and _ECO_1815(w_eco1815, sel_prim[2], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_1816(w_eco1816, !sel_prim[0], sel_prim[11], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1817(w_eco1817, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[5]);
	and _ECO_1818(w_eco1818, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1819(w_eco1819, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1820(w_eco1820, !sel_prim[0], !sel_prim[1], !sel_prim[2], sel_prim[11], !sel_prim[7], sel_prim[8]);
	and _ECO_1821(w_eco1821, sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], sel_prim[8], sel_prim[3]);
	and _ECO_1822(w_eco1822, sel_prim[1], !sel_prim[11], sel_prim[12], sel_prim[7], sel_prim[3]);
	and _ECO_1823(w_eco1823, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[8]);
	and _ECO_1824(w_eco1824, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1825(w_eco1825, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[8], sel_prim[3]);
	and _ECO_1826(w_eco1826, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_1827(w_eco1827, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1828(w_eco1828, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[5]);
	and _ECO_1829(w_eco1829, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1830(w_eco1830, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1831(w_eco1831, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[6]);
	and _ECO_1832(w_eco1832, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1833(w_eco1833, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], sel_prim[7]);
	and _ECO_1834(w_eco1834, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1835(w_eco1835, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1836(w_eco1836, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[7], !sel_prim[3], sel_prim[4]);
	and _ECO_1837(w_eco1837, !sel_prim[0], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], sel_prim[8], !sel_prim[3]);
	and _ECO_1838(w_eco1838, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1839(w_eco1839, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1840(w_eco1840, sel_prim[2], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1841(w_eco1841, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1842(w_eco1842, !sel_prim[0], sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1843(w_eco1843, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[4], sel_prim[6]);
	and _ECO_1844(w_eco1844, sel_prim[0], !sel_prim[11], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1845(w_eco1845, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1846(w_eco1846, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[7], !sel_prim[8], !sel_prim[9], sel_prim[10]);
	and _ECO_1847(w_eco1847, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1848(w_eco1848, sel_prim[2], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1849(w_eco1849, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1850(w_eco1850, !sel_prim[0], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9], sel_prim[3]);
	and _ECO_1851(w_eco1851, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[11], !sel_prim[7], !sel_prim[9], !sel_prim[10]);
	and _ECO_1852(w_eco1852, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[4]);
	and _ECO_1853(w_eco1853, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1854(w_eco1854, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1855(w_eco1855, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1856(w_eco1856, !sel_prim[0], sel_prim[1], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1857(w_eco1857, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1858(w_eco1858, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1859(w_eco1859, !sel_prim[0], sel_prim[15], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1860(w_eco1860, sel_prim[1], !sel_prim[15], !sel_prim[11], !sel_prim[13], sel_prim[14], sel_prim[7], sel_prim[3]);
	and _ECO_1861(w_eco1861, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1862(w_eco1862, !sel_prim[0], sel_prim[2], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[17], !sel_prim[18]);
	and _ECO_1863(w_eco1863, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4]);
	and _ECO_1864(w_eco1864, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_1865(w_eco1865, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1866(w_eco1866, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1867(w_eco1867, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[4], sel_prim[6]);
	and _ECO_1868(w_eco1868, sel_prim[1], !sel_prim[15], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1869(w_eco1869, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[12], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1870(w_eco1870, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1871(w_eco1871, sel_prim[0], !sel_prim[11], !sel_prim[13], sel_prim[7], !sel_prim[4], sel_prim[5]);
	and _ECO_1872(w_eco1872, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], sel_prim[7], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1873(w_eco1873, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1874(w_eco1874, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[3]);
	and _ECO_1875(w_eco1875, !sel_prim[0], sel_prim[1], !sel_prim[15], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], sel_prim[8], !sel_prim[17], !sel_prim[18]);
	and _ECO_1876(w_eco1876, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1877(w_eco1877, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], sel_prim[13], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10]);
	and _ECO_1878(w_eco1878, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[18]);
	and _ECO_1879(w_eco1879, !sel_prim[0], !sel_prim[1], !sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[13], !sel_prim[14], !sel_prim[7], !sel_prim[8], sel_prim[9]);
	and _ECO_1880(w_eco1880, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1881(w_eco1881, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1882(w_eco1882, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[7], !sel_prim[9], sel_prim[10], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1883(w_eco1883, !sel_prim[0], sel_prim[2], sel_prim[15], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1884(w_eco1884, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1885(w_eco1885, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[3]);
	and _ECO_1886(w_eco1886, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_1887(w_eco1887, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[17]);
	and _ECO_1888(w_eco1888, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[18]);
	and _ECO_1889(w_eco1889, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1890(w_eco1890, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[6]);
	and _ECO_1891(w_eco1891, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1892(w_eco1892, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1893(w_eco1893, !sel_prim[0], sel_prim[2], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1894(w_eco1894, !sel_prim[0], sel_prim[2], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1895(w_eco1895, !sel_prim[0], sel_prim[1], sel_prim[15], sel_prim[7], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1896(w_eco1896, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1897(w_eco1897, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1898(w_eco1898, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6]);
	and _ECO_1899(w_eco1899, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], sel_prim[4], !sel_prim[17], !sel_prim[18]);
	and _ECO_1900(w_eco1900, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], sel_prim[8], !sel_prim[3], sel_prim[17]);
	and _ECO_1901(w_eco1901, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_1902(w_eco1902, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[6]);
	and _ECO_1903(w_eco1903, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1904(w_eco1904, !sel_prim[0], sel_prim[1], !sel_prim[7], sel_prim[8], !sel_prim[3], !sel_prim[4], sel_prim[5]);
	and _ECO_1905(w_eco1905, !sel_prim[0], sel_prim[1], sel_prim[15], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[4], sel_prim[5]);
	and _ECO_1906(w_eco1906, !sel_prim[0], sel_prim[2], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1907(w_eco1907, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[5]);
	and _ECO_1908(w_eco1908, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_1909(w_eco1909, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[18]);
	and _ECO_1910(w_eco1910, !sel_prim[0], sel_prim[1], !sel_prim[11], !sel_prim[12], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], !sel_prim[4], sel_prim[6]);
	and _ECO_1911(w_eco1911, !sel_prim[0], sel_prim[2], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	and _ECO_1912(w_eco1912, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], !sel_prim[12], !sel_prim[14], !sel_prim[7], !sel_prim[8], !sel_prim[9], !sel_prim[10], sel_prim[17]);
	and _ECO_1913(w_eco1913, !sel_prim[0], sel_prim[1], !sel_prim[16], !sel_prim[11], sel_prim[12], !sel_prim[7], !sel_prim[9], !sel_prim[10], !sel_prim[3], !sel_prim[5], !sel_prim[6], !sel_prim[17], !sel_prim[18]);
	or _ECO_1914(w_eco1914, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913);
	xor _ECO_out26(prim_out[6], sub_wire26, w_eco1914);

endmodule