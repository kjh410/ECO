module ex5 (y,a,b,cin,cout);
	input [4:0] a,b;
	input cin;
	output cout;
	output [4:0] y;
	wire [24:0] w;
	
	xor xor_0 (w[0],a[4],b[4]);
	and and_0 (w[1],a[4],b[4]);
	xor xor_1 (w[2],w[0],cin);
	and and_1 (w[3],w[0],cin);
	or or_0 (w[4],w[3],w[1]);
	assign y[4]= w[2];
	xor xor_00(w[5],a[3],b[3]);
	and and_00(w[6],a[3],b[3]);
	xor xor_11(w[7],w[5],w[4]);
	and and_11(w[8],w[5],w[4]);
	or or_11(w[9],w[8],w[6]);
	assign y[3] = w[7];
	xor xor_000(w[10],a[2],b[2]);
	and and_000(w[11],a[2],b[2]);
	xor xor_111(w[12],w[10],w[9]);
	and and_111(w[13],w[10],w[9]);
	or or_111(w[14],w[13],w[11]);
	assign y[2] = w[12];
	xor xor_0000(w[15],a[1],b[1]);
	and and_0000(w[16],a[1],b[1]);
	xor xor_1111(w[17],w[15],w[14]);
	and and_1111(w[18],w[15],w[14]);
	or or_1111(w[19],w[18],w[16]);
	assign y[1] = w[17];
	or xor_00000(w[20],a[0],b[0]);
	and and_00000(w[21],a[0],b[0]);
	xor xor_11111(w[22],w[20],w[19]);
	and and_11111(w[23],w[20],w[19]);
	or or_11111(w[24],w[23],w[21]);
	assign y[0] = w[22];
	assign cout = w[24];
endmodule
