module top(a_gtet_b,a,b);
	input [7:0]a, b;
	output a_gtet_b;
	wire [7:0]a, b;
	wire a_gtet_b, n_8, n_13, n_43, n_52, n_59, n_64, n_67, n_149, n_156, n_158, n_171, n_403, n_407, n_410, n_415, n_425, n_432, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988;

	nand g47(n_52, n_8, a[2]);
	nand g58(n_149, n_485, n_496);
	nor g133(n_158, n_43, a[1]);
	not g468(n_442, a[2]);
	not g469(n_443, a[1]);
	not g470(n_444, b[2]);
	not g471(n_445, b[5]);
	not g472(n_446, a[5]);
	not g473(n_447, b[7]);
	not g474(n_448, a[7]);
	not g475(n_449, a[3]);
	not g476(n_450, b[4]);
	not g477(n_451, a[4]);
	not g478(n_452, b[6]);
	not g479(n_453, a[6]);
	not g480(n_454, b[1]);
	not g481(n_455, a[0]);
	nand g482(n_8, n_449, b[3]);
	not g483(n_456, n_8);
	nand g484(n_13, a[7], n_447);
	not g485(n_457, n_13);
	nor g486(n_458, a[6], n_452);
	not g487(n_459, n_458);
	nor g488(n_407, n_442, b[2]);
	not g489(n_460, n_407);
	nor g490(n_43, n_449, b[3]);
	not g491(n_461, n_43);
	not g492(n_462, n_158);
	nor g493(n_463, n_43, n_454);
	not g494(n_464, n_463);
	nand g495(n_465, n_462, n_464);
	nand g496(n_466, n_460, n_465, b[0]);
	nor g497(n_403, a[2], n_444);
	not g498(n_467, n_403);
	nand g499(n_410, n_467, n_8, n_454);
	not g500(n_468, n_410);
	nand g501(n_469, n_460, n_461, n_443);
	nor g502(n_470, n_468, n_469);
	not g503(n_471, n_470);
	nor g504(n_472, n_456, n_461);
	not g505(n_473, n_472);
	nor g506(n_474, n_456, b[2]);
	not g507(n_475, n_474);
	nand g508(n_476, n_52, n_473, n_475);
	nor g509(n_477, n_468, n_476);
	not g510(n_478, n_477);
	nand g511(n_59, n_466, n_471, n_478);
	not g512(n_479, n_59);
	nor g513(n_480, n_59, n_451);
	not g514(n_481, n_480);
	nor g515(n_482, n_479, a[4]);
	not g516(n_483, n_482);
	nand g517(n_484, n_483, n_450);
	nand g518(n_64, n_481, n_484);
	nand g519(n_485, n_13, n_459, n_64);
	nand g520(n_67, n_448, b[7]);
	not g521(n_486, n_67);
	nor g522(n_487, n_453, b[6]);
	not g523(n_488, n_487);
	nand g524(n_489, n_67, n_488, n_446);
	nor g525(n_415, n_486, a[6]);
	not g526(n_490, n_415);
	nand g527(n_425, n_13, n_490);
	not g528(n_491, n_425);
	nor g529(n_492, n_13, n_491);
	not g530(n_493, n_492);
	nor g531(n_494, n_491, n_452);
	not g532(n_495, n_494);
	nand g533(n_496, n_489, n_493, n_495);
	nor g534(n_497, a[5], n_445);
	not g535(n_498, n_497);
	nand g536(n_156, n_467, n_498);
	nor g537(n_499, n_156, n_453, n_455);
	not g538(n_500, n_499);
	nor g539(n_501, n_156, n_455, b[6]);
	not g540(n_502, n_501);
	nand g541(n_503, n_500, n_502);
	not g542(n_504, n_503);
	nor g543(n_505, a[4], n_450);
	not g544(n_506, n_505);
	nand g545(n_171, n_8, n_506);
	nor g546(n_507, n_457, n_171, n_443);
	not g547(n_508, n_507);
	nor g548(n_509, n_457, n_171, b[1]);
	not g549(n_510, n_509);
	nand g550(n_511, n_508, n_510);
	not g551(n_512, n_511);
	nor g552(n_513, n_504, n_512);
	not g553(n_514, n_513);
	nor g554(n_515, n_486, n_452, n_445);
	not g555(n_516, n_515);
	nor g556(n_517, n_490, n_445);
	not g557(n_518, n_517);
	nand g558(n_432, n_516, n_518);
	not g559(n_519, n_432);
	nor g560(n_520, n_519, a[5]);
	not g561(n_521, n_520);
	nor g562(n_522, n_519, n_64);
	not g563(n_523, n_522);
	nand g564(n_524, n_149, n_521, n_523);
	nand g565(sub_wire0, n_514, n_524);
	and _ECO_0(w_eco0, !a[2], b[2], !b[7], b[4], !a[4], !b[1], a[0], !b[0]);
	and _ECO_1(w_eco1, !b[7], !a[7], b[4], !a[4], !b[1], a[0], !b[0]);
	and _ECO_2(w_eco2, !a[2], b[2], !b[7], a[7], !b[1], a[0]);
	and _ECO_3(w_eco3, !a[2], a[1], b[2], !b[7], b[4], !a[4], a[0], !b[0]);
	and _ECO_4(w_eco4, a[1], !b[7], !a[7], b[4], !a[4], a[0], !b[0]);
	and _ECO_5(w_eco5, !a[1], b[5], b[7], !a[7], b[4], !a[4], b[1], !b[0]);
	and _ECO_6(w_eco6, !a[1], !b[2], !b[5], !b[7], !a[7], b[4], !a[4], b[1]);
	and _ECO_7(w_eco7, !b[5], !b[7], a[7], b[4], !a[4], !b[1], !a[0]);
	and _ECO_8(w_eco8, !a[2], !a[1], b[2], b[5], b[7], !a[7], b[4], b[1]);
	and _ECO_9(w_eco9, !a[2], !a[1], b[2], !b[5], !b[7], !a[7], b[4], b[1], b[0]);
	and _ECO_10(w_eco10, !a[1], b[2], b[5], b[7], !a[7], !a[4], b[1], b[0]);
	and _ECO_11(w_eco11, a[2], !a[1], !b[5], !b[7], !a[7], b[4], !a[4], b[1]);
	and _ECO_12(w_eco12, a[2], !b[5], !b[7], !a[7], b[4], !a[4], a[0]);
	and _ECO_13(w_eco13, !a[2], a[1], b[2], !b[7], a[7], a[0]);
	and _ECO_14(w_eco14, !a[2], !a[1], b[5], b[7], !a[7], b[4], !a[4], b[1]);
	and _ECO_15(w_eco15, !b[2], !b[5], !b[7], !a[7], b[4], !a[4], a[0]);
	and _ECO_16(w_eco16, !a[2], b[2], !b[5], !b[7], b[4], !a[4], !b[1], !b[0]);
	and _ECO_17(w_eco17, a[1], !b[5], !b[7], a[7], !a[4], !a[0], !b[0]);
	and _ECO_18(w_eco18, !a[1], b[5], b[7], b[4], !a[4], !a[6], b[1], !b[0]);
	and _ECO_19(w_eco19, !b[5], !b[7], b[4], !a[4], b[6]);
	and _ECO_20(w_eco20, !a[1], !b[2], !b[5], !a[5], b[7], !a[7], b[1], !b[0]);
	and _ECO_21(w_eco21, b[5], !a[5], !b[7], a[7], !b[1], a[0]);
	and _ECO_22(w_eco22, !b[7], a[7], b[4], !a[4], a[6], !b[1], !a[0]);
	and _ECO_23(w_eco23, b[5], b[7], !a[7], b[4], !a[4], b[6], !a[0], !b[0]);
	and _ECO_24(w_eco24, !a[1], b[5], !a[5], !b[7], !a[7], !b[4], a[4], !b[0]);
	and _ECO_25(w_eco25, !a[2], !a[1], b[2], !b[5], !b[7], !a[7], !a[4], b[1], b[0]);
	and _ECO_26(w_eco26, !a[2], !a[1], b[2], b[5], b[7], !a[7], !a[4], b[1]);
	and _ECO_27(w_eco27, !a[2], !a[1], b[2], b[5], b[7], b[4], !a[6], b[1]);
	and _ECO_28(w_eco28, b[2], !b[5], !b[7], a[7], b[4], b[6], b[1]);
	and _ECO_29(w_eco29, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], b[1], b[0]);
	and _ECO_30(w_eco30, !a[2], !a[1], b[2], b[5], !a[7], b[4], a[6], b[1], b[0]);
	and _ECO_31(w_eco31, b[2], !b[5], a[5], !b[7], !a[7], b[4], b[1]);
	and _ECO_32(w_eco32, a[2], !a[1], !b[2], b[5], !a[5], !b[7], !a[7], a[4], b[1], !b[0]);
	and _ECO_33(w_eco33, a[2], !a[1], !b[2], !b[5], !b[7], !a[7], b[4], a[6], b[1]);
	and _ECO_34(w_eco34, !a[1], b[2], b[5], b[7], b[4], !a[4], !a[6], b[1]);
	and _ECO_35(w_eco35, a[2], !a[1], b[2], !b[5], !a[5], b[7], !a[7], b[1]);
	and _ECO_36(w_eco36, !a[1], !b[7], !a[7], b[4], !a[4], a[6], b[1], b[0]);
	and _ECO_37(w_eco37, a[2], a[5], !b[7], !a[7], b[4], !a[4], !b[1], a[0]);
	and _ECO_38(w_eco38, b[2], b[5], b[7], !a[7], b[4], !a[4], b[6], !a[0]);
	and _ECO_39(w_eco39, !b[7], b[4], !a[4], !a[6], !b[1], a[0]);
	and _ECO_40(w_eco40, !a[1], b[5], b[7], !a[7], b[4], !a[4], b[1], b[3]);
	and _ECO_41(w_eco41, a[2], !b[2], b[5], a[5], b[7], a[7], b[4], !a[4], !b[1], a[0], b[0]);
	and _ECO_42(w_eco42, a[2], !b[2], !a[5], b[4], !a[4], !a[6], !b[1], a[0], b[0]);
	and _ECO_43(w_eco43, a[2], !b[2], !b[5], !a[5], a[7], b[4], !a[4], !b[1], !a[0], b[0]);
	and _ECO_44(w_eco44, !a[2], !a[1], b[5], b[7], b[4], !a[4], !a[6], b[1]);
	and _ECO_45(w_eco45, !a[2], b[5], b[7], !a[7], b[4], !a[4], b[6], !a[0]);
	and _ECO_46(w_eco46, !a[2], b[2], !b[7], b[4], !a[4], a[6], !b[1], !b[0]);
	and _ECO_47(w_eco47, a[1], b[5], !a[5], !b[7], a[7], a[0]);
	and _ECO_48(w_eco48, a[1], !b[7], a[7], !a[4], a[6], !a[0], !b[0]);
	and _ECO_49(w_eco49, !a[1], b[5], b[7], b[4], !a[4], !b[6], a[6], b[1]);
	and _ECO_50(w_eco50, !b[7], b[4], !a[4], b[6], a[6]);
	and _ECO_51(w_eco51, a[1], !b[7], a[7], !b[6], !a[0]);
	and _ECO_52(w_eco52, !a[1], !b[5], !a[5], b[7], a[7], !b[4], a[4], !a[6], b[1], !b[0]);
	and _ECO_53(w_eco53, b[5], !a[5], !b[7], a[7], !b[4], a[4], !a[6]);
	and _ECO_54(w_eco54, !b[5], a[5], !b[7], !a[7], a[6]);
	and _ECO_55(w_eco55, !a[2], !a[1], b[2], b[5], b[7], !a[4], !a[6], b[1]);
	and _ECO_56(w_eco56, b[2], !b[5], !b[7], a[7], !a[4], b[6], b[1]);
	and _ECO_57(w_eco57, !a[2], !a[1], b[2], b[5], !a[7], !a[4], a[6], b[1], b[0]);
	and _ECO_58(w_eco58, !a[2], b[2], b[5], b[7], !a[7], !b[4], !a[4], b[1], !b[3]);
	and _ECO_59(w_eco59, a[1], b[5], b[7], !a[7], !b[4], !a[4], !b[1], !b[3], !b[0]);
	and _ECO_60(w_eco60, a[2], !a[1], !b[2], b[5], !a[5], !b[7], !a[7], !b[4], b[1], !b[0]);
	and _ECO_61(w_eco61, !a[1], b[2], b[5], b[7], !a[7], !a[3], b[4], b[1], b[3]);
	and _ECO_62(w_eco62, !a[1], b[2], b[5], b[7], !a[7], a[3], b[4], b[1], !b[3]);
	and _ECO_63(w_eco63, a[2], b[2], b[5], b[7], !a[7], b[4], a[4], a[0], !b[3]);
	and _ECO_64(w_eco64, a[2], a[1], b[2], b[5], b[7], !a[7], b[4], a[4], !b[1], !b[3]);
	and _ECO_65(w_eco65, b[2], b[5], b[7], !a[7], b[4], a[4], b[1], a[0], !b[3]);
	and _ECO_66(w_eco66, !a[2], b[2], b[5], b[7], !a[7], b[4], a[4], b[1], !b[3]);
	and _ECO_67(w_eco67, !a[1], b[2], b[5], b[7], b[4], !b[6], a[6], b[1]);
	and _ECO_68(w_eco68, b[2], !b[7], a[7], b[4], b[6], a[6], b[1]);
	and _ECO_69(w_eco69, !a[2], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1]);
	and _ECO_70(w_eco70, !a[2], b[2], b[5], b[7], b[4], a[4], !a[6], b[1], !b[3]);
	and _ECO_71(w_eco71, !a[2], !b[5], !a[5], b[7], !a[7], a[4], !b[3], b[0]);
	and _ECO_72(w_eco72, !a[2], b[2], b[5], !a[7], b[4], a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_73(w_eco73, !a[2], b[2], !b[5], !a[5], !a[7], b[4], a[4], b[1], !b[3], b[0]);
	and _ECO_74(w_eco74, a[2], !a[1], !b[5], !a[5], b[7], !a[7], b[4], b[1], b[3]);
	and _ECO_75(w_eco75, !a[2], !a[1], b[5], b[7], !a[7], !a[3], b[4], b[1], b[3]);
	and _ECO_76(w_eco76, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], b[4], !a[6], b[1]);
	and _ECO_77(w_eco77, !a[2], !a[1], b[2], !b[7], !a[7], b[6], a[6], !b[0]);
	and _ECO_78(w_eco78, !a[2], b[2], !b[5], !b[7], !a[7], !a[4], !a[6], b[1]);
	and _ECO_79(w_eco79, !a[2], b[2], !b[5], !b[7], !a[7], b[4], !a[6], b[1]);
	and _ECO_80(w_eco80, a[1], b[5], b[7], !a[7], b[4], a[4], a[0], !b[3], !b[0]);
	and _ECO_81(w_eco81, a[1], b[5], b[7], !a[7], b[4], a[4], !b[1], !b[3], !b[0]);
	and _ECO_82(w_eco82, a[2], a[1], !b[2], b[5], b[7], !a[7], b[4], a[4], !b[3], !b[0]);
	and _ECO_83(w_eco83, a[2], !a[1], !b[2], !b[5], b[7], a[4], b[6], !a[6], b[1], !b[0]);
	and _ECO_84(w_eco84, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[4], !a[6], b[1]);
	and _ECO_85(w_eco85, a[2], !a[1], !b[2], !b[5], !b[7], !a[7], b[4], !b[6], !a[6]);
	and _ECO_86(w_eco86, a[1], !b[7], b[4], !a[4], !b[6], !a[6]);
	and _ECO_87(w_eco87, !b[7], b[4], !a[4], !b[6], !a[6], !b[1]);
	and _ECO_88(w_eco88, !b[2], b[5], a[5], !a[7], b[4], !a[4], a[6], a[0], !b[0]);
	and _ECO_89(w_eco89, !b[2], !b[5], !a[5], b[7], !a[7], a[6], a[0], !b[0]);
	and _ECO_90(w_eco90, b[5], b[7], b[4], !a[4], b[6], !a[6], !a[0], !b[0]);
	and _ECO_91(w_eco91, !b[2], !b[5], !a[5], b[7], !a[7], b[6], !a[0], !b[0]);
	and _ECO_92(w_eco92, a[2], b[2], b[5], a[5], !a[7], b[4], !a[4], a[6], a[0]);
	and _ECO_93(w_eco93, a[2], b[2], !b[5], !a[5], b[7], !a[7], a[6], a[0]);
	and _ECO_94(w_eco94, b[2], b[5], b[7], b[4], !a[4], b[6], !a[6], !a[0]);
	and _ECO_95(w_eco95, a[2], b[2], !b[5], !a[5], b[7], !a[7], b[6], !a[0]);
	and _ECO_96(w_eco96, !a[2], !b[5], !a[5], b[7], !a[7], b[6], !a[0], b[0]);
	and _ECO_97(w_eco97, !a[2], b[2], !b[5], !a[5], a[7], b[4], !a[4], !b[6], a[6], !b[1]);
	and _ECO_98(w_eco98, a[2], a[1], !b[2], b[5], a[5], b[7], a[7], b[4], !a[4], a[0], b[0]);
	and _ECO_99(w_eco99, a[2], a[1], !b[2], !a[5], b[4], !a[4], !a[6], a[0], b[0]);
	and _ECO_100(w_eco100, a[2], a[1], !b[2], !b[5], !a[5], a[7], b[4], !a[4], !a[0], b[0]);
	and _ECO_101(w_eco101, !a[1], b[5], b[7], b[4], !a[4], !a[6], b[1], b[3]);
	and _ECO_102(w_eco102, a[2], !b[2], !a[5], b[7], a[7], b[6], a[6], !b[1], b[0]);
	and _ECO_103(w_eco103, a[2], !b[2], b[5], b[4], !a[4], !a[6], !b[1], a[0], b[0]);
	and _ECO_104(w_eco104, a[2], !b[2], b[5], b[4], !a[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_105(w_eco105, !a[2], !b[2], b[5], a[5], !a[7], b[4], !a[4], a[6], a[0]);
	and _ECO_106(w_eco106, !a[2], !b[2], !b[5], !a[5], b[7], !a[7], a[6], a[0]);
	and _ECO_107(w_eco107, !a[2], b[5], b[7], b[4], !a[4], b[6], !a[6], !a[0]);
	and _ECO_108(w_eco108, !a[2], b[2], !b[5], !a[5], !a[7], b[4], !a[4], a[6], !b[1], !a[0], !b[0]);
	and _ECO_109(w_eco109, !b[2], b[5], a[5], b[7], b[4], !a[4], !b[6], a[6], a[0]);
	and _ECO_110(w_eco110, !b[5], !a[5], a[7], b[4], !a[4], !b[6], a[6], !b[1], !a[0]);
	and _ECO_111(w_eco111, b[5], !a[5], !b[7], b[4], !a[4], !b[6], !b[1], !b[0]);
	and _ECO_112(w_eco112, !a[1], b[2], !b[5], !a[5], b[7], a[7], !b[4], a[4], !a[6], b[1]);
	and _ECO_113(w_eco113, !a[1], a[5], b[7], !b[4], a[4], b[6], !a[6], b[1]);
	and _ECO_114(w_eco114, !a[1], b[5], !b[7], !a[7], !b[4], a[4], b[6], !a[6], b[1], b[0]);
	and _ECO_115(w_eco115, a[2], !b[2], b[5], !a[5], a[7], !b[4], a[4], !a[6], b[0]);
	and _ECO_116(w_eco116, a[2], !a[1], !b[5], !a[5], b[7], !a[7], !b[4], a[4], a[6], b[1]);
	and _ECO_117(w_eco117, !a[2], !a[1], !b[5], !a[5], b[7], a[7], !b[4], a[4], !a[6], b[1]);
	and _ECO_118(w_eco118, b[5], !a[5], !b[7], !a[7], !b[4], a[4], b[1], !b[0]);
	and _ECO_119(w_eco119, !a[2], !a[1], b[2], a[5], !b[7], !a[7], !b[4], a[4], !b[6], !b[0]);
	and _ECO_120(w_eco120, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[4], !b[1], !b[3]);
	and _ECO_121(w_eco121, a[2], b[2], b[5], b[7], !a[7], !b[4], !a[4], a[0], !b[3]);
	and _ECO_122(w_eco122, a[2], a[1], b[2], b[5], b[7], !a[7], !b[4], !a[4], !b[1], !b[3]);
	and _ECO_123(w_eco123, !a[1], b[2], b[5], b[7], !a[4], !b[6], a[6], b[1]);
	and _ECO_124(w_eco124, b[2], !b[7], a[7], !a[4], b[6], a[6], b[1]);
	and _ECO_125(w_eco125, a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[4], b[1], b[3]);
	and _ECO_126(w_eco126, !a[2], !a[1], b[5], b[7], !a[7], !a[3], !a[4], b[1], b[3]);
	and _ECO_127(w_eco127, !a[2], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1]);
	and _ECO_128(w_eco128, !a[2], b[2], b[5], b[7], !b[4], !a[4], !a[6], b[1], !b[3]);
	and _ECO_129(w_eco129, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[4], !a[6], b[1]);
	and _ECO_130(w_eco130, a[1], b[5], b[7], !a[7], a[3], !b[4], !a[4], !b[1], !b[0]);
	and _ECO_131(w_eco131, !a[2], a[1], !b[5], !a[5], b[7], !a[7], !b[4], !b[1], !b[3]);
	and _ECO_132(w_eco132, a[1], b[5], b[7], !a[7], !b[4], !a[4], a[0], !b[3], !b[0]);
	and _ECO_133(w_eco133, a[2], a[1], !b[2], b[5], b[7], !a[7], !b[4], !a[4], !b[3], !b[0]);
	and _ECO_134(w_eco134, a[2], !a[1], !b[2], !b[5], b[7], !b[4], b[6], !a[6], b[1], !b[0]);
	and _ECO_135(w_eco135, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[7], !b[4], !a[6], b[1]);
	and _ECO_136(w_eco136, a[2], !a[1], !b[2], !b[5], !b[7], !a[7], !a[4], a[6], b[1]);
	and _ECO_137(w_eco137, a[2], !a[1], !b[2], !b[5], !b[7], !a[7], !a[4], !b[6], !a[6]);
	and _ECO_138(w_eco138, b[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], a[0]);
	and _ECO_139(w_eco139, b[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], b[0]);
	and _ECO_140(w_eco140, b[2], b[5], b[7], !a[7], b[4], a[4], b[1], !b[3], b[0]);
	and _ECO_141(w_eco141, !a[1], b[2], b[5], b[7], !a[3], b[4], !a[6], b[1], b[3]);
	and _ECO_142(w_eco142, !a[1], b[2], b[5], !a[7], !a[3], b[4], a[6], b[1], b[3], b[0]);
	and _ECO_143(w_eco143, a[2], !a[1], b[2], !b[5], !a[5], !a[7], !a[3], b[4], b[1], b[3]);
	and _ECO_144(w_eco144, !a[1], b[2], b[5], b[7], a[3], b[4], !a[6], b[1], !b[3]);
	and _ECO_145(w_eco145, !a[1], b[2], b[5], !a[7], a[3], b[4], a[6], b[1], !b[3], b[0]);
	and _ECO_146(w_eco146, a[2], !a[1], b[2], !b[5], !a[5], !a[7], a[3], b[4], b[1], !b[3]);
	and _ECO_147(w_eco147, a[2], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], a[0]);
	and _ECO_148(w_eco148, a[2], a[1], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], !b[1]);
	and _ECO_149(w_eco149, a[1], !b[7], a[7], !a[6], a[0]);
	and _ECO_150(w_eco150, a[2], b[2], !b[5], !b[7], a[7], b[4], b[6], !b[3]);
	and _ECO_151(w_eco151, !a[1], b[2], !b[5], !b[7], a[7], b[4], !b[1], !a[0], b[3]);
	and _ECO_152(w_eco152, !a[1], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[3], b[0]);
	and _ECO_153(w_eco153, a[2], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], !b[3]);
	and _ECO_154(w_eco154, !a[1], b[2], b[5], b[7], !a[7], !a[3], b[4], a[4], !b[3], b[0]);
	and _ECO_155(w_eco155, b[2], b[5], b[7], b[4], a[4], !b[6], a[6], b[1], !b[3]);
	and _ECO_156(w_eco156, !a[2], !a[1], !b[5], !b[7], a[7], !a[3], b[4], !b[1], !a[0]);
	and _ECO_157(w_eco157, a[2], !a[1], !b[2], !b[5], b[7], b[4], a[4], b[6], !a[6], b[1], b[3]);
	and _ECO_158(w_eco158, a[2], !a[1], !b[2], b[5], !a[5], !b[7], b[4], a[4], !a[6], b[1]);
	and _ECO_159(w_eco159, a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[3], b[4], b[1]);
	and _ECO_160(w_eco160, !b[7], a[7], !a[6], !b[1], a[0]);
	and _ECO_161(w_eco161, !b[7], a[7], !b[6], !b[1], !a[0]);
	and _ECO_162(w_eco162, !a[2], !b[5], !a[5], b[7], a[7], !b[4], a[4], !a[6], !b[3]);
	and _ECO_163(w_eco163, a[5], b[7], !b[4], a[4], b[6], !a[6], !b[3]);
	and _ECO_164(w_eco164, b[5], !b[7], !a[7], !b[4], a[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_165(w_eco165, a[2], !b[5], !a[5], b[7], !a[7], !b[4], a[4], a[6], !b[3]);
	and _ECO_166(w_eco166, !a[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], a[0], b[3]);
	and _ECO_167(w_eco167, !a[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], b[3], b[0]);
	and _ECO_168(w_eco168, !a[2], b[5], b[7], !a[7], !a[3], b[4], a[4], b[1], a[0], !b[3]);
	and _ECO_169(w_eco169, !a[2], b[5], b[7], !a[7], !a[3], b[4], a[4], b[1], !b[3], b[0]);
	and _ECO_170(w_eco170, !a[2], !a[1], b[5], b[7], !a[3], b[4], !a[6], b[1], b[3]);
	and _ECO_171(w_eco171, !a[2], !a[1], !b[5], !b[7], a[7], !a[3], b[4], b[6]);
	and _ECO_172(w_eco172, !a[2], !a[1], b[5], !a[7], !a[3], b[4], a[6], b[1], b[3], b[0]);
	and _ECO_173(w_eco173, !a[2], !a[1], !b[2], !b[5], !a[5], !a[7], !a[3], b[4], b[1], b[3]);
	and _ECO_174(w_eco174, !a[2], !a[1], b[5], b[7], !a[7], a[3], b[4], a[4], a[0], b[3]);
	and _ECO_175(w_eco175, !a[2], !a[1], b[5], b[7], !a[7], a[3], b[4], a[4], b[3], b[0]);
	and _ECO_176(w_eco176, !a[2], !a[1], b[5], b[7], !a[7], !a[3], b[4], a[4], a[0], !b[3]);
	and _ECO_177(w_eco177, !a[2], !a[1], b[5], b[7], !a[7], !a[3], b[4], a[4], !b[3], b[0]);
	and _ECO_178(w_eco178, a[1], !b[7], !a[7], !a[3], b[4], b[1], a[0], b[3], !b[0]);
	and _ECO_179(w_eco179, !a[1], !b[7], !a[7], !a[3], b[4], !b[1], a[0], b[3], !b[0]);
	and _ECO_180(w_eco180, !a[2], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], b[1]);
	and _ECO_181(w_eco181, !a[2], a[1], !b[5], !a[5], b[7], !a[7], b[4], a[4], !a[6], !b[3]);
	and _ECO_182(w_eco182, !a[2], b[2], !b[7], !a[7], b[6], a[6], b[1], !b[0]);
	and _ECO_183(w_eco183, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], b[4], b[6], b[1]);
	and _ECO_184(w_eco184, a[1], b[5], b[7], !a[7], a[3], b[4], a[4], a[0], !b[0]);
	and _ECO_185(w_eco185, a[1], b[5], b[7], !a[7], a[3], b[4], a[4], !b[1], !b[0]);
	and _ECO_186(w_eco186, !a[2], a[1], b[2], !b[7], !a[3], a[0], b[3], !b[0]);
	and _ECO_187(w_eco187, a[1], !b[5], !b[7], a[7], b[4], b[6], !b[0]);
	and _ECO_188(w_eco188, b[2], b[5], b[7], !a[7], a[3], b[4], a[4], a[0], !b[0]);
	and _ECO_189(w_eco189, b[2], b[5], b[7], !a[7], a[3], b[4], a[4], !b[3], !b[0]);
	and _ECO_190(w_eco190, a[2], a[1], !b[2], b[5], b[7], !a[7], a[3], b[4], a[4], !b[0]);
	and _ECO_191(w_eco191, a[1], b[5], b[7], b[4], a[4], !a[6], b[1], a[0], !b[3], !b[0]);
	and _ECO_192(w_eco192, a[2], a[1], !b[5], !b[7], !a[7], b[4], b[1], a[0], !b[0]);
	and _ECO_193(w_eco193, a[2], a[1], !b[2], b[5], b[7], b[4], a[4], !a[6], b[1], !b[3], !b[0]);
	and _ECO_194(w_eco194, a[2], a[1], !b[2], !b[5], !a[5], !a[7], b[4], a[4], b[1], !b[3], !b[0]);
	and _ECO_195(w_eco195, !a[1], b[5], a[5], b[7], b[6], !a[6], b[1], !b[0]);
	and _ECO_196(w_eco196, a[2], !b[2], b[5], !a[5], !b[7], a[7], a[4], !b[6]);
	and _ECO_197(w_eco197, a[2], !a[1], !b[2], !b[7], !a[7], b[4], b[6], a[6]);
	and _ECO_198(w_eco198, a[2], !a[1], !b[2], !b[7], !a[7], b[4], a[4], !b[6], !a[6]);
	and _ECO_199(w_eco199, !a[1], b[5], a[5], b[7], b[6], !a[6], b[1], b[3]);
	and _ECO_200(w_eco200, a[1], b[5], b[7], !a[7], a[3], b[4], a[4], !b[3], !b[0]);
	and _ECO_201(w_eco201, !a[1], !b[2], b[5], !a[5], !b[7], !a[7], a[3], a[4], !b[3], !b[0]);
	and _ECO_202(w_eco202, a[1], !b[7], b[4], !a[4], b[6], a[0]);
	and _ECO_203(w_eco203, a[2], b[5], a[5], b[7], b[4], !a[4], !b[6], a[6], a[0]);
	and _ECO_204(w_eco204, !a[2], a[1], b[2], !b[5], !a[5], a[7], b[4], !a[4], !b[6], a[6]);
	and _ECO_205(w_eco205, a[2], a[1], !b[2], !a[5], b[7], a[7], b[6], a[6], b[0]);
	and _ECO_206(w_eco206, a[2], a[1], !b[2], b[5], b[4], !a[4], !a[6], a[0], b[0]);
	and _ECO_207(w_eco207, a[2], a[1], !b[2], b[5], !a[4], !b[6], !a[6], b[1], b[0]);
	and _ECO_208(w_eco208, !a[1], b[5], b[7], !a[3], b[4], !a[4], !a[6], b[1]);
	and _ECO_209(w_eco209, a[2], !b[2], b[5], !a[5], b[4], !a[4], b[6], !b[1], a[0], b[0]);
	and _ECO_210(w_eco210, a[2], !b[5], !a[5], !a[7], !b[6], a[6], a[0]);
	and _ECO_211(w_eco211, a[2], !b[2], b[5], a[7], b[4], !a[4], b[6], a[6], !b[1], b[0]);
	and _ECO_212(w_eco212, a[2], !b[2], !a[5], b[4], !a[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_213(w_eco213, !a[2], a[1], b[2], !b[5], !a[5], !a[7], b[4], !a[4], a[6], !a[0], !b[0]);
	and _ECO_214(w_eco214, !a[2], a[1], b[2], !b[7], b[4], !a[4], !b[6], !b[0]);
	and _ECO_215(w_eco215, !b[5], !a[5], !a[7], b[4], !a[4], !b[6], a[6], !b[1], a[0], !b[0]);
	and _ECO_216(w_eco216, !a[2], !b[5], !a[5], b[7], !a[7], b[6], !a[6], !a[0]);
	and _ECO_217(w_eco217, a[1], !b[5], !a[5], a[7], b[4], !a[4], !b[6], a[6], !a[0]);
	and _ECO_218(w_eco218, a[1], b[5], !a[5], !b[7], b[4], !a[4], !b[6], !b[0]);
	and _ECO_219(w_eco219, !a[1], !b[2], b[5], a[5], !a[7], b[4], !a[4], !b[6], a[6], b[1]);
	and _ECO_220(w_eco220, b[2], !b[5], !a[5], b[7], a[7], !a[3], !b[4], a[4], !b[1], !a[0], b[3]);
	and _ECO_221(w_eco221, b[2], !b[5], !a[5], b[7], a[7], !b[4], a[4], !a[6], !b[3]);
	and _ECO_222(w_eco222, a[2], b[2], !b[5], !a[5], b[7], !a[7], a[4], !b[3]);
	and _ECO_223(w_eco223, !a[5], b[7], a[7], !b[4], a[4], b[6], a[6]);
	and _ECO_224(w_eco224, !a[2], !a[1], b[2], b[5], !a[5], b[7], a[7], !b[6], !a[6], b[1]);
	and _ECO_225(w_eco225, b[5], !a[5], !b[7], a[7], !b[4], a[4], !b[6]);
	and _ECO_226(w_eco226, !b[5], a[5], !b[7], !a[7], !b[6]);
	and _ECO_227(w_eco227, !a[1], !b[5], !a[5], !a[7], !b[6], a[6], b[1], b[0]);
	and _ECO_228(w_eco228, b[5], !a[5], a[7], !b[4], a[4], !b[6], !a[6]);
	and _ECO_229(w_eco229, !a[2], !b[5], !a[5], b[7], !a[7], a[3], a[4], b[0]);
	and _ECO_230(w_eco230, !a[2], b[2], b[5], !a[7], a[3], b[4], a[4], a[6], b[1], b[0]);
	and _ECO_231(w_eco231, !a[2], !b[5], !a[5], b[7], a[7], a[3], !b[4], a[4], !a[6]);
	and _ECO_232(w_eco232, a[5], b[7], a[3], !b[4], a[4], b[6], !a[6]);
	and _ECO_233(w_eco233, b[5], !b[7], !a[7], a[3], !b[4], a[4], b[6], !a[6], b[0]);
	and _ECO_234(w_eco234, a[2], b[2], !b[5], !a[5], b[7], a[3], !b[4], a[4], !a[6]);
	and _ECO_235(w_eco235, !b[5], !a[5], !a[7], a[4], !b[6], a[6], !b[3], b[0]);
	and _ECO_236(w_eco236, b[2], b[5], b[7], a[3], b[4], a[4], !a[6], b[1], !b[3]);
	and _ECO_237(w_eco237, b[2], b[5], !a[7], a[3], b[4], a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_238(w_eco238, !a[5], b[7], a[7], !b[4], a[4], !b[6], !a[6]);
	and _ECO_239(w_eco239, a[2], !b[2], b[5], !a[5], !b[4], a[4], b[6], !a[6], b[0]);
	and _ECO_240(w_eco240, a[2], !a[1], !b[5], !a[5], b[7], !b[4], a[4], !b[6], !a[6], b[1]);
	and _ECO_241(w_eco241, a[2], !b[5], !a[5], b[7], !b[4], a[4], !b[6], !a[6], !b[3]);
	and _ECO_242(w_eco242, a[1], b[5], !b[7], !a[7], !b[4], a[4], b[6], !a[6], !b[1], !b[3]);
	and _ECO_243(w_eco243, !a[1], b[5], !a[5], b[7], !b[4], a[4], b[6], a[6], !b[0]);
	and _ECO_244(w_eco244, !a[1], b[5], !a[5], !b[4], a[4], !b[6], !a[6], !b[0]);
	and _ECO_245(w_eco245, !a[1], !b[2], !b[5], !a[5], !a[7], !b[6], a[6], b[1]);
	and _ECO_246(w_eco246, b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], a[0]);
	and _ECO_247(w_eco247, b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], b[0]);
	and _ECO_248(w_eco248, b[2], b[5], b[7], !a[7], !b[4], !a[4], b[1], !b[3], b[0]);
	and _ECO_249(w_eco249, !a[1], b[2], b[5], !a[7], !a[3], !a[4], a[6], b[1], b[3], b[0]);
	and _ECO_250(w_eco250, !a[1], b[2], b[5], b[7], a[3], !a[4], !a[6], b[1], !b[3]);
	and _ECO_251(w_eco251, !a[1], b[2], b[5], !a[7], a[3], !a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_252(w_eco252, a[2], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], a[0]);
	and _ECO_253(w_eco253, a[2], a[1], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], !b[1]);
	and _ECO_254(w_eco254, a[2], b[2], !b[5], !b[7], a[7], !a[4], b[6], !b[3]);
	and _ECO_255(w_eco255, !a[1], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[3], b[0]);
	and _ECO_256(w_eco256, a[2], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], !b[3]);
	and _ECO_257(w_eco257, !a[1], b[2], b[5], b[7], !a[7], !a[3], !b[4], !a[4], !b[3], b[0]);
	and _ECO_258(w_eco258, !a[2], !b[5], !a[5], b[7], !a[7], !b[4], !b[3], b[0]);
	and _ECO_259(w_eco259, !a[2], b[2], b[5], !a[7], !b[4], !a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_260(w_eco260, b[2], b[5], b[7], !b[4], !a[4], !b[6], a[6], b[1], !b[3]);
	and _ECO_261(w_eco261, !a[2], b[2], !a[5], !a[7], !b[4], !a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_262(w_eco262, a[2], !a[1], !b[2], !b[5], b[7], !b[4], !a[4], b[6], !a[6], b[1], b[3]);
	and _ECO_263(w_eco263, a[2], !a[1], !b[2], b[5], !a[5], !b[7], !b[4], !a[4], !a[6], b[1]);
	and _ECO_264(w_eco264, !a[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], a[0], b[3]);
	and _ECO_265(w_eco265, !a[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], b[3], b[0]);
	and _ECO_266(w_eco266, !a[2], b[5], b[7], !a[7], !a[3], !b[4], !a[4], b[1], a[0], !b[3]);
	and _ECO_267(w_eco267, !a[2], b[5], b[7], !a[7], !a[3], !b[4], !a[4], b[1], !b[3], b[0]);
	and _ECO_268(w_eco268, !a[2], !a[1], !b[5], !b[7], a[7], !a[3], !a[4], b[6]);
	and _ECO_269(w_eco269, !a[2], !a[1], b[5], !a[7], !a[3], !a[4], a[6], b[1], b[3], b[0]);
	and _ECO_270(w_eco270, !a[2], !a[1], b[5], b[7], !a[7], a[3], !b[4], !a[4], a[0], b[3]);
	and _ECO_271(w_eco271, !a[2], !a[1], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[3], b[0]);
	and _ECO_272(w_eco272, !a[2], !a[1], b[5], b[7], !a[7], !a[3], !b[4], !a[4], a[0], !b[3]);
	and _ECO_273(w_eco273, !a[2], !a[1], b[5], b[7], !a[7], !a[3], !b[4], !a[4], !b[3], b[0]);
	and _ECO_274(w_eco274, a[1], !b[7], !a[7], !a[3], !a[4], b[1], a[0], b[3], !b[0]);
	and _ECO_275(w_eco275, !a[1], !b[7], !a[7], !a[3], !a[4], !b[1], a[0], b[3], !b[0]);
	and _ECO_276(w_eco276, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[4], b[6], b[1]);
	and _ECO_277(w_eco277, a[1], b[5], a[5], b[7], !b[4], !a[4], !a[6], !b[3], !b[0]);
	and _ECO_278(w_eco278, a[1], b[5], !a[5], b[7], !b[4], !a[4], a[6], !b[1], !b[3], !b[0]);
	and _ECO_279(w_eco279, a[1], b[5], a[5], !a[7], !b[4], !a[4], !a[6], !b[1], !b[3], !b[0]);
	and _ECO_280(w_eco280, a[1], b[5], !a[5], !b[7], !a[4], !b[6], !b[1], !b[0]);
	and _ECO_281(w_eco281, b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], a[0], !b[0]);
	and _ECO_282(w_eco282, b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], !b[3], !b[0]);
	and _ECO_283(w_eco283, a[1], b[5], b[7], !a[7], a[3], !b[4], !a[4], a[0], !b[0]);
	and _ECO_284(w_eco284, a[2], a[1], !b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], !b[0]);
	and _ECO_285(w_eco285, a[2], a[1], !b[2], !b[5], !a[5], !a[7], !b[4], !a[4], b[1], !b[3], !b[0]);
	and _ECO_286(w_eco286, a[2], !b[2], b[5], !a[5], !b[7], a[7], !b[4], !b[6]);
	and _ECO_287(w_eco287, a[2], !a[1], !b[2], !b[7], !a[7], !a[4], b[6], a[6]);
	and _ECO_288(w_eco288, a[2], !a[1], !b[2], !b[7], !a[7], !b[4], !a[4], !b[6], !a[6]);
	and _ECO_289(w_eco289, !a[1], !b[2], b[5], !a[5], !b[7], !a[7], a[3], !b[4], !b[3], !b[0]);
	and _ECO_290(w_eco290, b[2], b[5], b[7], a[3], b[4], a[4], !a[6], b[1], a[0]);
	and _ECO_291(w_eco291, b[2], b[5], !a[7], a[3], b[4], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_292(w_eco292, a[2], a[1], b[2], a[5], !b[7], !a[7], !a[3], b[4], b[1], a[0], b[3]);
	and _ECO_293(w_eco293, a[1], !b[7], !a[3], b[4], !a[6], b[1], a[0], b[3]);
	and _ECO_294(w_eco294, b[2], b[5], b[7], !a[7], !a[3], b[4], b[6], b[1], !a[0], b[3]);
	and _ECO_295(w_eco295, b[2], !b[5], !b[7], !a[7], a[3], b[4], !a[6], b[1], !b[3]);
	and _ECO_296(w_eco296, b[2], b[5], b[7], b[4], a[4], !a[6], b[1], a[0], !b[3]);
	and _ECO_297(w_eco297, b[2], b[5], !a[7], b[4], a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_298(w_eco298, a[2], b[2], !b[5], !b[7], a[7], a[3], b[4], b[6]);
	and _ECO_299(w_eco299, a[1], b[2], !b[5], !a[5], b[7], a[7], !a[3], a[4], !b[1], !a[0], b[3], b[0]);
	and _ECO_300(w_eco300, a[2], b[2], b[5], a[5], b[7], b[4], a[4], !a[6], !b[3]);
	and _ECO_301(w_eco301, a[2], a[1], b[2], b[5], !a[5], b[7], b[4], a[4], a[6], !b[1], !b[3]);
	and _ECO_302(w_eco302, a[2], a[1], b[2], a[5], !b[7], b[4], !a[6], !b[1], a[0], !b[3]);
	and _ECO_303(w_eco303, a[2], a[1], b[2], b[5], !a[5], !b[7], b[4], a[4], !b[6], !b[1], !b[3]);
	and _ECO_304(w_eco304, a[2], b[2], !b[7], a[7], b[4], b[6], a[6], !b[3]);
	and _ECO_305(w_eco305, a[2], !a[1], b[2], b[5], !a[7], a[3], b[4], a[4], a[6], !b[3], b[0]);
	and _ECO_306(w_eco306, a[2], a[1], b[2], b[5], a[5], !a[7], b[4], a[4], !a[6], !b[1], !b[3]);
	and _ECO_307(w_eco307, a[2], b[2], !b[5], !b[7], b[4], b[6], !a[6], !b[3]);
	and _ECO_308(w_eco308, a[2], b[2], b[5], b[7], b[4], a[4], !b[6], a[6], !b[3]);
	and _ECO_309(w_eco309, a[2], a[1], b[5], !a[5], b[7], b[4], a[4], b[6], !a[6], !b[3]);
	and _ECO_310(w_eco310, a[1], !a[5], b[7], a[7], a[4], b[6], a[6], !b[1]);
	and _ECO_311(w_eco311, a[1], !b[5], !a[5], a[7], a[4], !b[6], !a[6], !b[1]);
	and _ECO_312(w_eco312, a[2], b[2], b[5], a[5], !a[7], b[4], a[4], !b[6], a[6], !b[3]);
	and _ECO_313(w_eco313, !a[1], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], a[0], b[3]);
	and _ECO_314(w_eco314, !a[1], b[2], b[5], !a[7], a[3], b[4], a[4], a[6], a[0], b[3], b[0]);
	and _ECO_315(w_eco315, a[2], !a[1], b[2], a[5], !b[7], !a[7], !a[3], b[4], !b[1], a[0], b[3]);
	and _ECO_316(w_eco316, !a[1], !b[7], !a[3], b[4], !a[6], !b[1], a[0], b[3]);
	and _ECO_317(w_eco317, !a[1], b[2], b[5], b[7], !a[7], !a[3], b[4], b[6], !a[0], b[0]);
	and _ECO_318(w_eco318, a[2], !a[1], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], !b[3]);
	and _ECO_319(w_eco319, !a[2], b[5], b[7], a[3], b[4], a[4], !b[6], a[6], b[1], b[3]);
	and _ECO_320(w_eco320, !a[2], b[2], !a[5], !a[7], a[3], b[4], a[4], a[6], b[1], b[0]);
	and _ECO_321(w_eco321, !a[2], a[1], !b[5], b[7], a[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_322(w_eco322, !a[2], a[1], b[5], !b[7], b[6], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_323(w_eco323, !a[2], a[1], b[5], !b[7], !a[7], a[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_324(w_eco324, !a[2], !a[1], !b[5], !a[5], !a[7], a[3], b[4], a[4], a[0], b[3], b[0]);
	and _ECO_325(w_eco325, !a[2], !a[1], b[5], b[7], !a[3], b[4], a[4], !a[6], a[0], !b[3]);
	and _ECO_326(w_eco326, !a[2], !a[1], b[5], !a[7], !a[3], b[4], a[4], a[6], a[0], !b[3], b[0]);
	and _ECO_327(w_eco327, a[2], a[1], !b[2], b[5], !a[3], b[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_328(w_eco328, a[2], a[1], b[5], !a[7], b[4], a[4], b[6], a[6], b[1], a[0], !b[3]);
	and _ECO_329(w_eco329, a[2], a[1], !b[2], b[5], b[4], !b[6], !a[6], b[1], b[0]);
	and _ECO_330(w_eco330, a[2], a[1], !b[2], b[5], !a[7], b[4], a[4], b[6], a[6], b[1], !a[0]);
	and _ECO_331(w_eco331, a[2], !b[2], b[5], !a[5], a[7], a[3], a[4], !a[6], !b[3], b[0]);
	and _ECO_332(w_eco332, a[2], !a[1], b[5], !a[5], b[7], a[3], b[4], a[4], !a[6], !b[3], b[0]);
	and _ECO_333(w_eco333, a[2], !a[1], !b[2], !b[5], b[7], !a[3], b[4], a[4], b[6], !a[6], b[1]);
	and _ECO_334(w_eco334, !a[1], b[5], a[5], b[7], !a[3], b[6], !a[6], b[1]);
	and _ECO_335(w_eco335, a[1], !b[2], a[5], b[7], a[3], a[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_336(w_eco336, a[1], !b[2], b[5], !b[7], !a[7], a[3], a[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_337(w_eco337, a[2], !a[1], !b[2], b[5], !a[3], b[4], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_338(w_eco338, !a[2], b[5], b[7], a[3], b[4], a[4], !a[6], b[1], a[0], b[3]);
	and _ECO_339(w_eco339, !a[2], b[5], !a[7], a[3], b[4], a[4], a[6], b[1], a[0], b[3], b[0]);
	and _ECO_340(w_eco340, !a[2], !b[2], !b[5], !b[7], !a[7], b[4], b[1], a[0], b[3]);
	and _ECO_341(w_eco341, !a[2], !b[5], !b[7], a[7], b[4], b[6], b[1], b[3]);
	and _ECO_342(w_eco342, !a[2], b[5], b[7], !a[7], !a[3], b[4], b[6], b[1], !a[0], b[3]);
	and _ECO_343(w_eco343, !a[2], b[5], b[7], !a[3], b[4], a[4], !a[6], b[1], a[0], !b[3]);
	and _ECO_344(w_eco344, !a[2], b[5], !a[7], !a[3], b[4], a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_345(w_eco345, !a[2], !b[5], !b[7], a[7], !a[3], b[4], b[6], b[1]);
	and _ECO_346(w_eco346, !a[2], !a[1], !b[2], !b[5], b[7], a[3], a[4], b[6], !a[6], !b[3]);
	and _ECO_347(w_eco347, !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], a[4], !a[6], !b[3]);
	and _ECO_348(w_eco348, !a[1], !b[2], b[5], !a[5], !b[7], a[3], b[4], a[4], !a[6], !b[3]);
	and _ECO_349(w_eco349, !a[2], !a[1], b[5], b[7], a[3], b[4], a[4], !a[6], a[0], b[3]);
	and _ECO_350(w_eco350, !a[2], !a[1], b[5], !a[7], a[3], b[4], a[4], a[6], a[0], b[3], b[0]);
	and _ECO_351(w_eco351, !a[2], !a[1], !b[5], !b[7], a[7], b[4], b[6], b[3]);
	and _ECO_352(w_eco352, !a[2], !a[1], b[5], b[7], !a[7], !a[3], b[4], b[6], !a[0], b[0]);
	and _ECO_353(w_eco353, b[2], b[5], a[5], b[7], !a[7], a[3], b[4], a[4], b[1]);
	and _ECO_354(w_eco354, a[2], !a[1], b[2], b[5], a[5], !a[7], !a[3], b[4], a[6], b[1], b[3]);
	and _ECO_355(w_eco355, !a[1], !b[7], !a[7], a[3], b[4], b[6], a[6], !b[3]);
	and _ECO_356(w_eco356, a[1], b[5], !a[5], !b[7], !a[3], a[0], b[3], !b[0]);
	and _ECO_357(w_eco357, !a[1], b[2], b[5], a[5], b[7], !a[7], a[3], b[4], a[4], b[3]);
	and _ECO_358(w_eco358, !a[2], a[1], b[2], !b[7], !a[3], !b[6], b[3], !b[0]);
	and _ECO_359(w_eco359, !a[2], a[1], !b[5], !a[5], b[7], !a[7], b[4], a[4], b[6], !b[3]);
	and _ECO_360(w_eco360, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], a[4], !b[1]);
	and _ECO_361(w_eco361, a[1], b[5], a[5], b[7], b[4], a[4], !a[6], !b[3], !b[0]);
	and _ECO_362(w_eco362, a[1], a[5], !b[7], b[4], !a[6], !b[1], a[0], !b[3], !b[0]);
	and _ECO_363(w_eco363, a[1], b[5], !a[5], !b[7], b[4], !b[6], !b[1], !b[0]);
	and _ECO_364(w_eco364, a[1], !b[7], a[7], b[4], b[6], a[6], !b[0]);
	and _ECO_365(w_eco365, a[1], b[5], a[5], b[7], a[3], b[4], a[4], !a[6], !b[0]);
	and _ECO_366(w_eco366, a[1], b[5], a[5], !a[7], a[3], b[4], a[4], !a[6], !b[1], !b[0]);
	and _ECO_367(w_eco367, !a[2], b[2], !b[7], !a[3], !b[6], !b[1], b[3], !b[0]);
	and _ECO_368(w_eco368, !a[1], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], a[0], !b[0]);
	and _ECO_369(w_eco369, !a[1], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], !b[3], !b[0]);
	and _ECO_370(w_eco370, b[2], !b[5], !b[7], a[7], b[4], b[6], !b[0]);
	and _ECO_371(w_eco371, !a[2], !a[1], b[5], a[5], b[7], !a[7], !a[3], b[4], a[4], !b[3]);
	and _ECO_372(w_eco372, a[2], a[1], !b[2], !b[5], !a[5], !a[7], a[3], b[4], a[4], b[1], !b[0]);
	and _ECO_373(w_eco373, a[1], b[5], b[7], b[4], a[4], !b[6], a[6], !b[3], !b[0]);
	and _ECO_374(w_eco374, !b[5], !b[7], a[7], !a[3], b[4], b[6], !b[1], b[3], !b[0]);
	and _ECO_375(w_eco375, a[2], !a[1], !b[2], b[5], b[7], !a[7], !a[3], b[4], b[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_376(w_eco376, a[1], !b[2], !b[5], !b[7], !a[7], b[4], b[1], a[0], !b[0]);
	and _ECO_377(w_eco377, a[1], !b[2], !b[5], !a[5], !a[7], a[3], b[4], a[4], b[1], !b[3], !b[0]);
	and _ECO_378(w_eco378, !a[2], !a[1], !b[2], !b[5], !b[7], !a[7], b[4], a[0], b[3]);
	and _ECO_379(w_eco379, !a[2], !a[1], b[5], a[5], b[7], !a[7], a[3], b[4], a[4], b[3]);
	and _ECO_380(w_eco380, !a[2], !a[1], !b[2], !b[5], !b[7], !a[7], !a[3], b[4], a[0]);
	and _ECO_381(w_eco381, a[2], a[1], !b[2], b[5], !a[5], !a[4], b[6], b[1], a[0], b[0]);
	and _ECO_382(w_eco382, a[2], b[5], a[5], !a[7], b[4], !a[4], !b[6], a[6], a[0]);
	and _ECO_383(w_eco383, a[2], a[1], !b[2], b[5], b[7], a[7], !a[4], b[6], a[6], b[1], b[0]);
	and _ECO_384(w_eco384, a[2], a[1], !b[2], !a[5], b[4], !a[4], !b[6], !a[6], b[0]);
	and _ECO_385(w_eco385, a[2], !a[1], !b[2], b[5], b[7], a[7], a[3], !a[4], b[6], a[6], !b[3], b[0]);
	and _ECO_386(w_eco386, a[2], !b[2], !b[5], !a[5], b[7], a[7], a[3], b[4], !a[4], !a[6], !b[3], b[0]);
	and _ECO_387(w_eco387, !a[1], b[5], !a[7], !a[3], b[4], !a[4], b[6], a[6], b[1]);
	and _ECO_388(w_eco388, a[1], !b[5], !a[5], !a[7], b[4], !a[4], !b[6], a[6], a[0], !b[0]);
	and _ECO_389(w_eco389, a[2], !b[5], !a[5], !a[7], a[3], a[4], !b[6], a[6]);
	and _ECO_390(w_eco390, !b[5], !b[7], !a[3], b[6], !a[6], !b[1], a[0], b[3]);
	and _ECO_391(w_eco391, a[5], b[7], !b[4], a[4], b[6], !a[6], !a[0]);
	and _ECO_392(w_eco392, b[5], !b[7], !a[7], !b[4], a[4], b[6], !a[6], !a[0], b[0]);
	and _ECO_393(w_eco393, !b[5], !a[5], !a[7], a[3], a[4], !b[6], a[6], b[0]);
	and _ECO_394(w_eco394, a[2], !b[5], !a[5], b[7], !b[4], a[4], b[6], a[6]);
	and _ECO_395(w_eco395, a[2], !b[5], !a[5], b[7], a[3], !b[4], a[4], !b[6], !a[6]);
	and _ECO_396(w_eco396, a[2], !b[2], !a[5], !a[3], b[6], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_397(w_eco397, a[1], b[5], !b[7], !a[7], a[3], !b[4], a[4], b[6], !a[6], !b[1]);
	and _ECO_398(w_eco398, b[5], !a[5], !b[7], !a[7], !a[3], !b[4], a[4], b[3], !b[0]);
	and _ECO_399(w_eco399, !a[2], b[2], a[5], !b[7], !a[7], !b[4], a[4], !b[6], b[1], !b[0]);
	and _ECO_400(w_eco400, !a[2], !a[1], !b[5], !a[5], b[7], !a[7], b[6], !a[6], b[1]);
	and _ECO_401(w_eco401, !a[2], !a[1], b[2], !b[5], !b[7], !a[7], !b[6], !a[6], !b[0]);
	and _ECO_402(w_eco402, !a[2], a[1], b[2], !b[5], !b[7], !b[6], a[6], !b[1], !b[0]);
	and _ECO_403(w_eco403, a[1], !b[5], !b[7], !a[4], b[6], !a[6], !b[0]);
	and _ECO_404(w_eco404, a[1], !b[5], !b[7], b[4], b[6], !a[6], !b[0]);
	and _ECO_405(w_eco405, a[2], a[1], b[5], a[5], !a[7], b[4], a[4], !b[6], a[6], !b[3], !b[0]);
	and _ECO_406(w_eco406, !a[2], !b[2], !b[5], !a[5], b[7], !a[7], a[4], !b[3]);
	and _ECO_407(w_eco407, !a[1], !b[2], !b[5], !b[7], !a[7], a[3], b[4], a[4], !b[6], !b[3]);
	and _ECO_408(w_eco408, b[5], !a[5], b[7], !b[4], a[4], b[6], a[6], b[1], !b[0]);
	and _ECO_409(w_eco409, b[5], !a[5], !b[4], a[4], !b[6], !a[6], b[1], !b[0]);
	and _ECO_410(w_eco410, !b[2], !b[5], !a[5], !a[7], a[4], !b[6], a[6], !b[3]);
	and _ECO_411(w_eco411, !b[5], b[7], !b[4], a[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_412(w_eco412, !a[2], b[2], !b[5], !b[7], !a[7], !b[6], !a[6], b[1], !b[0]);
	and _ECO_413(w_eco413, b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], a[0]);
	and _ECO_414(w_eco414, b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], a[0], b[0]);
	and _ECO_415(w_eco415, a[2], a[1], b[2], a[5], !b[7], !a[7], !a[3], !a[4], b[1], a[0], b[3]);
	and _ECO_416(w_eco416, a[1], !b[7], !a[3], !a[4], !a[6], b[1], a[0], b[3]);
	and _ECO_417(w_eco417, b[2], b[5], b[7], !a[7], !a[3], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_418(w_eco418, b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], !b[3]);
	and _ECO_419(w_eco419, b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], !b[3], b[0]);
	and _ECO_420(w_eco420, a[2], b[2], !b[5], !a[5], !a[7], a[3], !b[4], !a[4], b[1], !b[3]);
	and _ECO_421(w_eco421, b[2], b[5], b[7], !b[4], !a[4], !a[6], b[1], a[0], !b[3]);
	and _ECO_422(w_eco422, b[2], b[5], !a[7], !b[4], !a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_423(w_eco423, !a[1], b[2], b[5], b[7], !a[3], !a[4], !a[6], b[1], b[3]);
	and _ECO_424(w_eco424, b[2], !b[5], !b[7], !a[7], !a[3], !a[4], !a[6], b[1], b[3]);
	and _ECO_425(w_eco425, a[2], b[2], !b[5], !b[7], a[7], a[3], !a[4], b[6]);
	and _ECO_426(w_eco426, a[1], b[2], !b[5], !a[5], b[7], a[7], !a[3], !b[4], !b[1], !a[0], b[3], b[0]);
	and _ECO_427(w_eco427, a[2], b[2], b[5], a[5], b[7], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_428(w_eco428, a[2], a[1], b[2], b[5], !a[5], b[7], !b[4], !a[4], a[6], !b[1], !b[3]);
	and _ECO_429(w_eco429, a[1], b[2], !b[5], !a[5], b[7], !a[7], !b[4], !b[1], !b[3]);
	and _ECO_430(w_eco430, a[2], a[1], b[2], a[5], !b[7], !a[4], !a[6], !b[1], a[0], !b[3]);
	and _ECO_431(w_eco431, a[2], a[1], b[2], b[5], !a[5], !b[7], !b[4], !a[4], !b[6], !b[1], !b[3]);
	and _ECO_432(w_eco432, a[2], b[2], !b[7], a[7], !a[4], b[6], a[6], !b[3]);
	and _ECO_433(w_eco433, a[2], a[1], b[2], b[5], a[5], !a[7], !b[4], !a[4], !a[6], !b[1], !b[3]);
	and _ECO_434(w_eco434, !a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], a[0], b[3]);
	and _ECO_435(w_eco435, !a[1], b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], a[0], b[3], b[0]);
	and _ECO_436(w_eco436, a[2], !a[1], b[2], a[5], !b[7], !a[7], !a[3], !a[4], !b[1], a[0], b[3]);
	and _ECO_437(w_eco437, !a[1], b[2], !b[5], !b[7], a[7], !a[3], !a[4], b[6]);
	and _ECO_438(w_eco438, !a[1], b[2], b[5], b[7], !a[7], !a[3], !a[4], b[6], !a[0], b[0]);
	and _ECO_439(w_eco439, a[2], !a[1], b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], a[0], b[0]);
	and _ECO_440(w_eco440, a[2], !a[1], b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], !b[3], b[0]);
	and _ECO_441(w_eco441, a[2], !a[1], b[2], !b[5], !a[5], !a[7], a[3], !b[4], !a[4], !b[3]);
	and _ECO_442(w_eco442, a[2], !a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_443(w_eco443, a[2], b[2], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[6]);
	and _ECO_444(w_eco444, !a[1], b[2], b[5], !a[7], !a[3], !b[4], !a[4], a[6], a[0], !b[3], b[0]);
	and _ECO_445(w_eco445, !a[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4], b[0]);
	and _ECO_446(w_eco446, !a[2], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1]);
	and _ECO_447(w_eco447, !a[2], b[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], b[0]);
	and _ECO_448(w_eco448, !a[2], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[6], b[1], b[3]);
	and _ECO_449(w_eco449, !a[2], b[2], !a[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], b[0]);
	and _ECO_450(w_eco450, !a[2], a[1], !b[5], !a[5], b[7], !b[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_451(w_eco451, !a[2], a[1], a[5], b[7], !b[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_452(w_eco452, !a[2], a[1], b[5], !b[7], !a[7], !b[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_453(w_eco453, !a[2], !a[1], !b[5], !a[5], !a[7], a[3], !b[4], !a[4], a[0], b[3], b[0]);
	and _ECO_454(w_eco454, !a[2], !a[1], !b[5], !b[7], a[7], !a[4], b[6], b[3]);
	and _ECO_455(w_eco455, !a[1], !b[7], !a[3], !a[4], !a[6], !b[1], a[0], b[3]);
	and _ECO_456(w_eco456, !a[2], !a[1], b[5], b[7], !a[3], !b[4], !a[4], !a[6], a[0], !b[3]);
	and _ECO_457(w_eco457, !a[2], !a[1], !b[5], !a[5], !a[7], !a[3], !b[4], !a[4], a[0], !b[3], b[0]);
	and _ECO_458(w_eco458, a[2], a[1], !b[2], b[5], !a[5], b[7], !a[7], !b[4], !a[4], b[6], b[1], !a[0]);
	and _ECO_459(w_eco459, a[2], !b[2], b[5], !a[5], !b[7], !a[7], !b[4], !a[4], b[6], b[1], b[0]);
	and _ECO_460(w_eco460, a[2], !b[2], !b[5], !b[7], !a[7], !b[4], !a[4], a[6], b[1], !b[3]);
	and _ECO_461(w_eco461, a[2], !b[2], b[5], !a[5], a[7], a[3], !b[4], !a[6], !b[3], b[0]);
	and _ECO_462(w_eco462, a[2], !a[1], b[5], !a[5], b[7], a[3], !b[4], !a[4], !a[6], !b[3], b[0]);
	and _ECO_463(w_eco463, a[2], !a[1], !b[2], !b[5], b[7], !a[3], !b[4], !a[4], b[6], !a[6], b[1]);
	and _ECO_464(w_eco464, !a[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], a[0], b[3]);
	and _ECO_465(w_eco465, !a[2], b[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], a[0], b[3], b[0]);
	and _ECO_466(w_eco466, !a[2], !b[2], !b[5], !b[7], !a[7], !a[4], b[1], a[0], b[3]);
	and _ECO_467(w_eco467, !a[2], !b[5], !b[7], a[7], !a[4], b[6], b[1], b[3]);
	and _ECO_468(w_eco468, !a[2], b[5], b[7], !a[7], !a[3], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_469(w_eco469, !a[2], b[5], b[7], !a[3], !b[4], !a[4], !a[6], b[1], a[0], !b[3]);
	and _ECO_470(w_eco470, !a[2], b[5], !a[7], !a[3], !b[4], !a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_471(w_eco471, !a[2], !b[2], !b[5], !b[7], !a[7], !a[3], !a[4], b[1], a[0]);
	and _ECO_472(w_eco472, !a[2], !b[5], !b[7], a[7], !a[3], !a[4], b[6], b[1]);
	and _ECO_473(w_eco473, !a[2], !a[1], !b[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], !b[3]);
	and _ECO_474(w_eco474, !a[1], !b[2], b[5], !a[5], !b[7], a[7], a[3], !b[4], !a[6], !b[3]);
	and _ECO_475(w_eco475, !a[1], !b[2], b[5], !a[5], !b[7], a[3], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_476(w_eco476, !a[2], a[1], !b[5], !a[5], b[7], a[7], !a[3], !b[4], !b[1], !a[0], b[3], b[0]);
	and _ECO_477(w_eco477, !a[2], !a[1], b[5], b[7], a[3], !b[4], !a[4], !a[6], a[0], b[3]);
	and _ECO_478(w_eco478, !a[2], !a[1], b[5], !a[7], a[3], !b[4], !a[4], a[6], a[0], b[3], b[0]);
	and _ECO_479(w_eco479, !a[2], !a[1], b[5], b[7], !a[7], !a[3], !a[4], b[6], !a[0], b[0]);
	and _ECO_480(w_eco480, !a[1], !b[2], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], a[6], !b[3]);
	and _ECO_481(w_eco481, !a[2], !a[1], b[5], !a[7], !a[3], !b[4], !a[4], a[6], a[0], !b[3], b[0]);
	and _ECO_482(w_eco482, a[2], b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], !b[3]);
	and _ECO_483(w_eco483, a[2], !a[1], b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], a[6], !b[3]);
	and _ECO_484(w_eco484, !a[2], !b[5], !a[5], b[7], !a[7], !b[4], !a[4], !a[6], a[0], !b[3]);
	and _ECO_485(w_eco485, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !b[1]);
	and _ECO_486(w_eco486, a[1], b[5], a[5], b[7], a[3], !b[4], !a[4], !a[6], !b[0]);
	and _ECO_487(w_eco487, a[1], b[5], !a[5], b[7], a[3], !b[4], !a[4], a[6], !b[1], !b[0]);
	and _ECO_488(w_eco488, a[1], b[5], a[5], !a[7], a[3], !b[4], !a[4], !a[6], !b[1], !b[0]);
	and _ECO_489(w_eco489, !a[2], a[1], b[2], !b[5], !a[5], !a[3], !b[4], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_490(w_eco490, a[1], b[5], b[7], !b[4], !a[4], !b[6], a[6], !b[3], !b[0]);
	and _ECO_491(w_eco491, a[1], b[5], b[7], !b[4], !a[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_492(w_eco492, a[1], !a[5], b[7], a[7], !b[4], b[6], a[6], !b[1]);
	and _ECO_493(w_eco493, a[1], !b[5], !a[5], a[7], !b[4], !b[6], !a[6], !b[1]);
	and _ECO_494(w_eco494, !a[2], a[1], b[2], !b[7], !a[4], !b[6], a[6], !b[1], !b[0]);
	and _ECO_495(w_eco495, !a[2], !a[1], b[5], a[5], b[7], !a[7], a[3], !b[4], !a[4], b[3]);
	and _ECO_496(w_eco496, !a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], a[0], !b[0]);
	and _ECO_497(w_eco497, !a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], !b[3], !b[0]);
	and _ECO_498(w_eco498, b[2], !b[5], !b[7], a[7], !a[4], b[6], !b[0]);
	and _ECO_499(w_eco499, !a[2], !a[1], b[5], a[5], b[7], !a[7], !a[3], !b[4], !a[4], !b[3]);
	and _ECO_500(w_eco500, a[1], !b[7], a[7], !a[4], b[6], a[6], !b[0]);
	and _ECO_501(w_eco501, a[2], a[1], !b[2], b[5], a[5], !a[7], !b[4], !a[4], a[6], b[1], !b[3], !b[0]);
	and _ECO_502(w_eco502, a[2], a[1], !b[2], b[5], !a[5], a[7], !b[4], !b[6], !a[6], b[1], !b[3]);
	and _ECO_503(w_eco503, b[5], !a[5], !b[7], !a[7], b[6], a[6], b[1], !b[0]);
	and _ECO_504(w_eco504, a[1], !b[5], !a[5], b[7], !a[7], !b[4], !b[1], !b[3], !b[0]);
	and _ECO_505(w_eco505, !b[5], !b[7], a[7], !a[3], !a[4], b[6], !b[1], b[3], !b[0]);
	and _ECO_506(w_eco506, a[2], !a[1], !b[2], b[5], b[7], !a[7], !a[3], !a[4], b[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_507(w_eco507, a[1], b[5], !a[7], !b[4], !a[4], !b[6], !b[1], !b[3], !b[0]);
	and _ECO_508(w_eco508, a[1], !b[5], !a[5], !a[7], !b[4], !b[6], a[6], !b[1], !b[3]);
	and _ECO_509(w_eco509, a[1], !b[2], a[5], b[7], a[3], !b[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_510(w_eco510, a[1], !b[2], b[5], !b[7], !a[7], a[3], !b[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_511(w_eco511, !a[2], !a[1], !b[2], !b[5], !b[7], !a[7], !a[4], a[0], b[3]);
	and _ECO_512(w_eco512, !a[2], !a[1], !b[2], !b[5], !b[7], !a[7], !a[3], !a[4], a[0]);
	and _ECO_513(w_eco513, b[2], b[5], b[7], a[3], b[4], a[4], !b[6], a[6], b[1]);
	and _ECO_514(w_eco514, a[2], b[2], !b[5], !a[5], b[7], !a[7], a[3], a[4]);
	and _ECO_515(w_eco515, b[2], !b[5], !b[7], !a[7], b[4], !a[6], b[1], a[0]);
	and _ECO_516(w_eco516, b[2], b[5], a[5], b[7], a[3], b[4], a[4], !a[6], b[1]);
	and _ECO_517(w_eco517, a[2], b[2], b[5], !a[5], b[7], a[7], a[3], b[4], a[4], b[6], !a[0], b[3]);
	and _ECO_518(w_eco518, a[2], b[2], b[5], a[5], !a[7], a[3], b[4], a[4], !a[6], !a[0], b[3], b[0]);
	and _ECO_519(w_eco519, a[2], b[2], b[5], !a[7], a[3], b[4], a[4], !b[6], !a[0], b[3], b[0]);
	and _ECO_520(w_eco520, a[2], b[2], b[5], a[5], !a[7], b[4], a[6], b[1], a[0]);
	and _ECO_521(w_eco521, !b[7], !a[7], b[4], b[6], a[6], b[1], a[0]);
	and _ECO_522(w_eco522, a[2], a[1], !b[2], b[5], !a[5], b[7], a[3], b[4], a[4], !a[6], b[1]);
	and _ECO_523(w_eco523, a[1], b[5], b[7], a[3], b[4], a[4], !b[6], a[6], !b[0]);
	and _ECO_524(w_eco524, b[2], b[5], b[7], b[4], b[6], !a[6], b[1], !a[0]);
	and _ECO_525(w_eco525, !b[7], !a[7], !a[3], b[4], b[6], a[6], b[1], b[3]);
	and _ECO_526(w_eco526, a[1], !b[7], !a[3], b[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_527(w_eco527, a[2], b[2], b[5], a[5], !a[7], !a[3], b[4], a[4], !a[6], !a[0], !b[3], b[0]);
	and _ECO_528(w_eco528, a[2], b[2], b[5], !a[7], !a[3], b[4], a[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_529(w_eco529, a[2], b[2], b[5], a[5], b[7], a[3], b[4], a[4], !a[6]);
	and _ECO_530(w_eco530, a[2], a[1], b[2], a[5], !b[7], a[3], b[4], !a[6], !b[1], a[0]);
	and _ECO_531(w_eco531, a[2], a[1], b[2], b[5], !a[5], !b[7], a[3], b[4], a[4], !b[6], !b[1]);
	and _ECO_532(w_eco532, a[2], b[2], b[5], b[7], a[3], b[4], a[4], !b[6], a[6]);
	and _ECO_533(w_eco533, a[2], b[2], !b[7], a[7], a[3], b[4], b[6], a[6]);
	and _ECO_534(w_eco534, a[2], b[2], !b[5], !b[7], a[3], b[4], b[6], !a[6]);
	and _ECO_535(w_eco535, a[1], a[5], b[7], !a[3], a[4], b[6], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_536(w_eco536, a[1], b[5], !b[7], !a[7], !a[3], a[4], b[6], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_537(w_eco537, !a[1], b[2], !b[7], b[4], b[6], a[6], a[0]);
	and _ECO_538(w_eco538, a[2], !a[1], b[2], b[5], a[5], !a[7], b[4], a[6], a[0]);
	and _ECO_539(w_eco539, !a[1], b[2], b[5], !a[5], b[7], a[7], !a[3], b[4], a[4], !a[6], !a[0], b[3]);
	and _ECO_540(w_eco540, b[2], !b[5], !a[5], b[7], a[7], !a[3], a[4], a[6], !b[1], !a[0], b[3]);
	and _ECO_541(w_eco541, !a[1], b[2], !b[7], a[7], !a[3], b[4], b[6], a[6]);
	and _ECO_542(w_eco542, !a[1], b[2], !b[5], !b[7], !a[3], b[4], b[6], !a[6]);
	and _ECO_543(w_eco543, !a[1], !b[5], !b[7], !a[7], a[3], b[4], !b[6], !a[6], !b[3]);
	and _ECO_544(w_eco544, !a[1], b[2], b[5], b[7], !a[3], b[4], a[4], !a[6], a[0], !b[3]);
	and _ECO_545(w_eco545, !a[1], b[2], b[5], !a[5], b[7], a[7], !a[3], b[4], a[4], b[6], !b[1], !a[0]);
	and _ECO_546(w_eco546, !a[2], a[1], b[2], !b[5], !a[5], a[7], !a[3], !b[6], a[6], b[3]);
	and _ECO_547(w_eco547, !a[2], a[1], !b[5], b[7], a[3], a[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_548(w_eco548, !a[2], a[1], b[5], !b[7], a[3], b[6], !a[6], !b[1], a[0], b[0]);
	and _ECO_549(w_eco549, a[1], b[5], a[5], b[7], a[4], b[6], !a[6], !b[1], !b[3]);
	and _ECO_550(w_eco550, !a[2], a[1], !a[5], a[7], a[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_551(w_eco551, a[1], b[5], a[5], b[7], a[3], a[4], b[6], !a[6], !b[1]);
	and _ECO_552(w_eco552, !a[2], a[1], b[5], !a[5], !b[7], a[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_553(w_eco553, !a[2], !a[1], b[5], b[7], a[3], b[4], a[4], !b[6], a[6], b[3]);
	and _ECO_554(w_eco554, !a[2], !a[1], b[5], a[5], b[7], a[3], b[4], a[4], !a[6], b[3]);
	and _ECO_555(w_eco555, !a[2], !a[1], b[5], !a[5], b[7], a[7], b[4], a[4], b[6], !b[1], !a[0], b[3]);
	and _ECO_556(w_eco556, !a[2], !a[1], !b[7], a[7], b[4], b[6], a[6], b[3]);
	and _ECO_557(w_eco557, !a[2], !a[1], b[5], a[5], !a[7], a[3], b[4], a[4], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_558(w_eco558, !a[2], !a[1], b[5], !b[7], a[3], b[4], a[4], !b[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_559(w_eco559, !a[2], !a[1], !b[5], !b[7], b[4], b[6], !a[6], b[3]);
	and _ECO_560(w_eco560, !a[2], !a[1], b[5], b[7], !a[3], b[4], !b[6], a[6], b[1]);
	and _ECO_561(w_eco561, !a[2], !b[5], b[7], a[3], a[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_562(w_eco562, !a[2], !a[1], b[5], !a[5], !b[7], a[3], b[4], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_563(w_eco563, !a[2], !a[1], b[5], !a[5], !b[7], a[3], b[4], a[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_564(w_eco564, !a[2], b[5], a[5], b[7], a[3], a[4], b[6], !a[6]);
	and _ECO_565(w_eco565, !a[2], !a[1], !b[7], a[3], b[4], !b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_566(w_eco566, !a[2], !a[1], b[5], b[7], !a[3], b[4], a[4], !b[6], a[6], !b[3]);
	and _ECO_567(w_eco567, !a[2], !a[1], b[5], a[5], b[7], !a[3], b[4], a[4], !a[6], !b[3]);
	and _ECO_568(w_eco568, !a[2], !a[1], b[5], a[5], !a[7], !a[3], b[4], a[4], !a[6], !b[1], !a[0], !b[3], b[0]);
	and _ECO_569(w_eco569, !a[2], !a[1], b[5], !b[7], !a[3], b[4], a[4], !b[6], !b[1], !a[0], !b[3], b[0]);
	and _ECO_570(w_eco570, a[1], b[5], !a[7], a[3], b[4], a[4], b[6], a[6], b[1], a[0], b[3]);
	and _ECO_571(w_eco571, a[2], a[1], !b[2], !a[5], a[7], !a[3], !a[6], a[0], b[3], b[0]);
	and _ECO_572(w_eco572, a[2], a[1], !b[2], b[5], b[7], b[4], a[4], b[6], a[6], b[1], b[0]);
	and _ECO_573(w_eco573, a[2], !b[2], !b[5], !a[5], b[7], !a[7], !a[3], b[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_574(w_eco574, a[2], a[1], !b[2], !b[5], !a[5], a[7], !a[3], !b[6], !a[0], b[3], b[0]);
	and _ECO_575(w_eco575, a[2], !a[1], !b[2], b[5], b[7], a[7], a[3], b[4], b[6], a[6], !b[3], b[0]);
	and _ECO_576(w_eco576, a[2], !a[1], b[5], b[7], a[3], b[4], a[4], !b[6], !a[6], !b[3], b[0]);
	and _ECO_577(w_eco577, a[2], !a[1], b[5], !a[7], a[3], b[4], a[4], b[6], a[6], !b[3], b[0]);
	and _ECO_578(w_eco578, !a[1], !b[2], !b[5], a[5], b[7], a[3], a[4], b[6], !a[6], !b[3]);
	and _ECO_579(w_eco579, a[2], !b[2], !a[5], b[7], a[7], a[3], b[6], a[6], !b[3], b[0]);
	and _ECO_580(w_eco580, a[2], !b[2], !b[5], !a[5], b[7], a[7], a[3], !b[6], !a[6], !b[3], b[0]);
	and _ECO_581(w_eco581, a[2], a[1], !b[2], b[5], !a[5], a[7], !a[6], a[0], b[0]);
	and _ECO_582(w_eco582, a[2], a[1], !b[2], b[5], !a[5], a[7], a[4], !a[6], b[0]);
	and _ECO_583(w_eco583, a[1], !b[2], b[5], !b[7], !a[7], a[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_584(w_eco584, a[2], a[1], !b[2], b[5], !a[5], a[4], b[6], !a[6], b[0]);
	and _ECO_585(w_eco585, a[1], !b[5], !a[5], b[7], a[3], a[4], b[6], a[6], !b[1]);
	and _ECO_586(w_eco586, a[2], a[1], !b[2], !b[5], !a[5], b[7], a[3], !b[6], !a[6], !b[1], b[0]);
	and _ECO_587(w_eco587, a[2], a[1], !b[5], !a[5], b[7], a[4], b[6], a[6], !b[1]);
	and _ECO_588(w_eco588, a[1], !b[2], a[5], b[7], a[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_589(w_eco589, a[2], a[1], !b[2], !b[5], !a[5], b[7], !b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_590(w_eco590, a[2], !b[2], b[5], !a[5], a[7], !a[6], !b[1], a[0], b[0]);
	and _ECO_591(w_eco591, a[2], !a[1], !b[2], b[5], !a[5], b[4], !a[6], !b[1], a[0], b[0]);
	and _ECO_592(w_eco592, a[2], !b[2], b[5], !a[5], a[7], a[4], !a[6], !b[1], b[0]);
	and _ECO_593(w_eco593, !a[1], b[5], !a[5], b[7], !a[7], a[3], b[4], a[4], !a[6], !b[1], b[3], b[0]);
	and _ECO_594(w_eco594, a[2], !a[1], !b[2], b[5], b[7], b[4], a[4], b[6], a[6], !b[1], b[0]);
	and _ECO_595(w_eco595, a[2], !a[1], !b[2], !a[5], !a[3], b[4], !b[6], !a[6], !b[1], b[3], b[0]);
	and _ECO_596(w_eco596, !a[1], b[5], !a[5], b[7], !a[7], !a[3], b[4], a[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_597(w_eco597, !a[2], !b[2], b[5], !a[5], b[7], a[7], a[3], b[4], a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_598(w_eco598, !a[2], !b[7], a[7], b[4], b[6], a[6], b[1], b[3]);
	and _ECO_599(w_eco599, !a[2], !b[2], b[5], a[5], !a[7], a[3], b[4], a[4], !a[6], b[1], !a[0], b[3], b[0]);
	and _ECO_600(w_eco600, !a[2], !b[2], b[5], !a[7], a[3], b[4], a[4], !b[6], b[1], !a[0], b[3], b[0]);
	and _ECO_601(w_eco601, !a[2], !b[5], !b[7], b[4], b[6], !a[6], b[1], b[3]);
	and _ECO_602(w_eco602, !a[2], !b[2], b[5], a[5], !a[7], !a[3], b[4], a[6], b[1], a[0]);
	and _ECO_603(w_eco603, !a[2], b[5], b[7], !a[3], b[4], b[6], !a[6], b[1], !a[0]);
	and _ECO_604(w_eco604, !a[2], !b[2], !b[5], b[7], a[3], a[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_605(w_eco605, a[1], !b[2], b[5], !a[5], !b[7], a[3], b[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_606(w_eco606, !b[2], b[5], !a[5], !b[7], a[3], b[4], a[4], !a[6], b[1], !b[3], b[0]);
	and _ECO_607(w_eco607, !a[2], b[5], b[7], !a[3], b[4], a[4], !b[6], a[6], b[1], !b[3]);
	and _ECO_608(w_eco608, !a[2], !b[5], !b[7], !a[7], !a[3], b[4], !a[6], b[1], a[0]);
	and _ECO_609(w_eco609, !a[2], !b[7], a[7], !a[3], b[4], b[6], a[6], b[1]);
	and _ECO_610(w_eco610, !a[2], !b[2], b[5], a[5], !a[7], !a[3], b[4], a[4], !a[6], b[1], !a[0], !b[3], b[0]);
	and _ECO_611(w_eco611, !a[2], !b[2], b[5], !a[7], !a[3], b[4], a[4], !b[6], b[1], !a[0], !b[3], b[0]);
	and _ECO_612(w_eco612, !a[2], !b[5], !b[7], !a[3], b[4], b[6], !a[6], b[1]);
	and _ECO_613(w_eco613, !b[2], b[5], !a[5], !b[7], a[7], a[3], a[4], !b[6], !b[3]);
	and _ECO_614(w_eco614, !a[1], !b[2], !b[7], !a[7], a[3], b[4], a[4], !b[6], !a[6], !b[3]);
	and _ECO_615(w_eco615, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], b[4], a[6], a[0]);
	and _ECO_616(w_eco616, !a[2], !b[5], !a[5], b[7], a[7], !a[3], a[4], a[6], !b[1], !a[0], b[3]);
	and _ECO_617(w_eco617, !a[2], !a[1], b[5], !a[5], b[7], a[7], !a[3], b[4], a[4], b[6], !b[1], !a[0]);
	and _ECO_618(w_eco618, !a[2], !a[1], !b[7], a[7], !a[3], b[4], b[6], a[6]);
	and _ECO_619(w_eco619, !a[2], !a[1], !b[5], !b[7], !a[3], b[4], b[6], !a[6]);
	and _ECO_620(w_eco620, a[2], b[2], b[5], a[5], !a[7], a[3], b[4], a[4], !b[6], !a[0], b[3]);
	and _ECO_621(w_eco621, a[2], a[1], b[5], a[5], b[7], !a[7], b[4], a[6], a[0], !b[0]);
	and _ECO_622(w_eco622, a[1], b[5], !a[5], b[7], !a[3], b[4], a[4], !a[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_623(w_eco623, a[1], b[5], a[5], b[7], !a[7], b[4], b[6], !a[0], !b[0]);
	and _ECO_624(w_eco624, !a[1], b[2], b[5], a[5], b[7], !a[7], !a[3], b[4], b[6], !a[0]);
	and _ECO_625(w_eco625, !a[1], b[2], b[5], !a[5], b[7], !a[3], b[4], a[4], !a[6], !a[0], b[3], !b[0]);
	and _ECO_626(w_eco626, b[5], !a[5], !b[7], !a[7], !a[3], a[6], !b[1], b[3], !b[0]);
	and _ECO_627(w_eco627, !a[2], !b[5], !a[5], b[7], !a[7], a[3], b[4], a[4], !a[6], a[0]);
	and _ECO_628(w_eco628, !a[2], a[1], b[2], !b[5], !a[5], !a[7], !a[3], b[4], a[6], b[1], !a[0], b[3], !b[0]);
	and _ECO_629(w_eco629, a[1], b[5], b[7], a[3], b[4], a[4], b[6], !a[6], !b[0]);
	and _ECO_630(w_eco630, !a[2], a[1], b[2], !b[7], b[4], !b[6], a[6], !b[1], !b[0]);
	and _ECO_631(w_eco631, a[1], !b[5], !a[5], b[7], !a[7], a[4], a[6], !b[1], a[0], !b[0]);
	and _ECO_632(w_eco632, !a[2], b[2], !b[5], !a[5], !a[3], a[4], !b[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_633(w_eco633, a[1], b[5], a[5], !a[7], b[4], a[4], !a[6], !b[1], !b[3], !b[0]);
	and _ECO_634(w_eco634, a[1], !b[5], !a[5], b[7], !a[7], a[4], !b[1], !b[3], !b[0]);
	and _ECO_635(w_eco635, a[1], b[5], b[7], b[4], a[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_636(w_eco636, a[1], b[5], !a[7], b[4], a[4], !b[6], !b[1], !b[3], !b[0]);
	and _ECO_637(w_eco637, !a[2], b[2], !b[5], !a[5], !a[3], !b[6], a[6], !b[1], b[3], !b[0]);
	and _ECO_638(w_eco638, b[2], b[5], b[7], a[3], b[4], a[4], !b[6], a[6], !b[0]);
	and _ECO_639(w_eco639, b[2], !b[5], !b[7], b[4], b[6], !a[6], !b[0]);
	and _ECO_640(w_eco640, b[2], !b[7], a[7], b[4], b[6], a[6], !b[0]);
	and _ECO_641(w_eco641, !a[2], !b[5], !a[5], b[7], !a[7], b[4], a[4], !a[6], a[0], !b[3]);
	and _ECO_642(w_eco642, a[2], a[1], b[5], a[5], !a[7], a[3], b[4], a[4], !b[6], a[6], !b[0]);
	and _ECO_643(w_eco643, a[1], b[5], b[7], b[4], b[6], !a[6], !a[0], !b[0]);
	and _ECO_644(w_eco644, a[1], !b[5], !a[5], b[7], !a[7], a[3], a[4], !b[1], !b[0]);
	and _ECO_645(w_eco645, a[2], !a[1], !b[2], !b[5], b[7], a[3], a[4], b[6], !a[6], !b[0]);
	and _ECO_646(w_eco646, a[2], b[5], a[5], b[7], !a[7], !a[3], b[4], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_647(w_eco647, b[5], b[7], !a[3], b[4], b[6], !a[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_648(w_eco648, !b[7], a[7], !a[3], b[4], b[6], a[6], !b[1], b[3], !b[0]);
	and _ECO_649(w_eco649, !b[5], !b[7], !a[3], b[4], b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_650(w_eco650, b[5], a[5], b[7], a[3], a[4], b[6], !a[6], !b[0]);
	and _ECO_651(w_eco651, a[2], !b[5], !a[5], b[7], !a[7], a[3], a[4], !b[0]);
	and _ECO_652(w_eco652, a[2], !a[1], !b[2], !b[5], b[7], a[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_653(w_eco653, !a[2], !b[2], !b[5], !a[5], b[7], !a[7], a[3], a[4]);
	and _ECO_654(w_eco654, !a[2], !b[2], b[5], a[5], !a[7], a[3], b[4], a[4], !b[6], b[1], !a[0], b[3]);
	and _ECO_655(w_eco655, a[1], !b[2], b[5], a[5], !a[7], a[3], b[4], a[4], a[6], b[1], !b[3], !b[0]);
	and _ECO_656(w_eco656, !a[2], !b[2], b[5], a[5], !a[7], !a[3], b[4], a[4], !b[6], b[1], !a[0], !b[3]);
	and _ECO_657(w_eco657, a[1], b[5], !a[7], a[3], b[4], a[4], !b[6], !b[1], !b[0]);
	and _ECO_658(w_eco658, a[1], !b[5], !a[5], !a[7], a[3], a[4], !b[6], a[6], !b[1]);
	and _ECO_659(w_eco659, a[1], !b[2], b[5], a[5], b[7], !a[7], b[4], a[6], a[0], !b[0]);
	and _ECO_660(w_eco660, !a[2], !a[1], !b[2], b[5], a[5], !a[7], b[4], a[6], a[0], b[3]);
	and _ECO_661(w_eco661, !a[2], !a[1], !b[2], b[5], a[5], !a[7], a[3], b[4], a[4], !b[6], !a[0], b[3]);
	and _ECO_662(w_eco662, !a[2], !a[5], a[7], !a[3], a[4], !b[6], !a[6], !b[1], !a[0], b[3]);
	and _ECO_663(w_eco663, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], b[4], a[4], !b[6], !a[0], !b[3]);
	and _ECO_664(w_eco664, a[2], !a[1], b[2], b[5], a[5], !a[7], !a[4], !b[6], a[6], b[1]);
	and _ECO_665(w_eco665, a[1], !b[5], !b[7], !a[3], b[6], !a[6], a[0], b[3]);
	and _ECO_666(w_eco666, !a[5], !b[7], !a[3], b[6], !a[6], !b[1], a[0], b[3]);
	and _ECO_667(w_eco667, a[2], !a[1], !b[5], !a[5], !a[7], !b[6], a[6], b[1]);
	and _ECO_668(w_eco668, a[1], !b[5], !a[5], b[7], !a[7], !a[3], !b[4], a[4], a[6], a[0], b[3], !b[0]);
	and _ECO_669(w_eco669, !a[2], a[1], b[2], !b[5], !a[5], !a[3], !b[4], a[4], !b[6], b[3], !b[0]);
	and _ECO_670(w_eco670, !b[5], b[7], a[3], !b[4], a[4], b[6], !a[6], !b[0]);
	and _ECO_671(w_eco671, !b[2], !b[5], !a[5], !a[7], a[3], a[4], !b[6], a[6]);
	and _ECO_672(w_eco672, a[2], b[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4]);
	and _ECO_673(w_eco673, b[2], !b[5], !b[7], !a[7], !a[4], !a[6], b[1], a[0]);
	and _ECO_674(w_eco674, b[2], b[5], a[5], b[7], a[3], !b[4], !a[4], !a[6], b[1]);
	and _ECO_675(w_eco675, a[2], b[2], b[5], !a[5], b[7], a[7], a[3], !b[4], !a[4], b[6], !a[0], b[3]);
	and _ECO_676(w_eco676, a[2], b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], !a[6], !a[0], b[3], b[0]);
	and _ECO_677(w_eco677, a[2], b[2], b[5], !a[7], a[3], !b[4], !a[4], !b[6], !a[0], b[3], b[0]);
	and _ECO_678(w_eco678, a[2], b[2], b[5], a[5], !a[7], !a[4], a[6], b[1], a[0]);
	and _ECO_679(w_eco679, !b[7], !a[7], !a[4], b[6], a[6], b[1], a[0]);
	and _ECO_680(w_eco680, b[2], b[5], b[7], !a[4], b[6], !a[6], b[1], !a[0]);
	and _ECO_681(w_eco681, !b[7], !a[7], !a[3], !a[4], b[6], a[6], b[1], b[3]);
	and _ECO_682(w_eco682, a[1], !b[7], !a[3], !a[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_683(w_eco683, a[2], b[2], !b[5], !a[5], b[7], !a[7], !b[4], !b[3]);
	and _ECO_684(w_eco684, a[2], b[2], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !a[6], !a[0], !b[3], b[0]);
	and _ECO_685(w_eco685, a[2], b[2], b[5], !a[7], !a[3], !b[4], !a[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_686(w_eco686, !a[1], b[2], !b[5], !b[7], !a[4], b[6], !a[6], b[3]);
	and _ECO_687(w_eco687, !a[1], b[2], !b[5], !b[7], !a[3], !a[4], b[6], !a[6]);
	and _ECO_688(w_eco688, a[2], b[2], b[5], a[5], b[7], a[3], !b[4], !a[4], !a[6]);
	and _ECO_689(w_eco689, a[2], a[1], b[2], a[5], !b[7], a[3], !a[4], !a[6], !b[1], a[0]);
	and _ECO_690(w_eco690, a[2], a[1], b[2], b[5], !a[5], !b[7], a[3], !b[4], !a[4], !b[6], !b[1]);
	and _ECO_691(w_eco691, a[2], b[2], !b[7], a[7], a[3], !a[4], b[6], a[6]);
	and _ECO_692(w_eco692, a[1], a[5], b[7], !a[3], !b[4], b[6], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_693(w_eco693, a[1], b[5], !b[7], !a[7], !a[3], !b[4], b[6], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_694(w_eco694, a[2], b[2], !b[5], !b[7], a[3], !a[4], b[6], !a[6]);
	and _ECO_695(w_eco695, a[2], a[1], b[5], !a[5], b[7], a[3], !b[4], !a[4], b[6], !a[6]);
	and _ECO_696(w_eco696, a[2], b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], !b[6], a[6]);
	and _ECO_697(w_eco697, a[2], b[2], !b[5], !b[7], !a[4], b[6], !a[6], !b[3]);
	and _ECO_698(w_eco698, a[2], !a[1], b[2], b[5], a[5], !a[7], !a[4], a[6], a[0]);
	and _ECO_699(w_eco699, !a[1], !b[7], !a[7], !a[4], b[6], a[6], a[0]);
	and _ECO_700(w_eco700, !a[1], b[2], b[5], !a[5], b[7], a[7], !a[3], !b[4], !a[4], !a[6], !a[0], b[3]);
	and _ECO_701(w_eco701, b[2], !b[5], !a[5], b[7], a[7], !a[3], !b[4], a[6], !b[1], !a[0], b[3]);
	and _ECO_702(w_eco702, !a[1], b[2], !b[7], a[7], !a[3], !a[4], b[6], a[6]);
	and _ECO_703(w_eco703, !a[1], b[2], b[5], b[7], !a[3], !b[4], !a[4], !a[6], a[0], !b[3]);
	and _ECO_704(w_eco704, !a[1], b[2], b[5], b[7], !a[3], !b[4], !a[4], !b[6], a[6], !b[3]);
	and _ECO_705(w_eco705, !a[1], b[2], b[5], !a[5], b[7], a[7], !a[3], !b[4], !a[4], b[6], !b[1], !a[0]);
	and _ECO_706(w_eco706, !a[2], a[1], !b[5], b[7], a[3], !b[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_707(w_eco707, !a[2], a[1], !a[5], a[7], !b[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_708(w_eco708, !a[2], a[1], b[5], !a[5], !b[7], !b[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_709(w_eco709, a[1], b[5], a[5], b[7], a[3], !b[4], b[6], !a[6], !b[1]);
	and _ECO_710(w_eco710, a[1], !b[5], !a[5], !a[7], a[3], !b[4], !b[6], a[6], !b[1]);
	and _ECO_711(w_eco711, !a[2], !a[1], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[6], b[3]);
	and _ECO_712(w_eco712, !a[2], !a[1], b[5], a[5], b[7], a[3], !b[4], !a[4], !a[6], b[3]);
	and _ECO_713(w_eco713, !a[2], !a[1], b[5], !a[5], b[7], a[7], !b[4], !a[4], b[6], !b[1], !a[0], b[3]);
	and _ECO_714(w_eco714, !a[2], !a[1], !b[7], a[7], !a[4], b[6], a[6], b[3]);
	and _ECO_715(w_eco715, !a[2], !a[1], b[5], a[5], !a[7], a[3], !b[4], !a[4], !a[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_716(w_eco716, !a[2], !a[1], b[5], !b[7], a[3], !b[4], !a[4], !b[6], !b[1], !a[0], b[3], b[0]);
	and _ECO_717(w_eco717, !a[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_718(w_eco718, !a[2], !a[1], b[5], !a[5], !b[7], a[3], !a[4], !a[6], !b[1], a[0], !b[3], b[0]);
	and _ECO_719(w_eco719, !a[1], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], !b[6], a[0], b[0]);
	and _ECO_720(w_eco720, !a[2], !a[1], b[5], !a[5], !b[7], a[3], !b[4], !a[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_721(w_eco721, !a[1], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], a[6], !b[3], b[0]);
	and _ECO_722(w_eco722, !a[2], !a[1], b[5], a[5], b[7], !a[3], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_723(w_eco723, !a[2], !a[1], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !a[6], !b[1], !a[0], !b[3], b[0]);
	and _ECO_724(w_eco724, !a[2], !a[1], b[5], !b[7], !a[3], !b[4], !a[4], !b[6], !b[1], !a[0], !b[3], b[0]);
	and _ECO_725(w_eco725, a[2], !b[2], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], a[6], b[1]);
	and _ECO_726(w_eco726, a[2], a[1], !b[2], b[5], b[7], !a[3], !b[4], !a[4], b[6], b[1], a[0], b[3], b[0]);
	and _ECO_727(w_eco727, a[2], !b[2], !b[5], !a[5], b[7], !a[7], !a[3], !a[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_728(w_eco728, a[2], !a[1], b[5], b[7], a[3], !b[4], !a[4], !b[6], !a[6], !b[3], b[0]);
	and _ECO_729(w_eco729, a[2], !a[1], b[5], !a[7], a[3], !b[4], !a[4], b[6], a[6], !b[3], b[0]);
	and _ECO_730(w_eco730, !a[1], !b[2], !b[5], a[5], b[7], a[3], !b[4], b[6], !a[6], !b[3]);
	and _ECO_731(w_eco731, a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[3], a[6], b[1]);
	and _ECO_732(w_eco732, a[2], !a[1], !b[5], !a[5], b[7], !a[7], !a[3], !b[6], b[1]);
	and _ECO_733(w_eco733, a[2], a[1], !b[2], b[5], !a[5], a[7], !b[4], !a[6], b[0]);
	and _ECO_734(w_eco734, a[1], !b[2], a[5], b[7], !b[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_735(w_eco735, a[1], !b[2], b[5], !b[7], !a[7], !b[4], b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_736(w_eco736, a[1], !b[5], !a[5], b[7], a[3], !b[4], b[6], a[6], !b[1]);
	and _ECO_737(w_eco737, a[2], a[1], !b[2], b[5], !a[5], !b[4], b[6], !a[6], b[0]);
	and _ECO_738(w_eco738, a[2], a[1], !b[5], !a[5], b[7], !b[4], b[6], a[6], !b[1]);
	and _ECO_739(w_eco739, a[2], !a[1], !b[2], b[5], !a[5], !a[4], !a[6], !b[1], a[0], b[0]);
	and _ECO_740(w_eco740, a[2], !b[2], b[5], !a[5], a[7], !b[4], !a[6], !b[1], b[0]);
	and _ECO_741(w_eco741, !a[1], b[5], !a[5], b[7], !a[7], a[3], !b[4], !a[4], !a[6], !b[1], b[3], b[0]);
	and _ECO_742(w_eco742, a[2], !a[1], !b[2], b[5], !a[3], !a[4], !a[6], !b[1], a[0], b[3], b[0]);
	and _ECO_743(w_eco743, a[2], !a[1], !b[2], b[5], b[7], !b[4], !a[4], b[6], a[6], !b[1], b[0]);
	and _ECO_744(w_eco744, a[2], !a[1], !b[2], !a[5], !a[3], !a[4], !b[6], !a[6], !b[1], b[3], b[0]);
	and _ECO_745(w_eco745, !a[1], b[5], !a[5], b[7], !a[7], !a[3], !b[4], !a[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_746(w_eco746, !a[2], b[5], a[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], b[3]);
	and _ECO_747(w_eco747, !a[2], !b[2], b[5], !a[5], b[7], a[7], a[3], !b[4], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_748(w_eco748, !a[2], !b[7], a[7], !a[4], b[6], a[6], b[1], b[3]);
	and _ECO_749(w_eco749, !a[2], !b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], !a[6], b[1], !a[0], b[3], b[0]);
	and _ECO_750(w_eco750, !a[2], !b[2], b[5], !a[7], a[3], !b[4], !a[4], !b[6], b[1], !a[0], b[3], b[0]);
	and _ECO_751(w_eco751, !a[2], !b[2], b[5], a[5], !a[7], !a[3], !a[4], a[6], b[1], a[0]);
	and _ECO_752(w_eco752, !a[2], b[5], b[7], !a[3], !a[4], b[6], !a[6], b[1], !a[0]);
	and _ECO_753(w_eco753, !a[2], !a[1], b[5], b[7], !a[3], !a[4], !b[6], b[1], b[3]);
	and _ECO_754(w_eco754, !a[2], !b[5], !b[7], !a[3], !a[4], b[6], !a[6], b[1]);
	and _ECO_755(w_eco755, !a[2], !b[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_756(w_eco756, a[1], !b[2], b[5], !a[5], !b[7], a[3], !a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_757(w_eco757, !b[2], !b[5], !b[7], !a[7], !a[4], !b[6], b[1], a[0]);
	and _ECO_758(w_eco758, !b[2], b[5], !a[5], !b[7], a[3], !b[4], !a[4], !a[6], b[1], !b[3], b[0]);
	and _ECO_759(w_eco759, !b[2], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], a[6], b[1], !b[3]);
	and _ECO_760(w_eco760, !a[2], b[5], b[7], !a[3], !b[4], !a[4], !b[6], a[6], b[1], !b[3]);
	and _ECO_761(w_eco761, !a[2], !b[7], a[7], !a[3], !a[4], b[6], a[6], b[1]);
	and _ECO_762(w_eco762, !a[2], !b[2], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !a[6], b[1], !a[0], !b[3], b[0]);
	and _ECO_763(w_eco763, !a[2], !b[2], b[5], !a[7], !a[3], !b[4], !a[4], !b[6], b[1], !a[0], !b[3], b[0]);
	and _ECO_764(w_eco764, !a[2], !a[1], !b[5], !b[7], !a[4], b[6], !a[6], b[3]);
	and _ECO_765(w_eco765, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], !a[4], a[6], a[0]);
	and _ECO_766(w_eco766, !a[2], !b[5], !a[5], b[7], a[7], !a[3], !b[4], a[6], !b[1], !a[0], b[3]);
	and _ECO_767(w_eco767, !a[2], !a[1], b[5], b[7], !a[3], !b[4], !a[4], !b[6], a[6], !b[3]);
	and _ECO_768(w_eco768, !a[2], !a[1], b[5], !a[5], b[7], a[7], !a[3], !b[4], !a[4], b[6], !b[1], !a[0]);
	and _ECO_769(w_eco769, !a[2], !a[1], !b[7], a[7], !a[3], !a[4], b[6], a[6]);
	and _ECO_770(w_eco770, a[2], b[2], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !b[6], !a[0], !b[3]);
	and _ECO_771(w_eco771, a[2], a[1], b[5], a[5], b[7], !a[7], !a[4], a[6], a[0], !b[0]);
	and _ECO_772(w_eco772, a[1], b[5], !a[5], b[7], !a[3], !b[4], !a[4], !a[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_773(w_eco773, a[1], b[5], a[5], b[7], !a[7], !a[4], b[6], !a[0], !b[0]);
	and _ECO_774(w_eco774, !a[1], b[2], b[5], a[5], b[7], !a[7], !a[3], !a[4], b[6], !a[0]);
	and _ECO_775(w_eco775, !a[1], b[2], b[5], !a[5], b[7], !a[3], !b[4], !a[4], !a[6], !a[0], b[3], !b[0]);
	and _ECO_776(w_eco776, !a[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !a[4], !a[6], a[0]);
	and _ECO_777(w_eco777, !a[2], a[1], b[2], !b[5], !a[5], !a[7], !a[3], !a[4], a[6], b[1], !a[0], b[3], !b[0]);
	and _ECO_778(w_eco778, !a[2], !b[5], !a[5], b[7], !a[7], !b[4], !a[4], b[6], a[0], !b[3]);
	and _ECO_779(w_eco779, !a[2], a[1], !b[5], !a[5], b[7], !a[7], !a[4], b[6], !a[0], !b[3]);
	and _ECO_780(w_eco780, !a[2], a[1], !b[5], !a[5], b[7], !a[7], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_781(w_eco781, a[1], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[6], !b[0]);
	and _ECO_782(w_eco782, a[1], b[5], b[7], a[3], !b[4], !a[4], b[6], !a[6], !b[0]);
	and _ECO_783(w_eco783, b[2], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[6], !b[0]);
	and _ECO_784(w_eco784, b[2], !b[5], !b[7], !a[4], b[6], !a[6], !b[0]);
	and _ECO_785(w_eco785, b[2], !b[7], a[7], !a[4], b[6], a[6], !b[0]);
	and _ECO_786(w_eco786, a[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !b[0]);
	and _ECO_787(w_eco787, a[2], a[1], !b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], !b[0]);
	and _ECO_788(w_eco788, a[1], b[5], b[7], !a[4], b[6], !a[6], !a[0], !b[0]);
	and _ECO_789(w_eco789, a[1], b[5], !a[7], a[3], !b[4], !a[4], !b[6], !b[1], !b[0]);
	and _ECO_790(w_eco790, a[2], !a[1], !b[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], !b[0]);
	and _ECO_791(w_eco791, b[5], a[5], b[7], a[3], !b[4], b[6], !a[6], !b[0]);
	and _ECO_792(w_eco792, a[2], b[5], a[5], b[7], !a[7], !a[3], !a[4], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_793(w_eco793, b[5], b[7], !a[3], !a[4], b[6], !a[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_794(w_eco794, !a[2], b[2], !a[5], !a[3], !b[4], !b[6], !a[6], !b[1], !a[0], b[3], !b[0]);
	and _ECO_795(w_eco795, !b[7], a[7], !a[3], !a[4], b[6], a[6], !b[1], b[3], !b[0]);
	and _ECO_796(w_eco796, !b[5], !b[7], !a[3], !a[4], b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_797(w_eco797, a[2], !a[1], !b[2], !b[5], b[7], !b[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_798(w_eco798, a[2], !b[5], !a[5], b[7], !a[7], !b[4], !b[3], !b[0]);
	and _ECO_799(w_eco799, !a[2], !b[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4]);
	and _ECO_800(w_eco800, !a[2], !b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], !b[6], b[1], !a[0], b[3]);
	and _ECO_801(w_eco801, a[1], !b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], a[6], b[1], !b[3], !b[0]);
	and _ECO_802(w_eco802, !a[2], !b[2], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !b[6], b[1], !a[0], !b[3]);
	and _ECO_803(w_eco803, !b[2], !b[5], !a[5], !a[7], !b[4], !b[6], a[6], !b[3]);
	and _ECO_804(w_eco804, !a[2], !a[1], !b[5], !b[7], !a[3], !a[4], b[6], !a[6]);
	and _ECO_805(w_eco805, a[1], !b[2], b[5], a[5], b[7], !a[7], !a[4], a[6], a[0], !b[0]);
	and _ECO_806(w_eco806, !a[2], !a[1], !b[2], b[5], a[5], !a[7], a[3], !b[4], !a[4], !b[6], !a[0], b[3]);
	and _ECO_807(w_eco807, !a[2], !a[5], a[7], !a[3], !b[4], !b[6], !a[6], !b[1], !a[0], b[3]);
	and _ECO_808(w_eco808, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], !b[4], !a[4], !b[6], !a[0], !b[3]);
	and _ECO_809(w_eco809, a[2], b[2], !b[5], !a[5], b[7], a[3], a[4], b[6], a[6], !a[0], b[3]);
	and _ECO_810(w_eco810, a[2], b[2], !b[5], !a[5], b[7], a[3], a[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_811(w_eco811, a[2], b[2], b[5], a[5], b[7], b[4], !b[6], a[6], b[1], a[0]);
	and _ECO_812(w_eco812, a[1], !b[5], !a[5], a[7], !a[3], !b[6], a[6], !a[0], b[3]);
	and _ECO_813(w_eco813, b[2], !b[5], !b[7], b[4], b[6], !a[6], b[1]);
	and _ECO_814(w_eco814, !b[7], !a[7], a[3], b[4], b[6], a[6], b[1], !b[3]);
	and _ECO_815(w_eco815, a[2], b[2], !a[5], b[7], a[7], !a[3], a[4], b[6], a[6], !a[0], !b[3]);
	and _ECO_816(w_eco816, a[2], b[2], !b[5], !a[5], b[7], !a[3], a[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_817(w_eco817, !b[2], !b[5], a[5], b[7], a[3], a[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_818(w_eco818, !b[5], !b[7], !a[7], a[3], b[4], !b[6], !a[6], b[1], !b[3]);
	and _ECO_819(w_eco819, a[1], !b[2], !b[7], a[3], b[4], !b[6], !a[6], b[1], !b[3], b[0]);
	and _ECO_820(w_eco820, a[2], a[1], b[5], !a[5], b[7], a[3], b[4], a[4], b[6], !a[6]);
	and _ECO_821(w_eco821, a[2], b[2], b[5], a[5], !a[7], a[3], b[4], !b[6], a[6], a[0]);
	and _ECO_822(w_eco822, a[1], !a[5], a[7], !a[3], a[4], !b[6], !a[6], !b[1], b[3]);
	and _ECO_823(w_eco823, a[1], b[5], !a[5], !b[7], !a[3], a[4], b[6], !a[6], !b[1], b[3], b[0]);
	and _ECO_824(w_eco824, !a[1], !b[5], !b[7], !a[7], b[4], !b[6], !a[6], a[0]);
	and _ECO_825(w_eco825, a[2], !a[1], b[2], b[5], a[5], b[7], b[4], !b[6], a[6], a[0]);
	and _ECO_826(w_eco826, b[2], b[5], a[5], b[7], b[6], !a[6], !a[0]);
	and _ECO_827(w_eco827, b[2], !b[5], !a[5], a[7], !a[3], a[4], !b[6], !a[6], !b[1], !a[0]);
	and _ECO_828(w_eco828, b[2], b[5], a[5], !a[7], !a[3], a[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_829(w_eco829, !a[1], b[2], !a[5], !a[7], !a[3], b[4], a[4], !b[6], a[6], !b[3], b[0]);
	and _ECO_830(w_eco830, !a[2], !a[5], b[7], a[7], a[4], b[6], a[6], !b[1], !a[0], b[3]);
	and _ECO_831(w_eco831, !a[2], !b[5], !a[5], a[7], a[4], !b[6], !a[6], !b[1], !a[0], b[3]);
	and _ECO_832(w_eco832, !a[2], b[2], !b[5], !a[5], a[7], !a[3], !b[6], a[6], !b[1], b[3]);
	and _ECO_833(w_eco833, a[1], !a[5], !b[7], !a[3], b[6], !a[6], a[0], b[3]);
	and _ECO_834(w_eco834, b[2], !b[5], b[7], !b[4], a[4], b[6], !a[6], !a[0]);
	and _ECO_835(w_eco835, !a[2], !a[5], b[7], a[7], !a[3], a[4], b[6], a[6], !b[1], !a[0]);
	and _ECO_836(w_eco836, a[2], !b[2], !b[5], a[5], b[7], a[3], a[4], b[6], !a[6], b[0]);
	and _ECO_837(w_eco837, a[2], a[1], !b[2], !a[5], a[7], !b[6], !a[6], b[0]);
	and _ECO_838(w_eco838, a[2], !b[2], !b[5], a[5], b[7], !b[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_839(w_eco839, a[2], a[1], b[5], a[5], b[7], !a[7], !b[4], !a[4], b[6], a[6], b[1]);
	and _ECO_840(w_eco840, a[2], !b[2], !b[5], a[5], b[7], a[3], !b[4], b[6], !a[6], b[0]);
	and _ECO_841(w_eco841, a[2], !b[2], !b[7], !a[7], !a[4], b[6], a[6], b[1]);
	and _ECO_842(w_eco842, a[2], !b[2], !b[5], !b[7], !a[7], !a[4], !b[6], !a[6], b[1]);
	and _ECO_843(w_eco843, a[2], a[1], !b[2], b[5], !a[5], a[7], a[3], !b[4], !b[6], !a[6], b[1]);
	and _ECO_844(w_eco844, !b[5], !b[7], !a[7], b[4], !b[6], !a[6], b[1], a[0]);
	and _ECO_845(w_eco845, a[2], !b[2], !b[5], a[5], b[7], a[4], b[6], !a[6], !b[3], b[0]);
	and _ECO_846(w_eco846, a[2], !b[2], !b[7], !a[7], b[4], b[6], a[6], b[1]);
	and _ECO_847(w_eco847, a[2], !b[2], !b[5], !b[7], !a[7], b[4], !b[6], !a[6], b[1]);
	and _ECO_848(w_eco848, a[2], !b[2], !b[5], a[5], b[7], a[4], b[6], !a[6], !a[0], b[0]);
	and _ECO_849(w_eco849, a[2], !b[2], !b[5], !a[5], !a[7], !a[3], b[4], !b[6], !a[6], b[1], b[3], b[0]);
	and _ECO_850(w_eco850, a[2], !a[1], !b[2], b[5], b[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_851(w_eco851, a[2], !b[2], b[5], !a[5], a[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_852(w_eco852, a[2], !b[2], !a[5], a[7], !b[6], !a[6], !b[1], b[0]);
	and _ECO_853(w_eco853, a[2], !a[1], !b[2], b[5], !a[4], !b[6], !a[6], !b[1], b[0]);
	and _ECO_854(w_eco854, !b[5], !a[5], a[7], !a[3], !b[6], a[6], !b[1], !a[0], b[3]);
	and _ECO_855(w_eco855, a[1], b[5], a[5], b[7], a[3], b[4], a[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_856(w_eco856, !a[2], !b[2], !b[5], !a[5], b[7], a[3], a[4], b[6], a[6], !a[0], b[3]);
	and _ECO_857(w_eco857, !a[2], !b[2], !b[5], !a[5], b[7], a[3], a[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_858(w_eco858, !a[2], !b[2], b[5], a[5], b[7], !a[3], b[4], !b[6], a[6], b[1], a[0]);
	and _ECO_859(w_eco859, a[1], b[5], a[5], b[7], !a[3], b[4], a[4], !b[6], !a[6], b[1], !b[3]);
	and _ECO_860(w_eco860, !a[2], !b[2], !a[5], b[7], a[7], !a[3], a[4], b[6], a[6], !a[0], !b[3]);
	and _ECO_861(w_eco861, !a[2], !b[2], !b[5], !a[5], b[7], !a[3], a[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_862(w_eco862, !b[2], !b[5], !a[5], !a[7], !b[6], a[6], a[0]);
	and _ECO_863(w_eco863, a[1], !b[7], !a[3], b[6], !a[6], a[0], b[3], !b[0]);
	and _ECO_864(w_eco864, b[5], !a[5], b[7], !a[3], !b[4], a[4], b[6], a[6], b[3], !b[0]);
	and _ECO_865(w_eco865, a[1], b[5], !a[5], !a[3], a[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_866(w_eco866, !b[5], b[7], !b[4], a[4], b[6], !a[6], !a[0], !b[0]);
	and _ECO_867(w_eco867, !b[7], !a[3], b[6], !a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_868(w_eco868, !a[2], a[1], !b[5], b[7], a[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_869(w_eco869, !a[2], !a[1], !b[2], b[5], a[5], b[7], !a[3], b[4], !b[6], a[6], a[0]);
	and _ECO_870(w_eco870, !a[1], !b[7], !a[7], b[4], b[6], a[6], a[0]);
	and _ECO_871(w_eco871, !a[2], b[5], a[5], b[7], b[6], !a[6], !a[0]);
	and _ECO_872(w_eco872, !a[2], b[5], a[5], !a[7], !a[3], a[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_873(w_eco873, a[1], b[5], !a[5], !b[7], !a[3], !b[6], b[3], !b[0]);
	and _ECO_874(w_eco874, a[2], a[1], b[2], a[5], !b[7], !a[3], b[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_875(w_eco875, a[2], !b[5], !a[5], !a[7], a[4], !b[6], a[6], !b[3]);
	and _ECO_876(w_eco876, a[2], !a[1], a[5], !b[7], !a[7], !a[3], b[4], a[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_877(w_eco877, a[2], a[1], b[5], a[5], b[7], b[4], !b[6], a[6], a[0], !b[0]);
	and _ECO_878(w_eco878, a[1], b[5], !a[5], !a[3], a[4], b[6], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_879(w_eco879, a[1], !b[7], !a[7], !a[3], b[4], !b[6], a[6], a[0], b[3], !b[0]);
	and _ECO_880(w_eco880, !a[1], b[2], b[5], b[7], b[4], b[6], !a[6], !a[0], b[3]);
	and _ECO_881(w_eco881, !a[1], b[5], !a[5], !b[7], !a[7], b[6], a[6], !b[0]);
	and _ECO_882(w_eco882, b[5], !a[5], !b[7], !a[3], !b[6], !b[1], b[3], !b[0]);
	and _ECO_883(w_eco883, !a[1], b[2], b[5], b[7], !a[3], b[4], b[6], !a[6], !a[0]);
	and _ECO_884(w_eco884, !a[2], !b[5], !a[5], b[7], !a[7], a[3], b[4], a[4], b[6], a[0]);
	and _ECO_885(w_eco885, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], b[4], b[6], !a[0]);
	and _ECO_886(w_eco886, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], b[4], a[4], !a[6]);
	and _ECO_887(w_eco887, a[1], !b[5], !a[5], !a[7], !a[3], !b[6], a[6], a[0], b[3], !b[0]);
	and _ECO_888(w_eco888, !a[2], a[1], b[2], !b[5], !a[5], b[7], a[4], !b[6], !a[6], !b[1], !b[0]);
	and _ECO_889(w_eco889, !a[2], b[2], !b[7], !a[7], !a[3], b[6], a[6], b[3], !b[0]);
	and _ECO_890(w_eco890, !a[2], !b[5], !a[5], b[7], !a[7], a[3], b[4], b[6], !a[0], !b[3]);
	and _ECO_891(w_eco891, !a[2], !b[5], !a[5], b[7], !a[7], a[3], b[4], a[4], !a[6], !b[3]);
	and _ECO_892(w_eco892, !a[2], !b[5], !a[5], b[7], !a[7], b[4], a[4], b[6], a[0], !b[3]);
	and _ECO_893(w_eco893, a[2], !a[1], !b[2], b[5], !a[5], !b[7], !b[6], !b[1], !b[0]);
	and _ECO_894(w_eco894, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[3], a[4], b[6], !a[6]);
	and _ECO_895(w_eco895, b[5], a[5], b[7], b[6], !a[6], !a[0], !b[0]);
	and _ECO_896(w_eco896, a[2], !a[1], !b[2], b[5], !a[5], !b[7], !b[4], b[6], !a[6], !b[3]);
	and _ECO_897(w_eco897, b[5], a[5], b[7], !b[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_898(w_eco898, a[2], b[5], a[5], b[7], !a[3], b[4], !b[6], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_899(w_eco899, b[5], a[5], b[7], a[4], b[6], !a[6], !b[3], !b[0]);
	and _ECO_900(w_eco900, a[2], !b[5], !a[5], b[7], !a[7], a[4], !b[3], !b[0]);
	and _ECO_901(w_eco901, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[4], b[6], !a[6], !b[3]);
	and _ECO_902(w_eco902, !a[2], !b[2], b[5], a[5], !a[7], b[4], a[6], b[1], a[0], b[3]);
	and _ECO_903(w_eco903, a[1], b[5], !a[5], b[7], a[3], a[4], !b[6], !a[6], b[1], !b[3], !b[0]);
	and _ECO_904(w_eco904, !a[2], !a[1], b[5], b[7], b[4], b[6], !a[6], !a[0], b[3]);
	and _ECO_905(w_eco905, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], b[4], !b[6], a[6], b[1]);
	and _ECO_906(w_eco906, a[1], !b[2], b[5], a[5], b[7], b[4], !b[6], a[6], a[0], !b[0]);
	and _ECO_907(w_eco907, !a[2], !a[1], b[5], a[5], b[7], !a[7], !a[3], b[4], b[6], !a[0]);
	and _ECO_908(w_eco908, !a[2], !a[1], b[5], !a[5], b[7], !a[3], a[4], !b[6], !a[6], !a[0], b[3], !b[0]);
	and _ECO_909(w_eco909, !a[2], !a[1], b[5], b[7], !a[3], b[4], b[6], !a[6], !a[0]);
	and _ECO_910(w_eco910, a[2], a[1], !b[2], !a[5], !a[3], b[6], !a[6], a[0], b[3], b[0]);
	and _ECO_911(w_eco911, !a[2], !b[5], b[7], !b[4], a[4], b[6], !a[6], !a[0]);
	and _ECO_912(w_eco912, !a[5], b[7], !a[3], !b[4], a[4], b[6], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_913(w_eco913, !a[2], b[2], !a[5], !a[3], !b[4], a[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_914(w_eco914, a[2], b[2], !b[5], !a[5], b[7], a[3], !b[4], b[6], a[6], !a[0], b[3]);
	and _ECO_915(w_eco915, a[2], b[2], !b[5], !a[5], b[7], a[3], !b[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_916(w_eco916, a[2], !b[5], !a[5], !a[7], a[3], !b[4], !b[6], a[6]);
	and _ECO_917(w_eco917, a[2], !a[1], !b[2], b[5], !a[5], !b[7], a[3], !b[4], b[6], !a[6]);
	and _ECO_918(w_eco918, a[2], b[2], b[5], a[5], b[7], !a[4], !b[6], a[6], b[1], a[0]);
	and _ECO_919(w_eco919, a[2], b[2], !a[5], b[7], a[7], !a[3], !b[4], b[6], a[6], !a[0], !b[3]);
	and _ECO_920(w_eco920, a[2], b[2], !b[5], !a[5], b[7], !a[3], !b[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_921(w_eco921, a[2], !b[5], !a[5], !a[7], !b[4], !b[6], a[6], !b[3]);
	and _ECO_922(w_eco922, a[1], !a[5], a[7], !a[3], !b[4], !b[6], !a[6], !b[1], b[3]);
	and _ECO_923(w_eco923, a[1], b[5], !a[5], !b[7], !a[3], !b[4], b[6], !a[6], !b[1], b[3], b[0]);
	and _ECO_924(w_eco924, a[2], b[2], b[5], a[5], b[7], !a[4], !b[6], a[6], a[0], !b[3]);
	and _ECO_925(w_eco925, a[2], a[1], b[5], !a[5], b[7], !b[4], !a[4], b[6], !a[6], !b[3]);
	and _ECO_926(w_eco926, a[2], b[2], b[5], a[5], !a[7], !a[4], !b[6], a[6], a[0], !b[3]);
	and _ECO_927(w_eco927, a[2], b[2], b[5], b[7], !b[4], !a[4], !b[6], a[6], !b[3]);
	and _ECO_928(w_eco928, a[2], !a[1], b[2], b[5], a[5], b[7], !a[4], !b[6], a[6], a[0]);
	and _ECO_929(w_eco929, b[2], !b[5], !a[5], a[7], !a[3], !b[4], !b[6], !a[6], !b[1], !a[0]);
	and _ECO_930(w_eco930, b[2], b[5], a[5], !a[7], !a[3], !b[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_931(w_eco931, !a[1], !b[5], !b[7], !a[7], !a[4], !b[6], !a[6], a[0]);
	and _ECO_932(w_eco932, !a[2], !a[5], b[7], a[7], !b[4], b[6], a[6], !b[1], !a[0], b[3]);
	and _ECO_933(w_eco933, !a[2], !b[5], !a[5], a[7], !b[4], !b[6], !a[6], !b[1], !a[0], b[3]);
	and _ECO_934(w_eco934, !b[5], !a[5], !a[7], a[3], !b[4], !b[6], a[6], b[0]);
	and _ECO_935(w_eco935, !a[2], !b[5], !b[7], !a[4], b[6], !a[6], b[1], b[3]);
	and _ECO_936(w_eco936, !a[2], b[5], a[5], b[7], a[3], !b[4], b[6], !a[6]);
	and _ECO_937(w_eco937, !a[2], !a[1], !b[7], a[3], !a[4], !b[6], !a[6], !b[1], !b[3], b[0]);
	and _ECO_938(w_eco938, !a[1], !b[7], !a[7], a[3], !a[4], b[6], a[6], !b[3]);
	and _ECO_939(w_eco939, !a[2], !a[5], b[7], a[7], !a[3], !b[4], b[6], a[6], !b[1], !a[0]);
	and _ECO_940(w_eco940, !b[5], !a[5], !a[7], !b[4], !b[6], a[6], !b[3], b[0]);
	and _ECO_941(w_eco941, a[2], !b[2], !b[5], a[5], b[7], !b[4], b[6], !a[6], !a[0], b[0]);
	and _ECO_942(w_eco942, a[2], !b[2], b[5], !a[5], !b[4], b[6], !a[6], !b[1], b[0]);
	and _ECO_943(w_eco943, a[2], !b[2], !b[5], !a[5], !a[7], !a[3], !a[4], !b[6], !a[6], b[1], b[3], b[0]);
	and _ECO_944(w_eco944, !a[2], !b[2], !b[5], !a[5], b[7], a[3], !b[4], b[6], a[6], !a[0], b[3]);
	and _ECO_945(w_eco945, !a[2], !b[2], !b[5], !a[5], b[7], a[3], !b[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_946(w_eco946, !a[2], !b[2], b[5], a[5], b[7], !a[3], !a[4], !b[6], a[6], b[1], a[0]);
	and _ECO_947(w_eco947, a[1], !b[2], !b[7], a[3], !a[4], !b[6], !a[6], b[1], !b[3], b[0]);
	and _ECO_948(w_eco948, !b[7], !a[7], a[3], !a[4], b[6], a[6], b[1], !b[3]);
	and _ECO_949(w_eco949, a[1], b[5], a[5], b[7], !a[3], !b[4], !a[4], !b[6], !a[6], b[1], !b[3]);
	and _ECO_950(w_eco950, !a[2], !b[2], !a[5], b[7], a[7], !a[3], !b[4], b[6], a[6], !a[0], !b[3]);
	and _ECO_951(w_eco951, !a[2], !b[2], !b[5], !a[5], b[7], !a[3], !b[4], !b[6], !a[6], !a[0], !b[3]);
	and _ECO_952(w_eco952, !a[2], !a[1], b[5], b[7], !a[3], !a[4], b[6], !a[6], b[1]);
	and _ECO_953(w_eco953, !b[5], !b[7], !a[7], !a[3], !a[4], !b[6], !a[6], b[1], b[3]);
	and _ECO_954(w_eco954, !b[2], b[5], !a[5], !b[7], a[7], a[3], !b[4], !b[6], !b[3]);
	and _ECO_955(w_eco955, !a[1], !b[2], !b[7], !a[7], a[3], !b[4], !a[4], !b[6], !a[6], !b[3]);
	and _ECO_956(w_eco956, !a[2], !a[1], !b[2], b[5], a[5], b[7], !a[3], !a[4], !b[6], a[6], a[0]);
	and _ECO_957(w_eco957, !a[2], b[5], a[5], !a[7], !a[3], !b[4], b[6], !a[6], !b[1], !a[0], b[0]);
	and _ECO_958(w_eco958, a[2], a[1], b[2], a[5], !b[7], a[3], !a[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_959(w_eco959, !a[1], b[2], b[5], a[5], b[7], !a[7], !a[4], b[6], !a[0], b[3]);
	and _ECO_960(w_eco960, a[2], !a[1], a[5], !b[7], !a[7], a[3], !b[4], !a[4], !b[6], !a[6], !a[0], b[3]);
	and _ECO_961(w_eco961, !a[1], b[2], b[5], !a[5], !a[7], b[6], a[6], b[1], a[0], !b[0]);
	and _ECO_962(w_eco962, a[2], a[1], b[5], a[5], b[7], !a[4], !b[6], a[6], a[0], !b[0]);
	and _ECO_963(w_eco963, a[1], b[5], !a[5], !a[3], !b[4], b[6], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_964(w_eco964, !a[2], a[1], b[2], !a[5], !a[3], !b[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_965(w_eco965, a[1], b[5], !a[5], !a[3], !b[4], !b[6], !a[6], !b[1], b[3], !b[0]);
	and _ECO_966(w_eco966, a[1], !b[7], !a[7], !a[3], !a[4], !b[6], a[6], a[0], b[3], !b[0]);
	and _ECO_967(w_eco967, !a[1], b[2], b[5], b[7], !a[4], b[6], !a[6], !a[0], b[3]);
	and _ECO_968(w_eco968, !a[1], b[2], b[5], b[7], !a[3], !a[4], b[6], !a[6], !a[0]);
	and _ECO_969(w_eco969, !a[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !a[4], b[6], a[0]);
	and _ECO_970(w_eco970, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], !a[4], b[6], !a[0]);
	and _ECO_971(w_eco971, !a[2], a[1], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !a[4], !a[6]);
	and _ECO_972(w_eco972, !a[2], !b[5], !a[5], b[7], !a[7], a[3], !a[4], b[6], !a[0], !b[3]);
	and _ECO_973(w_eco973, !a[2], !b[5], !a[5], b[7], !a[7], a[3], !b[4], !a[4], !a[6], !b[3]);
	and _ECO_974(w_eco974, a[2], b[5], a[5], b[7], !a[3], !a[4], !b[6], a[6], !b[1], a[0], b[3], !b[0]);
	and _ECO_975(w_eco975, !a[2], !b[2], b[5], a[5], !a[7], !a[4], a[6], b[1], a[0], b[3]);
	and _ECO_976(w_eco976, !b[2], !b[5], !a[5], !a[7], a[3], !b[4], !b[6], a[6]);
	and _ECO_977(w_eco977, a[1], b[5], !a[5], b[7], a[3], !b[4], !b[6], !a[6], b[1], a[0], !b[0]);
	and _ECO_978(w_eco978, a[1], b[5], !a[5], b[7], a[3], !b[4], !b[6], !a[6], b[1], !b[3], !b[0]);
	and _ECO_979(w_eco979, a[1], b[5], !a[5], !a[7], a[3], b[6], a[6], b[1], !a[0], !b[3], !b[0]);
	and _ECO_980(w_eco980, !b[5], !b[7], !a[7], a[3], !a[4], !b[6], !a[6], b[1], !b[3]);
	and _ECO_981(w_eco981, !a[2], !a[1], b[5], b[7], !a[4], b[6], !a[6], !a[0], b[3]);
	and _ECO_982(w_eco982, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[3], !a[4], !b[6], a[6], b[1]);
	and _ECO_983(w_eco983, a[1], !b[2], b[5], a[5], b[7], !a[4], !b[6], a[6], a[0], !b[0]);
	and _ECO_984(w_eco984, !a[2], !a[1], !b[2], b[5], a[5], !a[7], !a[4], a[6], a[0], b[3]);
	and _ECO_985(w_eco985, !a[2], !a[1], b[5], a[5], b[7], !a[7], !a[3], !a[4], b[6], !a[0]);
	and _ECO_986(w_eco986, !a[2], !a[1], b[5], !a[5], b[7], !a[3], !b[4], !b[6], !a[6], !a[0], b[3], !b[0]);
	and _ECO_987(w_eco987, !a[2], !a[1], b[5], b[7], !a[3], !a[4], b[6], !a[6], !a[0]);
	or _ECO_988(w_eco988, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987);
	xor _ECO_out0(a_gtet_b, sub_wire0, w_eco988);

endmodule