module top(Sync,Gate,Done,cnt,clk,ena,rst,Tsync,Tgdel,Tgate,Tlen,prev_state,prev_cnt,prev_cnt_len);
	input clk, ena, rst;
	input [7:0]Tsync, Tgdel;
	input [15:0]Tgate, Tlen;
	input [4:0]prev_state;
	input [15:0]prev_cnt, prev_cnt_len;
	output Sync, Gate, Done;
	output [15:0]cnt;
	wire \mux_cnt_122_11_g657/w_0, \mux_cnt_122_11_g657/w_1, \mux_cnt_122_11_g657/w_2, \mux_cnt_122_11_g657/w_3, \mux_cnt_122_11_g657/w_4, \mux_cnt_122_11_g661/w_0, \mux_cnt_122_11_g661/w_1, \mux_cnt_122_11_g661/w_2, \mux_cnt_122_11_g661/w_3, \mux_cnt_122_11_g661/w_4, \mux_cnt_122_11_g665/w_0, \mux_cnt_122_11_g665/w_1, \mux_cnt_122_11_g665/w_2, \mux_cnt_122_11_g665/w_3, \mux_cnt_122_11_g665/w_4, \mux_cnt_122_11_g669/w_0, \mux_cnt_122_11_g669/w_1, \mux_cnt_122_11_g669/w_2, \mux_cnt_122_11_g669/w_3, \mux_cnt_122_11_g669/w_4, \mux_cnt_122_11_g673/w_0, \mux_cnt_122_11_g673/w_1, \mux_cnt_122_11_g673/w_2, \mux_cnt_122_11_g673/w_3, \mux_cnt_122_11_g673/w_4, \mux_cnt_122_11_g677/w_0, \mux_cnt_122_11_g677/w_1, \mux_cnt_122_11_g677/w_2, \mux_cnt_122_11_g677/w_3, \mux_cnt_122_11_g677/w_4, \mux_cnt_122_11_g681/w_0, \mux_cnt_122_11_g681/w_1, \mux_cnt_122_11_g681/w_2, \mux_cnt_122_11_g681/w_3, \mux_cnt_122_11_g681/w_4, \mux_cnt_122_11_g713/w_0, \mux_cnt_122_11_g713/w_1, \mux_cnt_122_11_g713/w_2, \mux_cnt_122_11_g713/w_3, \mux_cnt_122_11_g713/w_4, \mux_cnt_122_11_g653/w_0, \mux_cnt_122_11_g653/w_1, \mux_cnt_122_11_g653/w_2, \mux_cnt_122_11_g685/w_0, \mux_cnt_122_11_g685/w_1, \mux_cnt_122_11_g685/w_2, \mux_cnt_122_11_g689/w_0, \mux_cnt_122_11_g689/w_1, \mux_cnt_122_11_g689/w_2, \mux_cnt_122_11_g693/w_0, \mux_cnt_122_11_g693/w_1, \mux_cnt_122_11_g693/w_2, \mux_cnt_122_11_g697/w_0, \mux_cnt_122_11_g697/w_1, \mux_cnt_122_11_g697/w_2, \mux_cnt_122_11_g701/w_0, \mux_cnt_122_11_g701/w_1, \mux_cnt_122_11_g701/w_2, \mux_cnt_122_11_g705/w_0, \mux_cnt_122_11_g705/w_1, \mux_cnt_122_11_g705/w_2, \mux_cnt_122_11_g709/w_0, \mux_cnt_122_11_g709/w_1, \mux_cnt_122_11_g709/w_2, sub_111_47_n_67, sub_108_39_n_949, sub_108_39_n_166, sub_108_39_n_159, sub_108_39_n_151, sub_108_39_n_139, sub_108_39_n_119, sub_108_39_n_109, sub_108_39_n_103, sub_108_39_n_67, n_1387, n_1382, n_1257, n_1256, n_1255, n_1254, n_1253, n_1252, n_1251, n_1250, n_1249, n_1248, n_1247, n_1246, n_1245, n_1244, n_1243, n_1242, n_1241, n_1240, n_1239, n_1238, n_1237, n_1236, n_1235, n_1234, n_1233, n_1232, n_1231, n_1230, n_1229, n_1228, n_1227, n_1226, n_1225, n_1224, n_1223, n_1222, n_1220, n_1218, n_1217, n_1216, n_1215, n_1214, n_1213, n_1212, n_1211, n_1210, n_1209, n_1208, n_1207, n_1206, n_1205, n_1204, n_1203, n_1202, n_1201, n_1200, n_1199, n_1198, n_1197, n_1196, n_1195, n_1194, n_1193, n_1192, n_1191, n_1190, n_1189, n_1188, n_1187, n_1186, n_1185, n_1184, n_1183, n_1164, n_1162, n_1161, n_1160, n_1078, n_1069, n_1062, n_1052, n_1049, n_1043, n_995, n_977, n_976, n_975, n_941, n_746, n_744, n_741, n_732, n_326, n_45, n_44, n_43, Done, Gate, Sync, rst, ena, clk, \mux_cnt_122_11_g657/data0, \mux_cnt_122_11_g661/data0, \mux_cnt_122_11_g665/data0, \mux_cnt_122_11_g669/data0, \mux_cnt_122_11_g673/data0, \mux_cnt_122_11_g677/data0, \mux_cnt_122_11_g681/data0, \mux_cnt_122_11_g713/data0, \mux_cnt_122_11_g653/data0, \mux_cnt_122_11_g685/data0, \mux_cnt_122_11_g689/data0, \mux_cnt_122_11_g693/data0, \mux_cnt_122_11_g697/data0, \mux_cnt_122_11_g701/data0, \mux_cnt_122_11_g705/data0, \mux_cnt_122_11_g709/data0;
	wire [16:0]cnt_nxt;
	wire [15:0]cnt;
	wire [4:0]prev_state;
	wire [15:0]prev_cnt_len, prev_cnt, Tlen, Tgate;
	wire [7:0]Tgdel, Tsync;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, sub_wire1, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634, w_eco1635, sub_wire2, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, sub_wire3, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914, w_eco1915, w_eco1916, w_eco1917, w_eco1918, w_eco1919, w_eco1920, w_eco1921, w_eco1922, w_eco1923, w_eco1924, w_eco1925, w_eco1926, w_eco1927, w_eco1928, w_eco1929, w_eco1930, w_eco1931, w_eco1932, w_eco1933, w_eco1934, w_eco1935, w_eco1936, w_eco1937, w_eco1938, w_eco1939, w_eco1940, w_eco1941, w_eco1942, w_eco1943, w_eco1944, w_eco1945, w_eco1946, w_eco1947, w_eco1948, w_eco1949, w_eco1950, w_eco1951, w_eco1952, w_eco1953, w_eco1954, w_eco1955, w_eco1956, w_eco1957, w_eco1958, w_eco1959, w_eco1960, w_eco1961, w_eco1962, w_eco1963, w_eco1964, w_eco1965, w_eco1966, w_eco1967, w_eco1968, w_eco1969, w_eco1970, w_eco1971, w_eco1972, w_eco1973, w_eco1974, w_eco1975, w_eco1976, w_eco1977, w_eco1978, w_eco1979, w_eco1980, w_eco1981, w_eco1982, w_eco1983, w_eco1984, w_eco1985, w_eco1986, w_eco1987, w_eco1988, w_eco1989, w_eco1990, w_eco1991, w_eco1992, w_eco1993, w_eco1994, w_eco1995, w_eco1996, w_eco1997, w_eco1998, w_eco1999, w_eco2000, w_eco2001, w_eco2002, w_eco2003, w_eco2004, w_eco2005, w_eco2006, w_eco2007, w_eco2008, w_eco2009, w_eco2010, w_eco2011, w_eco2012, w_eco2013, w_eco2014, w_eco2015, w_eco2016, w_eco2017, w_eco2018, w_eco2019, w_eco2020, w_eco2021, w_eco2022, w_eco2023, w_eco2024, w_eco2025, w_eco2026, w_eco2027, w_eco2028, w_eco2029, w_eco2030, w_eco2031, w_eco2032, w_eco2033, w_eco2034, w_eco2035, w_eco2036, w_eco2037, w_eco2038, w_eco2039, w_eco2040, w_eco2041, w_eco2042, w_eco2043, w_eco2044, w_eco2045, w_eco2046, w_eco2047, w_eco2048, w_eco2049, w_eco2050, w_eco2051, w_eco2052, w_eco2053, w_eco2054, w_eco2055, w_eco2056, w_eco2057, w_eco2058, w_eco2059, w_eco2060, w_eco2061, w_eco2062, w_eco2063, w_eco2064, w_eco2065, w_eco2066, w_eco2067, w_eco2068, w_eco2069, w_eco2070, w_eco2071, w_eco2072, w_eco2073, w_eco2074, w_eco2075, w_eco2076, w_eco2077, w_eco2078, w_eco2079, w_eco2080, w_eco2081, w_eco2082, w_eco2083, w_eco2084, w_eco2085, w_eco2086, w_eco2087, w_eco2088, w_eco2089, w_eco2090, w_eco2091, w_eco2092, w_eco2093, w_eco2094, w_eco2095, w_eco2096, w_eco2097, w_eco2098, w_eco2099, w_eco2100, w_eco2101, w_eco2102, w_eco2103, w_eco2104, w_eco2105, w_eco2106, w_eco2107, w_eco2108, w_eco2109, w_eco2110, w_eco2111, w_eco2112, w_eco2113, w_eco2114, w_eco2115, w_eco2116, w_eco2117, w_eco2118, w_eco2119, w_eco2120, w_eco2121, w_eco2122, w_eco2123, w_eco2124, w_eco2125, w_eco2126, w_eco2127, w_eco2128, w_eco2129, w_eco2130, w_eco2131, w_eco2132, w_eco2133, w_eco2134, w_eco2135, w_eco2136, w_eco2137, w_eco2138, w_eco2139, w_eco2140, w_eco2141, w_eco2142, w_eco2143, w_eco2144, w_eco2145, w_eco2146, w_eco2147, w_eco2148, w_eco2149, w_eco2150, w_eco2151, w_eco2152, w_eco2153, w_eco2154, w_eco2155, w_eco2156, w_eco2157, w_eco2158, w_eco2159, w_eco2160, w_eco2161, w_eco2162, w_eco2163, w_eco2164, w_eco2165, w_eco2166, w_eco2167, w_eco2168, w_eco2169, w_eco2170, w_eco2171, w_eco2172, w_eco2173, w_eco2174, w_eco2175, w_eco2176, w_eco2177, w_eco2178, w_eco2179, w_eco2180, w_eco2181, w_eco2182, w_eco2183, w_eco2184, w_eco2185, w_eco2186, w_eco2187, w_eco2188, w_eco2189, w_eco2190, w_eco2191, w_eco2192, w_eco2193, w_eco2194, w_eco2195, w_eco2196, w_eco2197, w_eco2198, w_eco2199, w_eco2200, w_eco2201, w_eco2202, w_eco2203, w_eco2204, w_eco2205, w_eco2206, w_eco2207, w_eco2208, w_eco2209, w_eco2210, w_eco2211, w_eco2212, w_eco2213, w_eco2214, w_eco2215, w_eco2216, w_eco2217, w_eco2218, w_eco2219, w_eco2220, w_eco2221, w_eco2222, w_eco2223, w_eco2224, w_eco2225, w_eco2226, w_eco2227, w_eco2228, w_eco2229, w_eco2230, w_eco2231, w_eco2232, w_eco2233, w_eco2234, w_eco2235, w_eco2236, w_eco2237, w_eco2238, w_eco2239, w_eco2240, w_eco2241, w_eco2242, w_eco2243, w_eco2244, w_eco2245, w_eco2246, w_eco2247, w_eco2248, w_eco2249, w_eco2250, w_eco2251, w_eco2252, w_eco2253, w_eco2254, w_eco2255, w_eco2256, w_eco2257, w_eco2258, w_eco2259, w_eco2260, w_eco2261, w_eco2262, w_eco2263, w_eco2264, w_eco2265, w_eco2266, w_eco2267, w_eco2268, w_eco2269, w_eco2270, w_eco2271, w_eco2272, w_eco2273, w_eco2274, w_eco2275, w_eco2276, w_eco2277, w_eco2278, w_eco2279, w_eco2280, w_eco2281, w_eco2282, w_eco2283, w_eco2284, w_eco2285, w_eco2286, w_eco2287, w_eco2288, w_eco2289, w_eco2290, w_eco2291, w_eco2292, w_eco2293, w_eco2294, w_eco2295, w_eco2296, w_eco2297, w_eco2298, w_eco2299, w_eco2300, w_eco2301, w_eco2302, w_eco2303, w_eco2304, w_eco2305, w_eco2306, w_eco2307, w_eco2308, w_eco2309, w_eco2310, w_eco2311, w_eco2312, w_eco2313, w_eco2314, w_eco2315, w_eco2316, w_eco2317, w_eco2318, w_eco2319, w_eco2320, w_eco2321, w_eco2322, w_eco2323, w_eco2324, w_eco2325, w_eco2326, w_eco2327, w_eco2328, w_eco2329, w_eco2330, w_eco2331, w_eco2332, w_eco2333, w_eco2334, w_eco2335, w_eco2336, w_eco2337, w_eco2338, w_eco2339, w_eco2340, w_eco2341, w_eco2342, w_eco2343, w_eco2344, w_eco2345, w_eco2346, w_eco2347, w_eco2348, w_eco2349, w_eco2350, w_eco2351, w_eco2352, w_eco2353, w_eco2354, w_eco2355, w_eco2356, w_eco2357, w_eco2358, w_eco2359, w_eco2360, w_eco2361, w_eco2362, w_eco2363, w_eco2364, w_eco2365, w_eco2366, w_eco2367, w_eco2368, w_eco2369, w_eco2370, w_eco2371, w_eco2372, w_eco2373, w_eco2374, w_eco2375, w_eco2376, w_eco2377, w_eco2378, w_eco2379, w_eco2380, w_eco2381, w_eco2382, w_eco2383, w_eco2384, w_eco2385, w_eco2386, w_eco2387, w_eco2388, w_eco2389, w_eco2390, w_eco2391, w_eco2392, w_eco2393, w_eco2394, w_eco2395, w_eco2396, w_eco2397, w_eco2398, w_eco2399, w_eco2400, w_eco2401, w_eco2402, w_eco2403, w_eco2404, w_eco2405, w_eco2406, w_eco2407, w_eco2408, w_eco2409, w_eco2410, w_eco2411, w_eco2412, w_eco2413, w_eco2414, w_eco2415, w_eco2416, w_eco2417, w_eco2418, w_eco2419, w_eco2420, w_eco2421, w_eco2422, w_eco2423, w_eco2424, w_eco2425, w_eco2426, w_eco2427, w_eco2428, w_eco2429, w_eco2430, w_eco2431, w_eco2432, w_eco2433, w_eco2434, w_eco2435, w_eco2436, w_eco2437, w_eco2438, w_eco2439, w_eco2440, w_eco2441, w_eco2442, w_eco2443, w_eco2444, w_eco2445, w_eco2446, w_eco2447, w_eco2448, w_eco2449, w_eco2450, w_eco2451, w_eco2452, w_eco2453, w_eco2454, w_eco2455, w_eco2456, w_eco2457, w_eco2458, w_eco2459, w_eco2460, w_eco2461, w_eco2462, w_eco2463, w_eco2464, w_eco2465, w_eco2466, w_eco2467, w_eco2468, w_eco2469, w_eco2470, w_eco2471, w_eco2472, w_eco2473, w_eco2474, w_eco2475, w_eco2476, w_eco2477, w_eco2478, w_eco2479, w_eco2480, w_eco2481, w_eco2482, w_eco2483, w_eco2484, w_eco2485, w_eco2486, w_eco2487, w_eco2488, w_eco2489, w_eco2490, w_eco2491, w_eco2492, w_eco2493, w_eco2494, w_eco2495, w_eco2496, w_eco2497, w_eco2498, w_eco2499, w_eco2500, w_eco2501, w_eco2502, w_eco2503, w_eco2504, w_eco2505, w_eco2506, w_eco2507, w_eco2508, w_eco2509, w_eco2510, w_eco2511, w_eco2512, w_eco2513, w_eco2514, w_eco2515, w_eco2516, w_eco2517, w_eco2518, w_eco2519, w_eco2520, w_eco2521, w_eco2522, w_eco2523, w_eco2524, w_eco2525, w_eco2526, w_eco2527, w_eco2528, w_eco2529, w_eco2530, w_eco2531, w_eco2532, w_eco2533, w_eco2534, w_eco2535, w_eco2536, w_eco2537, w_eco2538, w_eco2539, w_eco2540, w_eco2541, w_eco2542, w_eco2543, w_eco2544, w_eco2545, w_eco2546, w_eco2547, w_eco2548, w_eco2549, w_eco2550, w_eco2551, w_eco2552, w_eco2553, w_eco2554, w_eco2555, w_eco2556, w_eco2557, w_eco2558, w_eco2559, w_eco2560, w_eco2561, w_eco2562, w_eco2563, w_eco2564, w_eco2565, w_eco2566, w_eco2567, w_eco2568, w_eco2569, w_eco2570, w_eco2571, w_eco2572, w_eco2573, w_eco2574, w_eco2575, w_eco2576, w_eco2577, w_eco2578, w_eco2579, w_eco2580, w_eco2581, w_eco2582, w_eco2583, w_eco2584, w_eco2585, w_eco2586, w_eco2587, w_eco2588, w_eco2589, w_eco2590, w_eco2591, w_eco2592, w_eco2593, w_eco2594, w_eco2595, w_eco2596, w_eco2597, w_eco2598, w_eco2599, w_eco2600, w_eco2601, w_eco2602, w_eco2603, w_eco2604, w_eco2605, w_eco2606, w_eco2607, w_eco2608, w_eco2609, w_eco2610, w_eco2611, w_eco2612, w_eco2613, w_eco2614, w_eco2615, w_eco2616, w_eco2617, w_eco2618, w_eco2619, w_eco2620, w_eco2621, w_eco2622, w_eco2623, w_eco2624, w_eco2625, w_eco2626, w_eco2627, w_eco2628, w_eco2629, w_eco2630, w_eco2631, w_eco2632, w_eco2633, w_eco2634, w_eco2635, w_eco2636, w_eco2637, w_eco2638, w_eco2639, w_eco2640, w_eco2641, w_eco2642, w_eco2643, w_eco2644, w_eco2645, w_eco2646, w_eco2647, w_eco2648, w_eco2649, w_eco2650, w_eco2651, w_eco2652, w_eco2653, w_eco2654, w_eco2655, w_eco2656, w_eco2657, w_eco2658, w_eco2659, w_eco2660, w_eco2661, w_eco2662, w_eco2663, w_eco2664, w_eco2665, w_eco2666, w_eco2667, w_eco2668, w_eco2669, w_eco2670, w_eco2671, w_eco2672, w_eco2673, w_eco2674, w_eco2675, w_eco2676, w_eco2677, w_eco2678, w_eco2679, w_eco2680, w_eco2681, w_eco2682, w_eco2683, w_eco2684, w_eco2685, w_eco2686, w_eco2687, w_eco2688, w_eco2689, w_eco2690, w_eco2691, w_eco2692, w_eco2693, w_eco2694, w_eco2695, w_eco2696, w_eco2697, w_eco2698, w_eco2699, w_eco2700, w_eco2701, w_eco2702, w_eco2703, w_eco2704, w_eco2705, w_eco2706, w_eco2707, w_eco2708, w_eco2709, w_eco2710, w_eco2711, w_eco2712, w_eco2713, w_eco2714, w_eco2715, w_eco2716, w_eco2717, w_eco2718, w_eco2719, w_eco2720, w_eco2721, w_eco2722, w_eco2723, w_eco2724, w_eco2725, w_eco2726, w_eco2727, w_eco2728, w_eco2729, w_eco2730, w_eco2731, w_eco2732, w_eco2733, w_eco2734, w_eco2735, w_eco2736, w_eco2737, w_eco2738, w_eco2739, w_eco2740, w_eco2741, w_eco2742, w_eco2743, w_eco2744, w_eco2745, w_eco2746, w_eco2747, w_eco2748, w_eco2749, w_eco2750, w_eco2751, w_eco2752, w_eco2753, w_eco2754, w_eco2755, w_eco2756, w_eco2757, w_eco2758, w_eco2759, w_eco2760, w_eco2761, w_eco2762, w_eco2763, w_eco2764, w_eco2765, w_eco2766, w_eco2767, w_eco2768, w_eco2769, w_eco2770, w_eco2771, w_eco2772, w_eco2773, w_eco2774, w_eco2775, w_eco2776, w_eco2777, w_eco2778, w_eco2779, w_eco2780, w_eco2781, w_eco2782, w_eco2783, w_eco2784, w_eco2785, w_eco2786, w_eco2787, w_eco2788, w_eco2789, w_eco2790, w_eco2791, w_eco2792, w_eco2793, w_eco2794, w_eco2795, w_eco2796, w_eco2797, w_eco2798, w_eco2799, w_eco2800, w_eco2801, w_eco2802, w_eco2803, w_eco2804, w_eco2805, w_eco2806, w_eco2807, w_eco2808, w_eco2809, w_eco2810, w_eco2811, w_eco2812, w_eco2813, w_eco2814, w_eco2815, w_eco2816, w_eco2817, w_eco2818, w_eco2819, w_eco2820, w_eco2821, w_eco2822, w_eco2823, w_eco2824, w_eco2825, w_eco2826, w_eco2827, w_eco2828, w_eco2829, w_eco2830, w_eco2831, w_eco2832, w_eco2833, w_eco2834, w_eco2835, w_eco2836, w_eco2837, w_eco2838, w_eco2839, w_eco2840, w_eco2841, w_eco2842, w_eco2843, w_eco2844, w_eco2845, w_eco2846, w_eco2847, w_eco2848, w_eco2849, w_eco2850, w_eco2851, w_eco2852, w_eco2853, w_eco2854, w_eco2855, w_eco2856, w_eco2857, w_eco2858, w_eco2859, w_eco2860, w_eco2861, w_eco2862, w_eco2863, w_eco2864, w_eco2865, w_eco2866, w_eco2867, w_eco2868, w_eco2869, w_eco2870, w_eco2871, w_eco2872, w_eco2873, w_eco2874, w_eco2875, w_eco2876, w_eco2877, w_eco2878, w_eco2879, w_eco2880, w_eco2881, w_eco2882, w_eco2883, w_eco2884, w_eco2885, w_eco2886, w_eco2887, w_eco2888, w_eco2889, w_eco2890, w_eco2891, w_eco2892, w_eco2893, w_eco2894, w_eco2895, w_eco2896, w_eco2897, w_eco2898, w_eco2899, w_eco2900, w_eco2901, w_eco2902, w_eco2903, w_eco2904, w_eco2905, w_eco2906, w_eco2907, w_eco2908, w_eco2909, w_eco2910, w_eco2911, w_eco2912, w_eco2913, w_eco2914, w_eco2915, w_eco2916, w_eco2917, w_eco2918, w_eco2919, w_eco2920, w_eco2921, w_eco2922, w_eco2923, w_eco2924, w_eco2925, w_eco2926, w_eco2927, w_eco2928, w_eco2929, w_eco2930, w_eco2931, w_eco2932, w_eco2933, w_eco2934, w_eco2935, w_eco2936, w_eco2937, w_eco2938, w_eco2939, w_eco2940, w_eco2941, w_eco2942, w_eco2943, w_eco2944, w_eco2945, w_eco2946, w_eco2947, w_eco2948, w_eco2949, w_eco2950, w_eco2951, w_eco2952, w_eco2953, w_eco2954, w_eco2955, w_eco2956, w_eco2957, w_eco2958, w_eco2959, w_eco2960, w_eco2961, w_eco2962, w_eco2963, w_eco2964, w_eco2965, w_eco2966, w_eco2967, w_eco2968, w_eco2969, w_eco2970, w_eco2971, w_eco2972, w_eco2973, w_eco2974, w_eco2975, w_eco2976, w_eco2977, w_eco2978, w_eco2979, w_eco2980, w_eco2981, w_eco2982, w_eco2983, w_eco2984, w_eco2985, w_eco2986, w_eco2987, w_eco2988, w_eco2989, w_eco2990, w_eco2991, w_eco2992, w_eco2993, w_eco2994, w_eco2995, w_eco2996, w_eco2997, w_eco2998, w_eco2999, w_eco3000, w_eco3001, w_eco3002, w_eco3003, w_eco3004, w_eco3005, w_eco3006, w_eco3007, w_eco3008, w_eco3009, w_eco3010, w_eco3011, w_eco3012, w_eco3013, w_eco3014, w_eco3015, w_eco3016, w_eco3017, w_eco3018, w_eco3019, w_eco3020, w_eco3021, w_eco3022, w_eco3023, w_eco3024, w_eco3025, w_eco3026, w_eco3027, w_eco3028, w_eco3029, w_eco3030, w_eco3031, w_eco3032, w_eco3033, w_eco3034, w_eco3035, w_eco3036, w_eco3037, w_eco3038, w_eco3039, w_eco3040, w_eco3041, w_eco3042, w_eco3043, w_eco3044, w_eco3045, w_eco3046, w_eco3047, w_eco3048, w_eco3049, w_eco3050, w_eco3051, w_eco3052, w_eco3053, w_eco3054, w_eco3055, w_eco3056, w_eco3057, w_eco3058, w_eco3059, w_eco3060, w_eco3061, w_eco3062, w_eco3063, w_eco3064, w_eco3065, w_eco3066, w_eco3067, w_eco3068, w_eco3069, w_eco3070, w_eco3071, w_eco3072, w_eco3073, w_eco3074, w_eco3075, w_eco3076, w_eco3077, w_eco3078, w_eco3079, w_eco3080, w_eco3081, w_eco3082, w_eco3083, w_eco3084, w_eco3085, w_eco3086, w_eco3087, w_eco3088, w_eco3089, w_eco3090, w_eco3091, w_eco3092, w_eco3093, w_eco3094, w_eco3095, w_eco3096, w_eco3097, w_eco3098, w_eco3099, w_eco3100, w_eco3101, w_eco3102, w_eco3103, w_eco3104, w_eco3105, w_eco3106, w_eco3107, w_eco3108, w_eco3109, w_eco3110, w_eco3111, w_eco3112, w_eco3113, w_eco3114, w_eco3115, w_eco3116, w_eco3117, w_eco3118, w_eco3119, w_eco3120, w_eco3121, w_eco3122, w_eco3123, w_eco3124, w_eco3125, w_eco3126, w_eco3127, w_eco3128, w_eco3129, w_eco3130, w_eco3131, w_eco3132, w_eco3133, w_eco3134, w_eco3135, w_eco3136, w_eco3137, w_eco3138, w_eco3139, w_eco3140, w_eco3141, w_eco3142, w_eco3143, w_eco3144, w_eco3145, w_eco3146, w_eco3147, w_eco3148, w_eco3149, w_eco3150, w_eco3151, w_eco3152, w_eco3153, w_eco3154, w_eco3155, w_eco3156, w_eco3157, w_eco3158, w_eco3159, w_eco3160, w_eco3161, w_eco3162, w_eco3163, w_eco3164, w_eco3165, w_eco3166, w_eco3167, w_eco3168, w_eco3169, w_eco3170, w_eco3171, w_eco3172, w_eco3173, w_eco3174, w_eco3175, w_eco3176, w_eco3177, w_eco3178, w_eco3179, w_eco3180, w_eco3181, w_eco3182, w_eco3183, w_eco3184, w_eco3185, w_eco3186, w_eco3187, w_eco3188, w_eco3189, w_eco3190, w_eco3191, w_eco3192, w_eco3193, w_eco3194, w_eco3195, w_eco3196, w_eco3197, w_eco3198, w_eco3199, w_eco3200, w_eco3201, w_eco3202, w_eco3203, w_eco3204, w_eco3205, w_eco3206, w_eco3207, w_eco3208, w_eco3209, w_eco3210, w_eco3211, w_eco3212, w_eco3213, w_eco3214, w_eco3215, w_eco3216, w_eco3217, w_eco3218, w_eco3219, w_eco3220, w_eco3221, w_eco3222, w_eco3223, w_eco3224, w_eco3225, w_eco3226, w_eco3227, w_eco3228, w_eco3229, w_eco3230, w_eco3231, w_eco3232, w_eco3233, w_eco3234, w_eco3235, w_eco3236, w_eco3237, w_eco3238, w_eco3239, w_eco3240, w_eco3241, w_eco3242, w_eco3243, w_eco3244, w_eco3245, w_eco3246, w_eco3247, w_eco3248, w_eco3249, w_eco3250, w_eco3251, w_eco3252, w_eco3253, w_eco3254, w_eco3255, w_eco3256, w_eco3257, w_eco3258, w_eco3259, w_eco3260, w_eco3261, w_eco3262, w_eco3263, w_eco3264, w_eco3265, w_eco3266, w_eco3267, w_eco3268, w_eco3269, w_eco3270, w_eco3271, w_eco3272, w_eco3273, w_eco3274, w_eco3275, w_eco3276, w_eco3277, w_eco3278, w_eco3279, w_eco3280, w_eco3281, w_eco3282, w_eco3283, w_eco3284, w_eco3285, w_eco3286, w_eco3287, w_eco3288, w_eco3289, w_eco3290, w_eco3291, w_eco3292, w_eco3293, w_eco3294, w_eco3295, w_eco3296, w_eco3297, w_eco3298, w_eco3299, w_eco3300, w_eco3301, w_eco3302, w_eco3303, w_eco3304, w_eco3305, w_eco3306, w_eco3307, w_eco3308, w_eco3309, w_eco3310, w_eco3311, w_eco3312, w_eco3313, w_eco3314, w_eco3315, w_eco3316, w_eco3317, w_eco3318, w_eco3319, w_eco3320, w_eco3321, w_eco3322, w_eco3323, w_eco3324, w_eco3325, w_eco3326, w_eco3327, w_eco3328, w_eco3329, w_eco3330, w_eco3331, w_eco3332, w_eco3333, w_eco3334, w_eco3335, w_eco3336, w_eco3337, w_eco3338, w_eco3339, w_eco3340, w_eco3341, w_eco3342, w_eco3343, w_eco3344, w_eco3345, w_eco3346, w_eco3347, w_eco3348, w_eco3349, w_eco3350, w_eco3351, w_eco3352, w_eco3353, w_eco3354, w_eco3355, w_eco3356, w_eco3357, w_eco3358, w_eco3359, w_eco3360, w_eco3361, w_eco3362, w_eco3363, w_eco3364, w_eco3365, w_eco3366, w_eco3367, w_eco3368, w_eco3369, w_eco3370, w_eco3371, w_eco3372, w_eco3373, w_eco3374, w_eco3375, w_eco3376, w_eco3377, w_eco3378, w_eco3379, w_eco3380, w_eco3381, w_eco3382, w_eco3383, w_eco3384, w_eco3385, w_eco3386, w_eco3387, w_eco3388, w_eco3389, w_eco3390, w_eco3391, w_eco3392, w_eco3393, w_eco3394, w_eco3395, w_eco3396, w_eco3397, w_eco3398, w_eco3399, w_eco3400, w_eco3401, w_eco3402, w_eco3403, w_eco3404, w_eco3405, w_eco3406, w_eco3407, w_eco3408, w_eco3409, w_eco3410, w_eco3411, w_eco3412, w_eco3413, w_eco3414, w_eco3415, w_eco3416, w_eco3417, w_eco3418, w_eco3419, w_eco3420, w_eco3421, w_eco3422, w_eco3423, w_eco3424, w_eco3425, w_eco3426, w_eco3427, w_eco3428, w_eco3429, w_eco3430, w_eco3431, w_eco3432, w_eco3433, w_eco3434, w_eco3435, w_eco3436, w_eco3437, w_eco3438, w_eco3439, w_eco3440, w_eco3441, w_eco3442, w_eco3443, w_eco3444, w_eco3445, w_eco3446, w_eco3447, w_eco3448, w_eco3449, w_eco3450, w_eco3451, w_eco3452, w_eco3453, w_eco3454, w_eco3455, w_eco3456, w_eco3457, w_eco3458, w_eco3459, w_eco3460, w_eco3461, w_eco3462, w_eco3463, w_eco3464, w_eco3465, w_eco3466, w_eco3467, w_eco3468, w_eco3469, w_eco3470, w_eco3471, w_eco3472, w_eco3473, w_eco3474, w_eco3475, w_eco3476, w_eco3477, w_eco3478, w_eco3479, w_eco3480, w_eco3481, w_eco3482, w_eco3483, w_eco3484, w_eco3485, w_eco3486, w_eco3487, w_eco3488, w_eco3489, w_eco3490, w_eco3491, w_eco3492, w_eco3493, w_eco3494, w_eco3495, w_eco3496, w_eco3497, w_eco3498, w_eco3499, w_eco3500, w_eco3501, w_eco3502, w_eco3503, w_eco3504, w_eco3505, w_eco3506, w_eco3507, w_eco3508, w_eco3509, w_eco3510, w_eco3511, w_eco3512, w_eco3513, w_eco3514, w_eco3515, w_eco3516, w_eco3517, w_eco3518, w_eco3519, w_eco3520, w_eco3521, w_eco3522, w_eco3523, w_eco3524, w_eco3525, w_eco3526, w_eco3527, w_eco3528, w_eco3529, w_eco3530, w_eco3531, w_eco3532, w_eco3533, w_eco3534, w_eco3535, w_eco3536, w_eco3537, w_eco3538, w_eco3539, w_eco3540, w_eco3541, w_eco3542, w_eco3543, w_eco3544, w_eco3545, w_eco3546, w_eco3547, w_eco3548, w_eco3549, w_eco3550, w_eco3551, w_eco3552, w_eco3553, w_eco3554, w_eco3555, w_eco3556, w_eco3557, w_eco3558, w_eco3559, w_eco3560, w_eco3561, w_eco3562, w_eco3563, w_eco3564, w_eco3565, w_eco3566, w_eco3567, w_eco3568, w_eco3569, w_eco3570, w_eco3571, w_eco3572, w_eco3573, w_eco3574, w_eco3575, w_eco3576, w_eco3577, w_eco3578, w_eco3579, w_eco3580, w_eco3581, w_eco3582, w_eco3583, w_eco3584, w_eco3585, w_eco3586, w_eco3587, w_eco3588, w_eco3589, w_eco3590, w_eco3591, w_eco3592, w_eco3593, w_eco3594, w_eco3595, w_eco3596, w_eco3597, w_eco3598, w_eco3599, w_eco3600, w_eco3601, w_eco3602, w_eco3603, w_eco3604, w_eco3605, w_eco3606, w_eco3607, w_eco3608, w_eco3609, w_eco3610, w_eco3611, w_eco3612, w_eco3613, w_eco3614, w_eco3615, w_eco3616, w_eco3617, w_eco3618, w_eco3619, w_eco3620, w_eco3621, w_eco3622, w_eco3623, w_eco3624, w_eco3625, w_eco3626, w_eco3627, w_eco3628, w_eco3629, w_eco3630, w_eco3631, w_eco3632, w_eco3633, w_eco3634, w_eco3635, w_eco3636, w_eco3637, w_eco3638, w_eco3639, w_eco3640, w_eco3641, w_eco3642, w_eco3643, w_eco3644, w_eco3645, w_eco3646, w_eco3647, w_eco3648, w_eco3649, w_eco3650, w_eco3651, w_eco3652, w_eco3653, w_eco3654, w_eco3655, w_eco3656, w_eco3657, w_eco3658, w_eco3659, w_eco3660, w_eco3661, w_eco3662, w_eco3663, w_eco3664, w_eco3665, w_eco3666, w_eco3667, w_eco3668, w_eco3669, w_eco3670, w_eco3671, w_eco3672, w_eco3673, w_eco3674, w_eco3675, w_eco3676, w_eco3677, w_eco3678, w_eco3679, w_eco3680, w_eco3681, w_eco3682, w_eco3683, w_eco3684, w_eco3685, w_eco3686, w_eco3687, w_eco3688, w_eco3689, w_eco3690, w_eco3691, w_eco3692, w_eco3693, w_eco3694, w_eco3695, w_eco3696, w_eco3697, w_eco3698, w_eco3699, w_eco3700, w_eco3701, w_eco3702, w_eco3703, w_eco3704, w_eco3705, w_eco3706, w_eco3707, w_eco3708, w_eco3709, w_eco3710, w_eco3711, w_eco3712, w_eco3713, w_eco3714, w_eco3715, w_eco3716, w_eco3717, w_eco3718, w_eco3719, w_eco3720, w_eco3721, w_eco3722, w_eco3723, w_eco3724, w_eco3725, w_eco3726, w_eco3727, w_eco3728, w_eco3729, w_eco3730, w_eco3731, w_eco3732, w_eco3733, w_eco3734, w_eco3735, w_eco3736, w_eco3737, w_eco3738, w_eco3739, w_eco3740, w_eco3741, w_eco3742, w_eco3743, w_eco3744, w_eco3745, w_eco3746, w_eco3747, w_eco3748, w_eco3749, w_eco3750, w_eco3751, w_eco3752, w_eco3753, w_eco3754, w_eco3755, w_eco3756, w_eco3757, w_eco3758, w_eco3759, w_eco3760, w_eco3761, w_eco3762, w_eco3763, w_eco3764, w_eco3765, w_eco3766, w_eco3767, w_eco3768, w_eco3769, w_eco3770, w_eco3771, w_eco3772, w_eco3773, w_eco3774, w_eco3775, w_eco3776, w_eco3777, w_eco3778, w_eco3779, w_eco3780, w_eco3781, w_eco3782, w_eco3783, w_eco3784, w_eco3785, w_eco3786, w_eco3787, w_eco3788, w_eco3789, w_eco3790, w_eco3791, w_eco3792, w_eco3793, w_eco3794, w_eco3795, w_eco3796, w_eco3797, w_eco3798, w_eco3799, w_eco3800, w_eco3801, w_eco3802, w_eco3803, w_eco3804, w_eco3805, w_eco3806, w_eco3807, w_eco3808, w_eco3809, w_eco3810, w_eco3811, w_eco3812, w_eco3813, w_eco3814, w_eco3815, w_eco3816, w_eco3817, w_eco3818, w_eco3819, w_eco3820, w_eco3821, w_eco3822, w_eco3823, w_eco3824, w_eco3825, w_eco3826, w_eco3827, w_eco3828, w_eco3829, w_eco3830, w_eco3831, w_eco3832, w_eco3833, w_eco3834, w_eco3835, w_eco3836, w_eco3837, w_eco3838, w_eco3839, w_eco3840, w_eco3841, w_eco3842, w_eco3843, w_eco3844, w_eco3845, w_eco3846, w_eco3847, w_eco3848, w_eco3849, w_eco3850, w_eco3851, w_eco3852, w_eco3853, w_eco3854, w_eco3855, w_eco3856, w_eco3857, w_eco3858, w_eco3859, w_eco3860, w_eco3861, w_eco3862, w_eco3863, w_eco3864, w_eco3865, w_eco3866, w_eco3867, w_eco3868, w_eco3869, w_eco3870, w_eco3871, w_eco3872, w_eco3873, w_eco3874, w_eco3875, w_eco3876, w_eco3877, w_eco3878, w_eco3879, w_eco3880, w_eco3881, w_eco3882, w_eco3883, w_eco3884, w_eco3885, w_eco3886, w_eco3887, w_eco3888, w_eco3889, w_eco3890, w_eco3891, w_eco3892, w_eco3893, w_eco3894, w_eco3895, w_eco3896, w_eco3897, w_eco3898, w_eco3899, w_eco3900, sub_wire4, w_eco3901, w_eco3902, w_eco3903, w_eco3904, w_eco3905, w_eco3906, w_eco3907, w_eco3908, w_eco3909, w_eco3910, w_eco3911, w_eco3912, w_eco3913, w_eco3914, w_eco3915, w_eco3916, w_eco3917, w_eco3918, w_eco3919, w_eco3920, w_eco3921, w_eco3922, w_eco3923, w_eco3924, w_eco3925, w_eco3926, w_eco3927, w_eco3928, w_eco3929, w_eco3930, w_eco3931, w_eco3932, w_eco3933, w_eco3934, w_eco3935, w_eco3936, w_eco3937, w_eco3938, w_eco3939, w_eco3940, w_eco3941, w_eco3942, w_eco3943, w_eco3944, w_eco3945, w_eco3946, w_eco3947, w_eco3948, w_eco3949, w_eco3950, w_eco3951, w_eco3952, w_eco3953, w_eco3954, w_eco3955, w_eco3956, w_eco3957, w_eco3958, w_eco3959, w_eco3960, w_eco3961, w_eco3962, w_eco3963, w_eco3964, w_eco3965, w_eco3966, w_eco3967, w_eco3968, w_eco3969, w_eco3970, w_eco3971, w_eco3972, w_eco3973, w_eco3974, w_eco3975, w_eco3976, w_eco3977, w_eco3978, w_eco3979, w_eco3980, w_eco3981, w_eco3982, w_eco3983, w_eco3984, w_eco3985, w_eco3986, w_eco3987, w_eco3988, w_eco3989, w_eco3990, w_eco3991, w_eco3992, w_eco3993, w_eco3994, w_eco3995, w_eco3996, w_eco3997, w_eco3998, w_eco3999, w_eco4000, w_eco4001, w_eco4002, w_eco4003, w_eco4004, w_eco4005, w_eco4006, w_eco4007, w_eco4008, w_eco4009, w_eco4010, w_eco4011, w_eco4012, w_eco4013, w_eco4014, w_eco4015, w_eco4016, w_eco4017, w_eco4018, w_eco4019, w_eco4020, w_eco4021, w_eco4022, w_eco4023, w_eco4024, w_eco4025, w_eco4026, w_eco4027, w_eco4028, w_eco4029, w_eco4030, w_eco4031, w_eco4032, w_eco4033, w_eco4034, w_eco4035, w_eco4036, w_eco4037, w_eco4038, w_eco4039, w_eco4040, w_eco4041, w_eco4042, w_eco4043, w_eco4044, w_eco4045, w_eco4046, w_eco4047, w_eco4048, w_eco4049, w_eco4050, w_eco4051, w_eco4052, w_eco4053, w_eco4054, w_eco4055, w_eco4056, w_eco4057, w_eco4058, w_eco4059, w_eco4060, w_eco4061, w_eco4062, w_eco4063, w_eco4064, w_eco4065, w_eco4066, w_eco4067, w_eco4068, w_eco4069, w_eco4070, w_eco4071, w_eco4072, w_eco4073, w_eco4074, w_eco4075, w_eco4076, w_eco4077, w_eco4078, w_eco4079, w_eco4080, w_eco4081, w_eco4082, w_eco4083, w_eco4084, w_eco4085, w_eco4086, w_eco4087, w_eco4088, w_eco4089, w_eco4090, w_eco4091, w_eco4092, w_eco4093, w_eco4094, w_eco4095, w_eco4096, w_eco4097, w_eco4098, w_eco4099, w_eco4100, w_eco4101, w_eco4102, w_eco4103, w_eco4104, w_eco4105, w_eco4106, w_eco4107, w_eco4108, w_eco4109, w_eco4110, w_eco4111, w_eco4112, w_eco4113, w_eco4114, w_eco4115, w_eco4116, w_eco4117, w_eco4118, w_eco4119, w_eco4120, w_eco4121, w_eco4122, w_eco4123, w_eco4124, w_eco4125, w_eco4126, w_eco4127, w_eco4128, w_eco4129, w_eco4130, w_eco4131, w_eco4132, w_eco4133, w_eco4134, w_eco4135, w_eco4136, w_eco4137, w_eco4138, w_eco4139, w_eco4140, w_eco4141, w_eco4142, w_eco4143, w_eco4144, w_eco4145, w_eco4146, w_eco4147, w_eco4148, w_eco4149, w_eco4150, w_eco4151, w_eco4152, w_eco4153, w_eco4154, w_eco4155, w_eco4156, w_eco4157, w_eco4158, w_eco4159, w_eco4160, w_eco4161, w_eco4162, w_eco4163, w_eco4164, w_eco4165, w_eco4166, w_eco4167, w_eco4168, w_eco4169, w_eco4170, w_eco4171, w_eco4172, w_eco4173, w_eco4174, w_eco4175, w_eco4176, w_eco4177, w_eco4178, w_eco4179, w_eco4180, w_eco4181, w_eco4182, w_eco4183, w_eco4184, w_eco4185, w_eco4186, w_eco4187, w_eco4188, w_eco4189, w_eco4190, w_eco4191, w_eco4192, w_eco4193, w_eco4194, w_eco4195, w_eco4196, w_eco4197, w_eco4198, w_eco4199, w_eco4200, w_eco4201, w_eco4202, w_eco4203, w_eco4204, w_eco4205, w_eco4206, w_eco4207, w_eco4208, w_eco4209, w_eco4210, w_eco4211, w_eco4212, w_eco4213, w_eco4214, w_eco4215, w_eco4216, w_eco4217, w_eco4218, w_eco4219, w_eco4220, w_eco4221, w_eco4222, w_eco4223, w_eco4224, w_eco4225, w_eco4226, w_eco4227, w_eco4228, w_eco4229, w_eco4230, w_eco4231, w_eco4232, w_eco4233, w_eco4234, w_eco4235, w_eco4236, w_eco4237, w_eco4238, w_eco4239, w_eco4240, w_eco4241, w_eco4242, w_eco4243, w_eco4244, w_eco4245, w_eco4246, w_eco4247, w_eco4248, w_eco4249, w_eco4250, w_eco4251, w_eco4252, w_eco4253, w_eco4254, w_eco4255, w_eco4256, w_eco4257, w_eco4258, w_eco4259, w_eco4260, w_eco4261, w_eco4262, w_eco4263, w_eco4264, w_eco4265, w_eco4266, w_eco4267, w_eco4268, w_eco4269, w_eco4270, w_eco4271, w_eco4272, w_eco4273, w_eco4274, w_eco4275, w_eco4276, w_eco4277, w_eco4278, w_eco4279, w_eco4280, w_eco4281, w_eco4282, w_eco4283, w_eco4284, w_eco4285, w_eco4286, w_eco4287, w_eco4288, w_eco4289, w_eco4290, w_eco4291, w_eco4292, w_eco4293, w_eco4294, w_eco4295, w_eco4296, w_eco4297, w_eco4298, w_eco4299, w_eco4300, w_eco4301, w_eco4302, w_eco4303, w_eco4304, w_eco4305, w_eco4306, w_eco4307, w_eco4308, w_eco4309, w_eco4310, w_eco4311, w_eco4312, w_eco4313, w_eco4314, w_eco4315, w_eco4316, w_eco4317, w_eco4318, w_eco4319, w_eco4320, w_eco4321, w_eco4322, w_eco4323, w_eco4324, w_eco4325, w_eco4326, w_eco4327, w_eco4328, w_eco4329, w_eco4330, w_eco4331, w_eco4332, w_eco4333, w_eco4334, w_eco4335, w_eco4336, w_eco4337, w_eco4338, w_eco4339, w_eco4340, w_eco4341, w_eco4342, w_eco4343, w_eco4344, w_eco4345, w_eco4346, w_eco4347, w_eco4348, w_eco4349, w_eco4350, w_eco4351, w_eco4352, w_eco4353, w_eco4354, w_eco4355, w_eco4356, w_eco4357, w_eco4358, w_eco4359, w_eco4360, w_eco4361, w_eco4362, w_eco4363, w_eco4364, w_eco4365, w_eco4366, w_eco4367, w_eco4368, w_eco4369, w_eco4370, w_eco4371, w_eco4372, w_eco4373, w_eco4374, w_eco4375, w_eco4376, w_eco4377, w_eco4378, w_eco4379, w_eco4380, w_eco4381, w_eco4382, w_eco4383, w_eco4384, w_eco4385, w_eco4386, w_eco4387, w_eco4388, w_eco4389, w_eco4390, w_eco4391, w_eco4392, w_eco4393, w_eco4394, w_eco4395, w_eco4396, w_eco4397, w_eco4398, w_eco4399, w_eco4400, w_eco4401, w_eco4402, w_eco4403, w_eco4404, w_eco4405, w_eco4406, w_eco4407, w_eco4408, w_eco4409, w_eco4410, w_eco4411, w_eco4412, w_eco4413, w_eco4414, w_eco4415, w_eco4416, w_eco4417, w_eco4418, w_eco4419, w_eco4420, w_eco4421, w_eco4422, w_eco4423, w_eco4424, w_eco4425, w_eco4426, w_eco4427, w_eco4428, w_eco4429, w_eco4430, w_eco4431, w_eco4432, w_eco4433, w_eco4434, w_eco4435, w_eco4436, w_eco4437, w_eco4438, w_eco4439, w_eco4440, w_eco4441, w_eco4442, w_eco4443, w_eco4444, w_eco4445, w_eco4446, w_eco4447, w_eco4448, w_eco4449, w_eco4450, w_eco4451, w_eco4452, w_eco4453, w_eco4454, w_eco4455, w_eco4456, w_eco4457, w_eco4458, w_eco4459, w_eco4460, w_eco4461, w_eco4462, w_eco4463, w_eco4464, w_eco4465, w_eco4466, w_eco4467, w_eco4468, w_eco4469, w_eco4470, w_eco4471, w_eco4472, w_eco4473, w_eco4474, w_eco4475, w_eco4476, w_eco4477, w_eco4478, w_eco4479, w_eco4480, w_eco4481, w_eco4482, w_eco4483, w_eco4484, w_eco4485, w_eco4486, w_eco4487, w_eco4488, w_eco4489, w_eco4490, w_eco4491, w_eco4492, w_eco4493, w_eco4494, w_eco4495, w_eco4496, w_eco4497, w_eco4498, w_eco4499, w_eco4500, w_eco4501, w_eco4502, w_eco4503, w_eco4504, w_eco4505, w_eco4506, w_eco4507, w_eco4508, w_eco4509, w_eco4510, w_eco4511, w_eco4512, w_eco4513, w_eco4514, w_eco4515, w_eco4516, w_eco4517, w_eco4518, w_eco4519, w_eco4520, w_eco4521, w_eco4522, w_eco4523, w_eco4524, w_eco4525, w_eco4526, w_eco4527, w_eco4528, w_eco4529, w_eco4530, w_eco4531, w_eco4532, w_eco4533, w_eco4534, w_eco4535, w_eco4536, w_eco4537, w_eco4538, w_eco4539, w_eco4540, w_eco4541, w_eco4542, w_eco4543, w_eco4544, w_eco4545, w_eco4546, w_eco4547, w_eco4548, w_eco4549, w_eco4550, w_eco4551, w_eco4552, w_eco4553, w_eco4554, w_eco4555, w_eco4556, w_eco4557, w_eco4558, w_eco4559, w_eco4560, w_eco4561, w_eco4562, w_eco4563, w_eco4564, w_eco4565, w_eco4566, w_eco4567, w_eco4568, w_eco4569, w_eco4570, w_eco4571, w_eco4572, w_eco4573, w_eco4574, w_eco4575, w_eco4576, w_eco4577, w_eco4578, w_eco4579, w_eco4580, w_eco4581, w_eco4582, w_eco4583, w_eco4584, w_eco4585, w_eco4586, w_eco4587, w_eco4588, w_eco4589, w_eco4590, w_eco4591, w_eco4592, w_eco4593, w_eco4594, w_eco4595, w_eco4596, w_eco4597, w_eco4598, w_eco4599, w_eco4600, w_eco4601, w_eco4602, w_eco4603, w_eco4604, w_eco4605, w_eco4606, w_eco4607, w_eco4608, w_eco4609, w_eco4610, w_eco4611, w_eco4612, w_eco4613, w_eco4614, w_eco4615, w_eco4616, w_eco4617, w_eco4618, w_eco4619, w_eco4620, w_eco4621, w_eco4622, w_eco4623, w_eco4624, w_eco4625, w_eco4626, w_eco4627, w_eco4628, w_eco4629, w_eco4630, w_eco4631, w_eco4632, w_eco4633, w_eco4634, w_eco4635, w_eco4636, w_eco4637, w_eco4638, w_eco4639, w_eco4640, w_eco4641, w_eco4642, w_eco4643, w_eco4644, w_eco4645, w_eco4646, w_eco4647, w_eco4648, w_eco4649, w_eco4650, w_eco4651, w_eco4652, w_eco4653, w_eco4654, w_eco4655, w_eco4656, w_eco4657, w_eco4658, w_eco4659, w_eco4660, w_eco4661, w_eco4662, w_eco4663, w_eco4664, w_eco4665, w_eco4666, w_eco4667, w_eco4668, w_eco4669, w_eco4670, w_eco4671, w_eco4672, w_eco4673, w_eco4674, w_eco4675, w_eco4676, w_eco4677, w_eco4678, w_eco4679, w_eco4680, w_eco4681, w_eco4682, w_eco4683, w_eco4684, w_eco4685, w_eco4686, w_eco4687, w_eco4688, w_eco4689, w_eco4690, w_eco4691, w_eco4692, w_eco4693, w_eco4694, w_eco4695, w_eco4696, w_eco4697, w_eco4698, w_eco4699, w_eco4700, w_eco4701, w_eco4702, w_eco4703, w_eco4704, w_eco4705, w_eco4706, w_eco4707, w_eco4708, w_eco4709, w_eco4710, w_eco4711, w_eco4712, w_eco4713, w_eco4714, w_eco4715, w_eco4716, w_eco4717, w_eco4718, w_eco4719, w_eco4720, w_eco4721, w_eco4722, w_eco4723, w_eco4724, w_eco4725, w_eco4726, w_eco4727, w_eco4728, w_eco4729, w_eco4730, w_eco4731, w_eco4732, w_eco4733, w_eco4734, w_eco4735, w_eco4736, w_eco4737, w_eco4738, w_eco4739, w_eco4740, w_eco4741, w_eco4742, w_eco4743, w_eco4744, w_eco4745, w_eco4746, w_eco4747, w_eco4748, w_eco4749, w_eco4750, w_eco4751, w_eco4752, w_eco4753, w_eco4754, w_eco4755, w_eco4756, w_eco4757, w_eco4758, w_eco4759, w_eco4760, w_eco4761, w_eco4762, w_eco4763, w_eco4764, w_eco4765, w_eco4766, w_eco4767, w_eco4768, w_eco4769, w_eco4770, w_eco4771, w_eco4772, w_eco4773, w_eco4774, w_eco4775, w_eco4776, w_eco4777, w_eco4778, w_eco4779, w_eco4780, w_eco4781, w_eco4782, w_eco4783, w_eco4784, w_eco4785, w_eco4786, w_eco4787, w_eco4788, w_eco4789, w_eco4790, w_eco4791, w_eco4792, w_eco4793, w_eco4794, w_eco4795, w_eco4796, w_eco4797, w_eco4798, w_eco4799, w_eco4800, w_eco4801, w_eco4802, w_eco4803, w_eco4804, w_eco4805, w_eco4806, w_eco4807, w_eco4808, w_eco4809, w_eco4810, w_eco4811, w_eco4812, w_eco4813, w_eco4814, w_eco4815, w_eco4816, w_eco4817, w_eco4818, w_eco4819, w_eco4820, w_eco4821, w_eco4822, w_eco4823, w_eco4824, w_eco4825, w_eco4826, w_eco4827, w_eco4828, w_eco4829, w_eco4830, w_eco4831, w_eco4832, w_eco4833, w_eco4834, w_eco4835, w_eco4836, w_eco4837, w_eco4838, w_eco4839, w_eco4840, w_eco4841, w_eco4842, w_eco4843, w_eco4844, w_eco4845, w_eco4846, w_eco4847, w_eco4848, w_eco4849, w_eco4850, w_eco4851, w_eco4852, w_eco4853, w_eco4854, w_eco4855, w_eco4856, w_eco4857, w_eco4858, w_eco4859, w_eco4860, w_eco4861, w_eco4862, w_eco4863, w_eco4864, w_eco4865, w_eco4866, w_eco4867, w_eco4868, w_eco4869, w_eco4870, w_eco4871, w_eco4872, w_eco4873, w_eco4874, w_eco4875, w_eco4876, w_eco4877, w_eco4878, w_eco4879, w_eco4880, w_eco4881, w_eco4882, w_eco4883, w_eco4884, w_eco4885, w_eco4886, w_eco4887, w_eco4888, w_eco4889, w_eco4890, w_eco4891, w_eco4892, w_eco4893, w_eco4894, w_eco4895, w_eco4896, w_eco4897, w_eco4898, w_eco4899, w_eco4900, w_eco4901, w_eco4902, w_eco4903, w_eco4904, w_eco4905, w_eco4906, w_eco4907, w_eco4908, w_eco4909, w_eco4910, w_eco4911, w_eco4912, w_eco4913, w_eco4914, w_eco4915, w_eco4916, w_eco4917, w_eco4918, w_eco4919, w_eco4920, w_eco4921, w_eco4922, w_eco4923, w_eco4924, w_eco4925, w_eco4926, w_eco4927, w_eco4928, w_eco4929, w_eco4930, w_eco4931, w_eco4932, w_eco4933, w_eco4934, w_eco4935, w_eco4936, w_eco4937, w_eco4938, w_eco4939, w_eco4940, w_eco4941, w_eco4942, w_eco4943, w_eco4944, w_eco4945, w_eco4946, w_eco4947, w_eco4948, w_eco4949, w_eco4950, w_eco4951, w_eco4952, w_eco4953, w_eco4954, w_eco4955, w_eco4956, w_eco4957, w_eco4958, w_eco4959, w_eco4960, w_eco4961, w_eco4962, w_eco4963, w_eco4964, w_eco4965, w_eco4966, w_eco4967, w_eco4968, w_eco4969, w_eco4970, w_eco4971, w_eco4972, w_eco4973, w_eco4974, w_eco4975, w_eco4976, w_eco4977, w_eco4978, w_eco4979, w_eco4980, w_eco4981, w_eco4982, w_eco4983, w_eco4984, w_eco4985, w_eco4986, w_eco4987, w_eco4988, w_eco4989, w_eco4990, w_eco4991, w_eco4992, w_eco4993, w_eco4994, w_eco4995, w_eco4996, w_eco4997, w_eco4998, w_eco4999, w_eco5000, w_eco5001, w_eco5002, w_eco5003, w_eco5004, w_eco5005, w_eco5006, w_eco5007, w_eco5008, w_eco5009, w_eco5010, w_eco5011, w_eco5012, w_eco5013, w_eco5014, w_eco5015, w_eco5016, w_eco5017, w_eco5018, w_eco5019, w_eco5020, w_eco5021, w_eco5022, w_eco5023, w_eco5024, w_eco5025, w_eco5026, w_eco5027, w_eco5028, w_eco5029, w_eco5030, w_eco5031, w_eco5032, w_eco5033, w_eco5034, w_eco5035, w_eco5036, w_eco5037, w_eco5038, w_eco5039, w_eco5040, w_eco5041, w_eco5042, w_eco5043, w_eco5044, w_eco5045, w_eco5046, w_eco5047, w_eco5048, w_eco5049, w_eco5050, w_eco5051, w_eco5052, w_eco5053, w_eco5054, w_eco5055, w_eco5056, w_eco5057, w_eco5058, w_eco5059, w_eco5060, w_eco5061, w_eco5062, w_eco5063, w_eco5064, w_eco5065, w_eco5066, w_eco5067, w_eco5068, w_eco5069, w_eco5070, w_eco5071, w_eco5072, w_eco5073, w_eco5074, w_eco5075, w_eco5076, w_eco5077, w_eco5078, w_eco5079, w_eco5080, w_eco5081, w_eco5082, w_eco5083, w_eco5084, w_eco5085, w_eco5086, w_eco5087, w_eco5088, w_eco5089, w_eco5090, w_eco5091, w_eco5092, w_eco5093, w_eco5094, w_eco5095, w_eco5096, w_eco5097, w_eco5098, w_eco5099, w_eco5100, w_eco5101, w_eco5102, w_eco5103, w_eco5104, w_eco5105, w_eco5106, w_eco5107, w_eco5108, w_eco5109, w_eco5110, w_eco5111, w_eco5112, w_eco5113, w_eco5114, w_eco5115, w_eco5116, w_eco5117, w_eco5118, w_eco5119, w_eco5120, w_eco5121, w_eco5122, w_eco5123, w_eco5124, w_eco5125, w_eco5126, w_eco5127, w_eco5128, w_eco5129, w_eco5130, w_eco5131, w_eco5132, w_eco5133, w_eco5134, w_eco5135, w_eco5136, w_eco5137, w_eco5138, w_eco5139, w_eco5140, w_eco5141, w_eco5142, w_eco5143, w_eco5144, w_eco5145, w_eco5146, w_eco5147, w_eco5148, w_eco5149, w_eco5150, w_eco5151, w_eco5152, w_eco5153, w_eco5154, w_eco5155, w_eco5156, w_eco5157, w_eco5158, w_eco5159, w_eco5160, w_eco5161, w_eco5162, w_eco5163, w_eco5164, w_eco5165, w_eco5166, w_eco5167, w_eco5168, w_eco5169, w_eco5170, w_eco5171, w_eco5172, w_eco5173, w_eco5174, w_eco5175, w_eco5176, w_eco5177, w_eco5178, w_eco5179, w_eco5180, w_eco5181, w_eco5182, w_eco5183, w_eco5184, w_eco5185, w_eco5186, w_eco5187, w_eco5188, w_eco5189, w_eco5190, w_eco5191, w_eco5192, w_eco5193, w_eco5194, w_eco5195, w_eco5196, w_eco5197, w_eco5198, w_eco5199, w_eco5200, w_eco5201, w_eco5202, w_eco5203, w_eco5204, w_eco5205, w_eco5206, w_eco5207, w_eco5208, w_eco5209, w_eco5210, w_eco5211, w_eco5212, w_eco5213, w_eco5214, w_eco5215, w_eco5216, w_eco5217, w_eco5218, w_eco5219, w_eco5220, w_eco5221, w_eco5222, w_eco5223, w_eco5224, w_eco5225, w_eco5226, w_eco5227, w_eco5228, w_eco5229, w_eco5230, w_eco5231, w_eco5232, w_eco5233, w_eco5234, w_eco5235, w_eco5236, w_eco5237, w_eco5238, w_eco5239, w_eco5240, w_eco5241, w_eco5242, w_eco5243, w_eco5244, w_eco5245, w_eco5246, w_eco5247, w_eco5248, w_eco5249, w_eco5250, w_eco5251, w_eco5252, w_eco5253, w_eco5254, w_eco5255, w_eco5256, w_eco5257, w_eco5258, w_eco5259, w_eco5260, w_eco5261, w_eco5262, w_eco5263, w_eco5264, w_eco5265, w_eco5266, w_eco5267, w_eco5268, w_eco5269, w_eco5270, w_eco5271, w_eco5272, w_eco5273, w_eco5274, w_eco5275, w_eco5276, w_eco5277, w_eco5278, w_eco5279, w_eco5280, w_eco5281, w_eco5282, w_eco5283, w_eco5284, w_eco5285, w_eco5286, w_eco5287, w_eco5288, w_eco5289, w_eco5290, w_eco5291, w_eco5292, w_eco5293, w_eco5294, w_eco5295, w_eco5296, w_eco5297, w_eco5298, w_eco5299, w_eco5300, w_eco5301, w_eco5302, w_eco5303, w_eco5304, w_eco5305, w_eco5306, w_eco5307, w_eco5308, w_eco5309, w_eco5310, w_eco5311, w_eco5312, w_eco5313, w_eco5314, w_eco5315, w_eco5316, w_eco5317, w_eco5318, w_eco5319, w_eco5320, w_eco5321, w_eco5322, w_eco5323, w_eco5324, w_eco5325, w_eco5326, w_eco5327, w_eco5328, w_eco5329, w_eco5330, w_eco5331, w_eco5332, w_eco5333, w_eco5334, w_eco5335, w_eco5336, w_eco5337, w_eco5338, w_eco5339, w_eco5340, w_eco5341, w_eco5342, w_eco5343, w_eco5344, w_eco5345, w_eco5346, w_eco5347, w_eco5348, w_eco5349, w_eco5350, w_eco5351, w_eco5352, w_eco5353, w_eco5354, w_eco5355, w_eco5356, w_eco5357, w_eco5358, w_eco5359, w_eco5360, w_eco5361, w_eco5362, w_eco5363, w_eco5364, w_eco5365, w_eco5366, w_eco5367, w_eco5368, w_eco5369, w_eco5370, w_eco5371, w_eco5372, w_eco5373, w_eco5374, w_eco5375, w_eco5376, w_eco5377, w_eco5378, w_eco5379, w_eco5380, w_eco5381, w_eco5382, w_eco5383, w_eco5384, w_eco5385, w_eco5386, w_eco5387, w_eco5388, w_eco5389, w_eco5390, w_eco5391, w_eco5392, w_eco5393, w_eco5394, w_eco5395, w_eco5396, w_eco5397, w_eco5398, w_eco5399, w_eco5400, w_eco5401, w_eco5402, w_eco5403, w_eco5404, w_eco5405, w_eco5406, w_eco5407, w_eco5408, w_eco5409, w_eco5410, w_eco5411, w_eco5412, w_eco5413, w_eco5414, w_eco5415, w_eco5416, w_eco5417, w_eco5418, w_eco5419, w_eco5420, w_eco5421, w_eco5422, w_eco5423, w_eco5424, w_eco5425, w_eco5426, w_eco5427, w_eco5428, w_eco5429, w_eco5430, w_eco5431, w_eco5432, w_eco5433, w_eco5434, w_eco5435, w_eco5436, w_eco5437, w_eco5438, w_eco5439, w_eco5440, w_eco5441, w_eco5442, w_eco5443, w_eco5444, w_eco5445, w_eco5446, w_eco5447, w_eco5448, w_eco5449, w_eco5450, w_eco5451, w_eco5452, w_eco5453, w_eco5454, w_eco5455, w_eco5456, w_eco5457, w_eco5458, w_eco5459, w_eco5460, w_eco5461, w_eco5462, w_eco5463, w_eco5464, w_eco5465, w_eco5466, w_eco5467, w_eco5468, w_eco5469, w_eco5470, w_eco5471, w_eco5472, w_eco5473, w_eco5474, w_eco5475, w_eco5476, w_eco5477, w_eco5478, w_eco5479, w_eco5480, sub_wire5, w_eco5481, w_eco5482, w_eco5483, w_eco5484, w_eco5485, w_eco5486, w_eco5487, w_eco5488, w_eco5489, w_eco5490, w_eco5491, w_eco5492, w_eco5493, w_eco5494, w_eco5495, w_eco5496, w_eco5497, w_eco5498, w_eco5499, w_eco5500, w_eco5501, w_eco5502, w_eco5503, w_eco5504, w_eco5505, w_eco5506, w_eco5507, w_eco5508, w_eco5509, w_eco5510, w_eco5511, w_eco5512, w_eco5513, w_eco5514, w_eco5515, w_eco5516, w_eco5517, w_eco5518, w_eco5519, w_eco5520, w_eco5521, w_eco5522, w_eco5523, w_eco5524, w_eco5525, w_eco5526, w_eco5527, w_eco5528, w_eco5529, w_eco5530, w_eco5531, w_eco5532, w_eco5533, w_eco5534, w_eco5535, w_eco5536, w_eco5537, w_eco5538, w_eco5539, w_eco5540, w_eco5541, w_eco5542, w_eco5543, w_eco5544, w_eco5545, w_eco5546, w_eco5547, w_eco5548, w_eco5549, w_eco5550, w_eco5551, w_eco5552, w_eco5553, w_eco5554, w_eco5555, w_eco5556, w_eco5557, w_eco5558, w_eco5559, w_eco5560, w_eco5561, w_eco5562, w_eco5563, w_eco5564, w_eco5565, w_eco5566, w_eco5567, w_eco5568, w_eco5569, w_eco5570, w_eco5571, w_eco5572, w_eco5573, w_eco5574, w_eco5575, w_eco5576, w_eco5577, w_eco5578, w_eco5579, w_eco5580, w_eco5581, w_eco5582, w_eco5583, w_eco5584, w_eco5585, w_eco5586, w_eco5587, w_eco5588, w_eco5589, w_eco5590, w_eco5591, w_eco5592, w_eco5593, w_eco5594, w_eco5595, w_eco5596, w_eco5597, w_eco5598, w_eco5599, w_eco5600, w_eco5601, w_eco5602, w_eco5603, w_eco5604, w_eco5605, w_eco5606, w_eco5607, w_eco5608, w_eco5609, w_eco5610, w_eco5611, w_eco5612, w_eco5613, w_eco5614, w_eco5615, w_eco5616, w_eco5617, w_eco5618, w_eco5619, w_eco5620, w_eco5621, w_eco5622, w_eco5623, w_eco5624, w_eco5625, w_eco5626, w_eco5627, w_eco5628, w_eco5629, w_eco5630, w_eco5631, w_eco5632, w_eco5633, w_eco5634, w_eco5635, w_eco5636, w_eco5637, w_eco5638, w_eco5639, w_eco5640, w_eco5641, w_eco5642, w_eco5643, w_eco5644, w_eco5645, w_eco5646, w_eco5647, w_eco5648, w_eco5649, w_eco5650, w_eco5651, w_eco5652, w_eco5653, w_eco5654, w_eco5655, w_eco5656, w_eco5657, w_eco5658, w_eco5659, w_eco5660, w_eco5661, w_eco5662, w_eco5663, w_eco5664, w_eco5665, w_eco5666, w_eco5667, w_eco5668, w_eco5669, w_eco5670, w_eco5671, w_eco5672, w_eco5673, w_eco5674, w_eco5675, w_eco5676, w_eco5677, w_eco5678, w_eco5679, w_eco5680, w_eco5681, w_eco5682, w_eco5683, w_eco5684, w_eco5685, w_eco5686, w_eco5687, w_eco5688, w_eco5689, w_eco5690, w_eco5691, w_eco5692, w_eco5693, w_eco5694, w_eco5695, w_eco5696, w_eco5697, w_eco5698, w_eco5699, w_eco5700, w_eco5701, w_eco5702, w_eco5703, w_eco5704, w_eco5705, w_eco5706, w_eco5707, w_eco5708, w_eco5709, w_eco5710, w_eco5711, w_eco5712, w_eco5713, w_eco5714, w_eco5715, w_eco5716, w_eco5717, w_eco5718, w_eco5719, w_eco5720, w_eco5721, w_eco5722, w_eco5723, w_eco5724, w_eco5725, w_eco5726, w_eco5727, w_eco5728, w_eco5729, w_eco5730, w_eco5731, w_eco5732, w_eco5733, w_eco5734, w_eco5735, w_eco5736, w_eco5737, w_eco5738, w_eco5739, w_eco5740, w_eco5741, w_eco5742, w_eco5743, w_eco5744, w_eco5745, w_eco5746, w_eco5747, w_eco5748, w_eco5749, w_eco5750, w_eco5751, w_eco5752, w_eco5753, w_eco5754, w_eco5755, w_eco5756, w_eco5757, w_eco5758, w_eco5759, w_eco5760, w_eco5761, w_eco5762, w_eco5763, w_eco5764, w_eco5765, w_eco5766, w_eco5767, w_eco5768, w_eco5769, w_eco5770, w_eco5771, w_eco5772, w_eco5773, w_eco5774, w_eco5775, w_eco5776, w_eco5777, w_eco5778, w_eco5779, w_eco5780, w_eco5781, w_eco5782, w_eco5783, w_eco5784, w_eco5785, w_eco5786, w_eco5787, w_eco5788, w_eco5789, w_eco5790, w_eco5791, w_eco5792, w_eco5793, w_eco5794, w_eco5795, w_eco5796, w_eco5797, w_eco5798, w_eco5799, w_eco5800, w_eco5801, w_eco5802, w_eco5803, w_eco5804, w_eco5805, w_eco5806, w_eco5807, w_eco5808, w_eco5809, w_eco5810, w_eco5811, w_eco5812, w_eco5813, w_eco5814, w_eco5815, w_eco5816, w_eco5817, w_eco5818, w_eco5819, w_eco5820, w_eco5821, w_eco5822, w_eco5823, w_eco5824, w_eco5825, w_eco5826, w_eco5827, w_eco5828, w_eco5829, w_eco5830, w_eco5831, w_eco5832, w_eco5833, w_eco5834, w_eco5835, w_eco5836, w_eco5837, w_eco5838, w_eco5839, w_eco5840, w_eco5841, w_eco5842, w_eco5843, w_eco5844, w_eco5845, w_eco5846, w_eco5847, w_eco5848, w_eco5849, w_eco5850, w_eco5851, w_eco5852, w_eco5853, w_eco5854, w_eco5855, w_eco5856, w_eco5857, w_eco5858, w_eco5859, w_eco5860, w_eco5861, w_eco5862, w_eco5863, w_eco5864, w_eco5865, w_eco5866, w_eco5867, w_eco5868, w_eco5869, w_eco5870, w_eco5871, w_eco5872, w_eco5873, w_eco5874, w_eco5875, w_eco5876, w_eco5877, w_eco5878, w_eco5879, w_eco5880, w_eco5881, w_eco5882, w_eco5883, w_eco5884, w_eco5885, w_eco5886, w_eco5887, w_eco5888, w_eco5889, w_eco5890, w_eco5891, w_eco5892, w_eco5893, w_eco5894, w_eco5895, w_eco5896, w_eco5897, w_eco5898, w_eco5899, w_eco5900, w_eco5901, w_eco5902, w_eco5903, w_eco5904, w_eco5905, w_eco5906, w_eco5907, w_eco5908, w_eco5909, w_eco5910, w_eco5911, w_eco5912, w_eco5913, w_eco5914, w_eco5915, w_eco5916, w_eco5917, w_eco5918, w_eco5919, w_eco5920, w_eco5921, w_eco5922, w_eco5923, w_eco5924, w_eco5925, w_eco5926, w_eco5927, w_eco5928, w_eco5929, w_eco5930, w_eco5931, w_eco5932, w_eco5933, w_eco5934, w_eco5935, w_eco5936, w_eco5937, w_eco5938, w_eco5939, w_eco5940, w_eco5941, w_eco5942, w_eco5943, w_eco5944, w_eco5945, w_eco5946, w_eco5947, w_eco5948, w_eco5949, w_eco5950, w_eco5951, w_eco5952, w_eco5953, w_eco5954, w_eco5955, w_eco5956, w_eco5957, w_eco5958, w_eco5959, w_eco5960, w_eco5961, w_eco5962, w_eco5963, w_eco5964, w_eco5965, w_eco5966, w_eco5967, w_eco5968, w_eco5969, w_eco5970, w_eco5971, w_eco5972, w_eco5973, w_eco5974, w_eco5975, w_eco5976, w_eco5977, w_eco5978, w_eco5979, w_eco5980, w_eco5981, w_eco5982, w_eco5983, w_eco5984, w_eco5985, w_eco5986, w_eco5987, w_eco5988, w_eco5989, w_eco5990, w_eco5991, w_eco5992, w_eco5993, w_eco5994, w_eco5995, w_eco5996, w_eco5997, w_eco5998, w_eco5999, w_eco6000, w_eco6001, w_eco6002, w_eco6003, w_eco6004, w_eco6005, w_eco6006, w_eco6007, w_eco6008, w_eco6009, w_eco6010, w_eco6011, w_eco6012, w_eco6013, w_eco6014, w_eco6015, w_eco6016, w_eco6017, w_eco6018, w_eco6019, w_eco6020, w_eco6021, w_eco6022, w_eco6023, w_eco6024, w_eco6025, w_eco6026, w_eco6027, w_eco6028, w_eco6029, w_eco6030, w_eco6031, w_eco6032, w_eco6033, w_eco6034, w_eco6035, w_eco6036, w_eco6037, w_eco6038, w_eco6039, w_eco6040, w_eco6041, w_eco6042, w_eco6043, w_eco6044, w_eco6045, w_eco6046, w_eco6047, w_eco6048, w_eco6049, w_eco6050, w_eco6051, w_eco6052, w_eco6053, w_eco6054, w_eco6055, w_eco6056, w_eco6057, w_eco6058, w_eco6059, w_eco6060, w_eco6061, w_eco6062, w_eco6063, w_eco6064, w_eco6065, w_eco6066, w_eco6067, w_eco6068, w_eco6069, w_eco6070, w_eco6071, w_eco6072, w_eco6073, w_eco6074, w_eco6075, w_eco6076, w_eco6077, w_eco6078, w_eco6079, w_eco6080, w_eco6081, w_eco6082, w_eco6083, w_eco6084, w_eco6085, w_eco6086, w_eco6087, w_eco6088, w_eco6089, w_eco6090, w_eco6091, w_eco6092, w_eco6093, w_eco6094, w_eco6095, w_eco6096, w_eco6097, w_eco6098, w_eco6099, w_eco6100, w_eco6101, w_eco6102, w_eco6103, w_eco6104, w_eco6105, w_eco6106, w_eco6107, w_eco6108, w_eco6109, w_eco6110, w_eco6111, w_eco6112, w_eco6113, w_eco6114, w_eco6115, w_eco6116, w_eco6117, w_eco6118, w_eco6119, w_eco6120, w_eco6121, w_eco6122, w_eco6123, w_eco6124, w_eco6125, w_eco6126, w_eco6127, w_eco6128, w_eco6129, w_eco6130, w_eco6131, w_eco6132, w_eco6133, w_eco6134, w_eco6135, w_eco6136, w_eco6137, w_eco6138, w_eco6139, w_eco6140, w_eco6141, w_eco6142, w_eco6143, w_eco6144, w_eco6145, w_eco6146, w_eco6147, w_eco6148, w_eco6149, w_eco6150, w_eco6151, w_eco6152, w_eco6153, w_eco6154, w_eco6155, w_eco6156, w_eco6157, w_eco6158, w_eco6159, w_eco6160, w_eco6161, w_eco6162, w_eco6163, w_eco6164, w_eco6165, w_eco6166, w_eco6167, w_eco6168, w_eco6169, w_eco6170, w_eco6171, w_eco6172, w_eco6173, w_eco6174, w_eco6175, w_eco6176, w_eco6177, w_eco6178, w_eco6179, w_eco6180, w_eco6181, w_eco6182, w_eco6183, w_eco6184, w_eco6185, w_eco6186, w_eco6187, w_eco6188, w_eco6189, w_eco6190, w_eco6191, w_eco6192, w_eco6193, w_eco6194, w_eco6195, w_eco6196, w_eco6197, w_eco6198, w_eco6199, w_eco6200, w_eco6201, w_eco6202, w_eco6203, w_eco6204, w_eco6205, w_eco6206, w_eco6207, w_eco6208, w_eco6209, w_eco6210, w_eco6211, w_eco6212, w_eco6213, w_eco6214, w_eco6215, w_eco6216, w_eco6217, w_eco6218, w_eco6219, w_eco6220, w_eco6221, w_eco6222, w_eco6223, w_eco6224, w_eco6225, w_eco6226, w_eco6227, w_eco6228, w_eco6229, w_eco6230, w_eco6231, w_eco6232, w_eco6233, w_eco6234, w_eco6235, w_eco6236, w_eco6237, w_eco6238, w_eco6239, w_eco6240, w_eco6241, w_eco6242, w_eco6243, w_eco6244, w_eco6245, w_eco6246, w_eco6247, w_eco6248, w_eco6249, w_eco6250, w_eco6251, w_eco6252, w_eco6253, w_eco6254, w_eco6255, w_eco6256, w_eco6257, w_eco6258, w_eco6259, w_eco6260, w_eco6261, w_eco6262, w_eco6263, w_eco6264, w_eco6265, w_eco6266, w_eco6267, w_eco6268, w_eco6269, w_eco6270, w_eco6271, w_eco6272, w_eco6273, w_eco6274, w_eco6275, w_eco6276, w_eco6277, w_eco6278, w_eco6279, w_eco6280, w_eco6281, w_eco6282, w_eco6283, w_eco6284, w_eco6285, w_eco6286, w_eco6287, w_eco6288, w_eco6289, w_eco6290, w_eco6291, w_eco6292, w_eco6293, w_eco6294, w_eco6295, w_eco6296, w_eco6297, w_eco6298, w_eco6299, w_eco6300, w_eco6301, w_eco6302, w_eco6303, w_eco6304, w_eco6305, w_eco6306, w_eco6307, w_eco6308, w_eco6309, w_eco6310, w_eco6311, w_eco6312, w_eco6313, w_eco6314, w_eco6315, w_eco6316, w_eco6317, w_eco6318, w_eco6319, w_eco6320, w_eco6321, w_eco6322, w_eco6323, w_eco6324, w_eco6325, w_eco6326, w_eco6327, w_eco6328, w_eco6329, w_eco6330, w_eco6331, w_eco6332, w_eco6333, w_eco6334, w_eco6335, w_eco6336, w_eco6337, w_eco6338, w_eco6339, w_eco6340, w_eco6341, w_eco6342, w_eco6343, w_eco6344, w_eco6345, w_eco6346, w_eco6347, w_eco6348, w_eco6349, w_eco6350, w_eco6351, w_eco6352, w_eco6353, w_eco6354, w_eco6355, w_eco6356, w_eco6357, w_eco6358, w_eco6359, w_eco6360, w_eco6361, w_eco6362, w_eco6363, w_eco6364, w_eco6365, w_eco6366, w_eco6367, w_eco6368, w_eco6369, w_eco6370, w_eco6371, w_eco6372, w_eco6373, w_eco6374, w_eco6375, w_eco6376, w_eco6377, w_eco6378, w_eco6379, w_eco6380, w_eco6381, w_eco6382, w_eco6383, w_eco6384, w_eco6385, w_eco6386, w_eco6387, w_eco6388, w_eco6389, w_eco6390, w_eco6391, w_eco6392, w_eco6393, w_eco6394, w_eco6395, w_eco6396, w_eco6397, w_eco6398, w_eco6399, w_eco6400, w_eco6401, w_eco6402, w_eco6403, w_eco6404, w_eco6405, w_eco6406, w_eco6407, w_eco6408, w_eco6409, w_eco6410, w_eco6411, w_eco6412, w_eco6413, w_eco6414, w_eco6415, w_eco6416, w_eco6417, w_eco6418, w_eco6419, w_eco6420, w_eco6421, w_eco6422, w_eco6423, w_eco6424, w_eco6425, w_eco6426, w_eco6427, w_eco6428, w_eco6429, w_eco6430, w_eco6431, w_eco6432, w_eco6433, w_eco6434, w_eco6435, w_eco6436, w_eco6437, w_eco6438, w_eco6439, w_eco6440, w_eco6441, w_eco6442, w_eco6443, w_eco6444, w_eco6445, w_eco6446, w_eco6447, w_eco6448, w_eco6449, w_eco6450, w_eco6451, w_eco6452, w_eco6453, w_eco6454, w_eco6455, w_eco6456, w_eco6457, w_eco6458, w_eco6459, w_eco6460, w_eco6461, w_eco6462, w_eco6463, w_eco6464, w_eco6465, w_eco6466, w_eco6467, w_eco6468, w_eco6469, w_eco6470, w_eco6471, w_eco6472, w_eco6473, w_eco6474, w_eco6475, w_eco6476, w_eco6477, w_eco6478, w_eco6479, w_eco6480, w_eco6481, w_eco6482, w_eco6483, w_eco6484, w_eco6485, w_eco6486, w_eco6487, w_eco6488, w_eco6489, w_eco6490, w_eco6491, w_eco6492, w_eco6493, w_eco6494, w_eco6495, w_eco6496, w_eco6497, w_eco6498, w_eco6499, w_eco6500, w_eco6501, w_eco6502, w_eco6503, w_eco6504, w_eco6505, w_eco6506, w_eco6507, w_eco6508, w_eco6509, w_eco6510, w_eco6511, w_eco6512, w_eco6513, w_eco6514, w_eco6515, w_eco6516, w_eco6517, w_eco6518, w_eco6519, w_eco6520, w_eco6521, w_eco6522, w_eco6523, w_eco6524, w_eco6525, w_eco6526, w_eco6527, w_eco6528, w_eco6529, w_eco6530, w_eco6531, w_eco6532, w_eco6533, w_eco6534, w_eco6535, w_eco6536, w_eco6537, w_eco6538, w_eco6539, w_eco6540, w_eco6541, w_eco6542, w_eco6543, w_eco6544, w_eco6545, w_eco6546, w_eco6547, w_eco6548, w_eco6549, w_eco6550, w_eco6551, w_eco6552, w_eco6553, w_eco6554, w_eco6555, w_eco6556, w_eco6557, w_eco6558, w_eco6559, w_eco6560, w_eco6561, w_eco6562, w_eco6563, w_eco6564, w_eco6565, w_eco6566, w_eco6567, w_eco6568, w_eco6569, w_eco6570, w_eco6571, w_eco6572, w_eco6573, w_eco6574, w_eco6575, w_eco6576, w_eco6577, w_eco6578, w_eco6579, w_eco6580, w_eco6581, w_eco6582, w_eco6583, w_eco6584, w_eco6585, w_eco6586, w_eco6587, w_eco6588, w_eco6589, w_eco6590, w_eco6591, w_eco6592, w_eco6593, w_eco6594, w_eco6595, w_eco6596, w_eco6597, w_eco6598, w_eco6599, w_eco6600, w_eco6601, w_eco6602, w_eco6603, w_eco6604, w_eco6605, w_eco6606, w_eco6607, w_eco6608, w_eco6609, w_eco6610, w_eco6611, w_eco6612, w_eco6613, w_eco6614, w_eco6615, w_eco6616, w_eco6617, w_eco6618, w_eco6619, w_eco6620, w_eco6621, w_eco6622, w_eco6623, w_eco6624, w_eco6625, w_eco6626, w_eco6627, w_eco6628, w_eco6629, w_eco6630, w_eco6631, w_eco6632, w_eco6633, w_eco6634, w_eco6635, w_eco6636, w_eco6637, w_eco6638, w_eco6639, w_eco6640, w_eco6641, w_eco6642, w_eco6643, w_eco6644, w_eco6645, w_eco6646, w_eco6647, w_eco6648, w_eco6649, w_eco6650, w_eco6651, w_eco6652, w_eco6653, w_eco6654, w_eco6655, w_eco6656, w_eco6657, w_eco6658, w_eco6659, w_eco6660, w_eco6661, w_eco6662, w_eco6663, w_eco6664, w_eco6665, w_eco6666, w_eco6667, w_eco6668, w_eco6669, w_eco6670, w_eco6671, w_eco6672, w_eco6673, w_eco6674, w_eco6675, w_eco6676, w_eco6677, w_eco6678, w_eco6679, w_eco6680, w_eco6681, w_eco6682, w_eco6683, w_eco6684, w_eco6685, w_eco6686, w_eco6687, w_eco6688, w_eco6689, w_eco6690, w_eco6691, w_eco6692, w_eco6693, w_eco6694, w_eco6695, w_eco6696, w_eco6697, w_eco6698, w_eco6699, w_eco6700, w_eco6701, w_eco6702, w_eco6703, w_eco6704, w_eco6705, w_eco6706, w_eco6707, w_eco6708, w_eco6709, w_eco6710, w_eco6711, w_eco6712, w_eco6713, w_eco6714, w_eco6715, w_eco6716, w_eco6717, w_eco6718, w_eco6719, w_eco6720, w_eco6721, w_eco6722, w_eco6723, w_eco6724, w_eco6725, w_eco6726, w_eco6727, w_eco6728, w_eco6729, w_eco6730, w_eco6731, w_eco6732, w_eco6733, w_eco6734, w_eco6735, w_eco6736, w_eco6737, w_eco6738, w_eco6739, w_eco6740, w_eco6741, w_eco6742, w_eco6743, w_eco6744, w_eco6745, w_eco6746, w_eco6747, w_eco6748, w_eco6749, w_eco6750, w_eco6751, w_eco6752, w_eco6753, w_eco6754, w_eco6755, w_eco6756, w_eco6757, w_eco6758, w_eco6759, w_eco6760, w_eco6761, w_eco6762, w_eco6763, w_eco6764, w_eco6765, w_eco6766, w_eco6767, w_eco6768, w_eco6769, w_eco6770, w_eco6771, w_eco6772, w_eco6773, w_eco6774, w_eco6775, w_eco6776, w_eco6777, w_eco6778, w_eco6779, w_eco6780, w_eco6781, w_eco6782, w_eco6783, w_eco6784, w_eco6785, w_eco6786, w_eco6787, w_eco6788, w_eco6789, w_eco6790, w_eco6791, w_eco6792, w_eco6793, w_eco6794, w_eco6795, w_eco6796, w_eco6797, w_eco6798, w_eco6799, w_eco6800, w_eco6801, w_eco6802, w_eco6803, w_eco6804, w_eco6805, w_eco6806, w_eco6807, w_eco6808, w_eco6809, w_eco6810, w_eco6811, w_eco6812, w_eco6813, w_eco6814, w_eco6815, w_eco6816, w_eco6817, w_eco6818, w_eco6819, w_eco6820, w_eco6821, w_eco6822, w_eco6823, w_eco6824, w_eco6825, w_eco6826, w_eco6827, w_eco6828, w_eco6829, w_eco6830, w_eco6831, w_eco6832, w_eco6833, w_eco6834, w_eco6835, w_eco6836, w_eco6837, w_eco6838, w_eco6839, w_eco6840, w_eco6841, w_eco6842, w_eco6843, w_eco6844, w_eco6845, w_eco6846, w_eco6847, w_eco6848, w_eco6849, w_eco6850, w_eco6851, w_eco6852, w_eco6853, w_eco6854, w_eco6855, w_eco6856, w_eco6857, w_eco6858, w_eco6859, w_eco6860, w_eco6861, w_eco6862, w_eco6863, w_eco6864, w_eco6865, w_eco6866, w_eco6867, w_eco6868, w_eco6869, w_eco6870, w_eco6871, w_eco6872, w_eco6873, w_eco6874, w_eco6875, w_eco6876, w_eco6877, w_eco6878, w_eco6879, w_eco6880, w_eco6881, w_eco6882, w_eco6883, w_eco6884, w_eco6885, w_eco6886, w_eco6887, w_eco6888, w_eco6889, w_eco6890, w_eco6891, w_eco6892, w_eco6893, w_eco6894, w_eco6895, w_eco6896, w_eco6897, w_eco6898, w_eco6899, w_eco6900, w_eco6901, w_eco6902, w_eco6903, w_eco6904, w_eco6905, w_eco6906, w_eco6907, w_eco6908, w_eco6909, w_eco6910, w_eco6911, w_eco6912, w_eco6913, w_eco6914, w_eco6915, w_eco6916, w_eco6917, w_eco6918, w_eco6919, w_eco6920, w_eco6921, w_eco6922, w_eco6923, w_eco6924, w_eco6925, w_eco6926, w_eco6927, w_eco6928, w_eco6929, w_eco6930, w_eco6931, w_eco6932, w_eco6933, w_eco6934, w_eco6935, w_eco6936, w_eco6937, w_eco6938, w_eco6939, w_eco6940, w_eco6941, w_eco6942, w_eco6943, w_eco6944, w_eco6945, w_eco6946, w_eco6947, w_eco6948, w_eco6949, w_eco6950, w_eco6951, w_eco6952, w_eco6953, w_eco6954, w_eco6955, w_eco6956, w_eco6957, w_eco6958, w_eco6959, w_eco6960, w_eco6961, w_eco6962, w_eco6963, w_eco6964, w_eco6965, w_eco6966, w_eco6967, w_eco6968, w_eco6969, w_eco6970, w_eco6971, w_eco6972, w_eco6973, w_eco6974, w_eco6975, w_eco6976, w_eco6977, w_eco6978, w_eco6979, w_eco6980, w_eco6981, w_eco6982, w_eco6983, w_eco6984, w_eco6985, w_eco6986, w_eco6987, w_eco6988, w_eco6989, w_eco6990, w_eco6991, w_eco6992, w_eco6993, w_eco6994, w_eco6995, w_eco6996, w_eco6997, w_eco6998, w_eco6999, w_eco7000, w_eco7001, w_eco7002, w_eco7003, w_eco7004, w_eco7005, w_eco7006, w_eco7007, w_eco7008, w_eco7009, w_eco7010, w_eco7011, w_eco7012, w_eco7013, w_eco7014, w_eco7015, w_eco7016, w_eco7017, w_eco7018, w_eco7019, w_eco7020, w_eco7021, w_eco7022, w_eco7023, w_eco7024, w_eco7025, w_eco7026, w_eco7027, w_eco7028, w_eco7029, w_eco7030, w_eco7031, w_eco7032, w_eco7033, w_eco7034, w_eco7035, w_eco7036, w_eco7037, w_eco7038, w_eco7039, w_eco7040, w_eco7041, w_eco7042, w_eco7043, w_eco7044, w_eco7045, w_eco7046, w_eco7047, w_eco7048, w_eco7049, w_eco7050, w_eco7051, w_eco7052, w_eco7053, w_eco7054, w_eco7055, w_eco7056, w_eco7057, w_eco7058, w_eco7059, w_eco7060, w_eco7061, w_eco7062, w_eco7063, w_eco7064, w_eco7065, w_eco7066, w_eco7067, w_eco7068, w_eco7069, w_eco7070, w_eco7071, w_eco7072, w_eco7073, w_eco7074, w_eco7075, w_eco7076, w_eco7077, w_eco7078, w_eco7079, w_eco7080, w_eco7081, w_eco7082, w_eco7083, w_eco7084, w_eco7085, w_eco7086, w_eco7087, w_eco7088, w_eco7089, w_eco7090, w_eco7091, w_eco7092, w_eco7093, w_eco7094, w_eco7095, w_eco7096, w_eco7097, w_eco7098, w_eco7099, w_eco7100, w_eco7101, w_eco7102, w_eco7103, w_eco7104, w_eco7105, w_eco7106, w_eco7107, w_eco7108, w_eco7109, w_eco7110, w_eco7111, w_eco7112, w_eco7113, w_eco7114, w_eco7115, w_eco7116, w_eco7117, w_eco7118, w_eco7119, w_eco7120, w_eco7121, w_eco7122, w_eco7123, w_eco7124, w_eco7125, w_eco7126, w_eco7127, w_eco7128, w_eco7129, w_eco7130, w_eco7131, w_eco7132, w_eco7133, w_eco7134, w_eco7135, w_eco7136, w_eco7137, w_eco7138, w_eco7139, w_eco7140, w_eco7141, w_eco7142, w_eco7143, w_eco7144, w_eco7145, w_eco7146, w_eco7147, w_eco7148, w_eco7149, w_eco7150, w_eco7151, w_eco7152, w_eco7153, w_eco7154, w_eco7155, w_eco7156, w_eco7157, w_eco7158, w_eco7159, w_eco7160, w_eco7161, w_eco7162, w_eco7163, w_eco7164, w_eco7165, w_eco7166, w_eco7167, w_eco7168, w_eco7169, w_eco7170, w_eco7171, w_eco7172, w_eco7173, w_eco7174, w_eco7175, w_eco7176, w_eco7177, w_eco7178, w_eco7179, w_eco7180, w_eco7181, w_eco7182, w_eco7183, w_eco7184, w_eco7185, w_eco7186, w_eco7187, w_eco7188, w_eco7189, w_eco7190, w_eco7191, w_eco7192, w_eco7193, w_eco7194, w_eco7195, w_eco7196, w_eco7197, w_eco7198, w_eco7199, w_eco7200, w_eco7201, w_eco7202, w_eco7203, w_eco7204, w_eco7205, w_eco7206, w_eco7207, w_eco7208, w_eco7209, w_eco7210, w_eco7211, w_eco7212, w_eco7213, w_eco7214, w_eco7215, w_eco7216, w_eco7217, w_eco7218, w_eco7219, w_eco7220, w_eco7221, w_eco7222, w_eco7223, w_eco7224, w_eco7225, w_eco7226, w_eco7227, w_eco7228, w_eco7229, w_eco7230, w_eco7231, w_eco7232, w_eco7233, w_eco7234, w_eco7235, w_eco7236, w_eco7237, w_eco7238, w_eco7239, w_eco7240, w_eco7241, w_eco7242, w_eco7243, w_eco7244, w_eco7245, w_eco7246, w_eco7247, w_eco7248, w_eco7249, w_eco7250, w_eco7251, w_eco7252, w_eco7253, w_eco7254, w_eco7255, w_eco7256, w_eco7257, w_eco7258, w_eco7259, w_eco7260, w_eco7261, w_eco7262, w_eco7263, w_eco7264, w_eco7265, w_eco7266, w_eco7267, w_eco7268, w_eco7269, w_eco7270, w_eco7271, w_eco7272, w_eco7273, w_eco7274, w_eco7275, w_eco7276, w_eco7277, w_eco7278, w_eco7279, w_eco7280, w_eco7281, w_eco7282, w_eco7283, w_eco7284, w_eco7285, w_eco7286, w_eco7287, w_eco7288, w_eco7289, w_eco7290, w_eco7291, w_eco7292, w_eco7293, w_eco7294, w_eco7295, w_eco7296, w_eco7297, w_eco7298, w_eco7299, w_eco7300, w_eco7301, w_eco7302, w_eco7303, w_eco7304, w_eco7305, w_eco7306, w_eco7307, w_eco7308, w_eco7309, w_eco7310, w_eco7311, w_eco7312, w_eco7313, w_eco7314, w_eco7315, w_eco7316, w_eco7317, w_eco7318, w_eco7319, w_eco7320, w_eco7321, w_eco7322, w_eco7323, w_eco7324, w_eco7325, w_eco7326, w_eco7327, w_eco7328, w_eco7329, w_eco7330, w_eco7331, w_eco7332, w_eco7333, w_eco7334, w_eco7335, w_eco7336, w_eco7337, w_eco7338, w_eco7339, w_eco7340, w_eco7341, w_eco7342, w_eco7343, w_eco7344, w_eco7345, w_eco7346, w_eco7347, w_eco7348, w_eco7349, w_eco7350, w_eco7351, w_eco7352, w_eco7353, w_eco7354, w_eco7355, w_eco7356, w_eco7357, w_eco7358, w_eco7359, w_eco7360, w_eco7361, w_eco7362, w_eco7363, w_eco7364, w_eco7365, w_eco7366, w_eco7367, w_eco7368, w_eco7369, w_eco7370, w_eco7371, w_eco7372, w_eco7373, w_eco7374, w_eco7375, w_eco7376, w_eco7377, w_eco7378, w_eco7379, w_eco7380, w_eco7381, w_eco7382, w_eco7383, w_eco7384, w_eco7385, w_eco7386, w_eco7387, w_eco7388, w_eco7389, w_eco7390, w_eco7391, w_eco7392, w_eco7393, w_eco7394, w_eco7395, w_eco7396, w_eco7397, w_eco7398, w_eco7399, w_eco7400, w_eco7401, w_eco7402, w_eco7403, w_eco7404, w_eco7405, w_eco7406, w_eco7407, w_eco7408, w_eco7409, w_eco7410, w_eco7411, w_eco7412, w_eco7413, w_eco7414, w_eco7415, w_eco7416, w_eco7417, w_eco7418, w_eco7419, w_eco7420, w_eco7421, w_eco7422, w_eco7423, w_eco7424, w_eco7425, w_eco7426, w_eco7427, w_eco7428, w_eco7429, w_eco7430, w_eco7431, w_eco7432, w_eco7433, w_eco7434, w_eco7435, w_eco7436, w_eco7437, w_eco7438, w_eco7439, w_eco7440, w_eco7441, w_eco7442, w_eco7443, w_eco7444, w_eco7445, w_eco7446, w_eco7447, w_eco7448, w_eco7449, w_eco7450, w_eco7451, w_eco7452, w_eco7453, w_eco7454, w_eco7455, w_eco7456, w_eco7457, w_eco7458, w_eco7459, w_eco7460, w_eco7461, w_eco7462, w_eco7463, w_eco7464, w_eco7465, w_eco7466, w_eco7467, w_eco7468, w_eco7469, w_eco7470, w_eco7471, w_eco7472, w_eco7473, w_eco7474, w_eco7475, w_eco7476, w_eco7477, w_eco7478, w_eco7479, w_eco7480, w_eco7481, w_eco7482, w_eco7483, w_eco7484, w_eco7485, w_eco7486, w_eco7487, w_eco7488, w_eco7489, w_eco7490, w_eco7491, w_eco7492, w_eco7493, w_eco7494, w_eco7495, w_eco7496, w_eco7497, w_eco7498, w_eco7499, w_eco7500, w_eco7501, w_eco7502, w_eco7503, w_eco7504, w_eco7505, w_eco7506, w_eco7507, w_eco7508, w_eco7509, w_eco7510, w_eco7511, w_eco7512, w_eco7513, w_eco7514, w_eco7515, w_eco7516, w_eco7517, w_eco7518, w_eco7519, w_eco7520, w_eco7521, w_eco7522, w_eco7523, w_eco7524, w_eco7525, w_eco7526, w_eco7527, w_eco7528, w_eco7529, w_eco7530, w_eco7531, w_eco7532, w_eco7533, w_eco7534, w_eco7535, w_eco7536, w_eco7537, w_eco7538, w_eco7539, w_eco7540, w_eco7541, w_eco7542, w_eco7543, w_eco7544, w_eco7545, w_eco7546, w_eco7547, w_eco7548, w_eco7549, w_eco7550, w_eco7551, w_eco7552, w_eco7553, w_eco7554, w_eco7555, w_eco7556, w_eco7557, w_eco7558, w_eco7559, w_eco7560, w_eco7561, w_eco7562, w_eco7563, w_eco7564, w_eco7565, w_eco7566, w_eco7567, w_eco7568, w_eco7569, w_eco7570, w_eco7571, w_eco7572, w_eco7573, w_eco7574, w_eco7575, w_eco7576, w_eco7577, w_eco7578, w_eco7579, w_eco7580, w_eco7581, w_eco7582, w_eco7583, w_eco7584, w_eco7585, w_eco7586, w_eco7587, w_eco7588, w_eco7589, w_eco7590, w_eco7591, w_eco7592, w_eco7593, w_eco7594, w_eco7595, w_eco7596, w_eco7597, w_eco7598, w_eco7599, w_eco7600, w_eco7601, w_eco7602, w_eco7603, w_eco7604, w_eco7605, w_eco7606, w_eco7607, w_eco7608, w_eco7609, w_eco7610, w_eco7611, w_eco7612, w_eco7613, w_eco7614, w_eco7615, w_eco7616, w_eco7617, w_eco7618, w_eco7619, w_eco7620, w_eco7621, w_eco7622, w_eco7623, w_eco7624, w_eco7625, w_eco7626, w_eco7627, w_eco7628, w_eco7629, w_eco7630, w_eco7631, w_eco7632, w_eco7633, w_eco7634, w_eco7635, w_eco7636, w_eco7637, w_eco7638, w_eco7639, w_eco7640, w_eco7641, w_eco7642, w_eco7643, w_eco7644, w_eco7645, w_eco7646, w_eco7647, w_eco7648, w_eco7649, w_eco7650, w_eco7651, w_eco7652, w_eco7653, w_eco7654, w_eco7655, w_eco7656, w_eco7657, w_eco7658, w_eco7659, w_eco7660, w_eco7661, w_eco7662, w_eco7663, w_eco7664, w_eco7665, w_eco7666, w_eco7667, w_eco7668, w_eco7669, w_eco7670, w_eco7671, w_eco7672, w_eco7673, w_eco7674, w_eco7675, w_eco7676, w_eco7677, w_eco7678, w_eco7679, w_eco7680, w_eco7681, w_eco7682, w_eco7683, w_eco7684, w_eco7685, w_eco7686, w_eco7687, w_eco7688, w_eco7689, w_eco7690, w_eco7691, w_eco7692, w_eco7693, w_eco7694, w_eco7695, w_eco7696, w_eco7697, w_eco7698, w_eco7699, w_eco7700, w_eco7701, w_eco7702, w_eco7703, w_eco7704, w_eco7705, w_eco7706, w_eco7707, w_eco7708, w_eco7709, w_eco7710, w_eco7711, w_eco7712, w_eco7713, w_eco7714, w_eco7715, w_eco7716, w_eco7717, w_eco7718, w_eco7719, w_eco7720, w_eco7721, w_eco7722, w_eco7723, w_eco7724, w_eco7725, w_eco7726, w_eco7727, w_eco7728, w_eco7729, w_eco7730, w_eco7731, w_eco7732, w_eco7733, w_eco7734, w_eco7735, w_eco7736, w_eco7737, w_eco7738, w_eco7739, w_eco7740, w_eco7741, w_eco7742, w_eco7743, w_eco7744, w_eco7745, w_eco7746, w_eco7747, w_eco7748, w_eco7749, w_eco7750, w_eco7751, w_eco7752, w_eco7753, w_eco7754, w_eco7755, w_eco7756, w_eco7757, w_eco7758, w_eco7759, w_eco7760, w_eco7761, w_eco7762, w_eco7763, w_eco7764, w_eco7765, w_eco7766, w_eco7767, w_eco7768, w_eco7769, w_eco7770, w_eco7771, w_eco7772, w_eco7773, w_eco7774, w_eco7775, w_eco7776, w_eco7777, w_eco7778, w_eco7779, w_eco7780, w_eco7781, w_eco7782, w_eco7783, w_eco7784, w_eco7785, w_eco7786, w_eco7787, w_eco7788, w_eco7789, w_eco7790, w_eco7791, w_eco7792, w_eco7793, w_eco7794, w_eco7795, w_eco7796, w_eco7797, w_eco7798, w_eco7799, sub_wire6, w_eco7800, w_eco7801, w_eco7802, w_eco7803, w_eco7804, w_eco7805, w_eco7806, w_eco7807, w_eco7808, w_eco7809, w_eco7810, w_eco7811, w_eco7812, w_eco7813, w_eco7814, w_eco7815, w_eco7816, w_eco7817, w_eco7818, w_eco7819, w_eco7820, w_eco7821, w_eco7822, w_eco7823, w_eco7824, w_eco7825, w_eco7826, w_eco7827, w_eco7828, w_eco7829, w_eco7830, w_eco7831, w_eco7832, w_eco7833, w_eco7834, w_eco7835, w_eco7836, w_eco7837, w_eco7838, w_eco7839, w_eco7840, w_eco7841, w_eco7842, w_eco7843, w_eco7844, w_eco7845, w_eco7846, w_eco7847, w_eco7848, w_eco7849, w_eco7850, w_eco7851, w_eco7852, w_eco7853, w_eco7854, w_eco7855, w_eco7856, w_eco7857, w_eco7858, w_eco7859, w_eco7860, w_eco7861, w_eco7862, w_eco7863, w_eco7864, w_eco7865, w_eco7866, w_eco7867, w_eco7868, w_eco7869, w_eco7870, w_eco7871, w_eco7872, w_eco7873, w_eco7874, w_eco7875, w_eco7876, w_eco7877, w_eco7878, w_eco7879, w_eco7880, w_eco7881, w_eco7882, w_eco7883, w_eco7884, w_eco7885, w_eco7886, w_eco7887, w_eco7888, w_eco7889, w_eco7890, w_eco7891, w_eco7892, w_eco7893, w_eco7894, w_eco7895, w_eco7896, w_eco7897, w_eco7898, w_eco7899, w_eco7900, w_eco7901, w_eco7902, w_eco7903, w_eco7904, w_eco7905, w_eco7906, w_eco7907, w_eco7908, w_eco7909, w_eco7910, w_eco7911, w_eco7912, w_eco7913, w_eco7914, w_eco7915, w_eco7916, w_eco7917, w_eco7918, w_eco7919, w_eco7920, w_eco7921, w_eco7922, w_eco7923, w_eco7924, w_eco7925, w_eco7926, w_eco7927, w_eco7928, w_eco7929, w_eco7930, w_eco7931, w_eco7932, w_eco7933, w_eco7934, w_eco7935, w_eco7936, w_eco7937, w_eco7938, w_eco7939, w_eco7940, w_eco7941, w_eco7942, w_eco7943, w_eco7944, w_eco7945, w_eco7946, w_eco7947, w_eco7948, w_eco7949, w_eco7950, w_eco7951, w_eco7952, w_eco7953, w_eco7954, w_eco7955, w_eco7956, w_eco7957, w_eco7958, w_eco7959, w_eco7960, w_eco7961, w_eco7962, w_eco7963, w_eco7964, w_eco7965, w_eco7966, w_eco7967, w_eco7968, w_eco7969, w_eco7970, w_eco7971, w_eco7972, w_eco7973, w_eco7974, w_eco7975, w_eco7976, w_eco7977, w_eco7978, w_eco7979, w_eco7980, w_eco7981, w_eco7982, w_eco7983, w_eco7984, w_eco7985, w_eco7986, w_eco7987, w_eco7988, w_eco7989, w_eco7990, w_eco7991, w_eco7992, w_eco7993, w_eco7994, w_eco7995, w_eco7996, w_eco7997, w_eco7998, w_eco7999, w_eco8000, w_eco8001, w_eco8002, w_eco8003, w_eco8004, w_eco8005, w_eco8006, w_eco8007, w_eco8008, w_eco8009, w_eco8010, w_eco8011, w_eco8012, w_eco8013, w_eco8014, w_eco8015, w_eco8016, w_eco8017, w_eco8018, w_eco8019, w_eco8020, w_eco8021, w_eco8022, w_eco8023, w_eco8024, w_eco8025, w_eco8026, w_eco8027, w_eco8028, w_eco8029, w_eco8030, w_eco8031, w_eco8032, w_eco8033, w_eco8034, w_eco8035, w_eco8036, w_eco8037, w_eco8038, w_eco8039, w_eco8040, w_eco8041, w_eco8042, w_eco8043, w_eco8044, w_eco8045, w_eco8046, w_eco8047, w_eco8048, w_eco8049, w_eco8050, w_eco8051, w_eco8052, w_eco8053, w_eco8054, w_eco8055, w_eco8056, w_eco8057, w_eco8058, w_eco8059, w_eco8060, w_eco8061, w_eco8062, w_eco8063, w_eco8064, w_eco8065, w_eco8066, w_eco8067, w_eco8068, w_eco8069, w_eco8070, w_eco8071, w_eco8072, w_eco8073, w_eco8074, w_eco8075, w_eco8076, w_eco8077, w_eco8078, w_eco8079, w_eco8080, w_eco8081, w_eco8082, w_eco8083, w_eco8084, w_eco8085, w_eco8086, w_eco8087, w_eco8088, w_eco8089, w_eco8090, w_eco8091, w_eco8092, w_eco8093, w_eco8094, w_eco8095, w_eco8096, w_eco8097, w_eco8098, w_eco8099, w_eco8100, w_eco8101, w_eco8102, w_eco8103, w_eco8104, w_eco8105, w_eco8106, w_eco8107, w_eco8108, w_eco8109, w_eco8110, w_eco8111, w_eco8112, w_eco8113, w_eco8114, w_eco8115, w_eco8116, w_eco8117, w_eco8118, w_eco8119, w_eco8120, w_eco8121, w_eco8122, w_eco8123, w_eco8124, w_eco8125, w_eco8126, w_eco8127, w_eco8128, w_eco8129, w_eco8130, w_eco8131, w_eco8132, w_eco8133, w_eco8134, w_eco8135, w_eco8136, w_eco8137, w_eco8138, w_eco8139, w_eco8140, w_eco8141, w_eco8142, w_eco8143, w_eco8144, w_eco8145, w_eco8146, w_eco8147, w_eco8148, w_eco8149, w_eco8150, w_eco8151, w_eco8152, w_eco8153, w_eco8154, w_eco8155, w_eco8156, w_eco8157, w_eco8158, w_eco8159, w_eco8160, w_eco8161, w_eco8162, w_eco8163, w_eco8164, w_eco8165, w_eco8166, w_eco8167, w_eco8168, w_eco8169, w_eco8170, w_eco8171, w_eco8172, w_eco8173, w_eco8174, w_eco8175, w_eco8176, w_eco8177, w_eco8178, w_eco8179, w_eco8180, w_eco8181, w_eco8182, w_eco8183, w_eco8184, w_eco8185, w_eco8186, w_eco8187, w_eco8188, w_eco8189, w_eco8190, w_eco8191, w_eco8192, w_eco8193, w_eco8194, w_eco8195, w_eco8196, w_eco8197, w_eco8198, w_eco8199, w_eco8200, w_eco8201, w_eco8202, w_eco8203, w_eco8204, w_eco8205, w_eco8206, w_eco8207, w_eco8208, w_eco8209, w_eco8210, w_eco8211, w_eco8212, w_eco8213, w_eco8214, w_eco8215, w_eco8216, w_eco8217, w_eco8218, w_eco8219, w_eco8220, w_eco8221, w_eco8222, w_eco8223, w_eco8224, w_eco8225, w_eco8226, w_eco8227, w_eco8228, w_eco8229, w_eco8230, w_eco8231, w_eco8232, w_eco8233, w_eco8234, w_eco8235, w_eco8236, w_eco8237, w_eco8238, w_eco8239, w_eco8240, w_eco8241, w_eco8242, w_eco8243, w_eco8244, w_eco8245, w_eco8246, w_eco8247, w_eco8248, w_eco8249, w_eco8250, w_eco8251, w_eco8252, w_eco8253, w_eco8254, w_eco8255, w_eco8256, w_eco8257, w_eco8258, w_eco8259, w_eco8260, w_eco8261, w_eco8262, w_eco8263, w_eco8264, w_eco8265, w_eco8266, w_eco8267, w_eco8268, w_eco8269, w_eco8270, w_eco8271, w_eco8272, w_eco8273, w_eco8274, w_eco8275, w_eco8276, w_eco8277, w_eco8278, w_eco8279, w_eco8280, w_eco8281, w_eco8282, w_eco8283, w_eco8284, w_eco8285, w_eco8286, w_eco8287, w_eco8288, w_eco8289, w_eco8290, w_eco8291, w_eco8292, w_eco8293, w_eco8294, w_eco8295, w_eco8296, w_eco8297, w_eco8298, w_eco8299, w_eco8300, w_eco8301, w_eco8302, w_eco8303, w_eco8304, w_eco8305, w_eco8306, w_eco8307, w_eco8308, w_eco8309, w_eco8310, w_eco8311, w_eco8312, w_eco8313, w_eco8314, w_eco8315, w_eco8316, w_eco8317, w_eco8318, w_eco8319, w_eco8320, w_eco8321, w_eco8322, w_eco8323, w_eco8324, w_eco8325, w_eco8326, w_eco8327, w_eco8328, w_eco8329, w_eco8330, w_eco8331, w_eco8332, w_eco8333, w_eco8334, w_eco8335, w_eco8336, w_eco8337, w_eco8338, w_eco8339, w_eco8340, w_eco8341, w_eco8342, w_eco8343, w_eco8344, w_eco8345, w_eco8346, w_eco8347, w_eco8348, w_eco8349, w_eco8350, w_eco8351, w_eco8352, w_eco8353, w_eco8354, w_eco8355, w_eco8356, w_eco8357, w_eco8358, w_eco8359, w_eco8360, w_eco8361, w_eco8362, w_eco8363, w_eco8364, w_eco8365, w_eco8366, w_eco8367, w_eco8368, w_eco8369, w_eco8370, w_eco8371, w_eco8372, w_eco8373, w_eco8374, w_eco8375, w_eco8376, w_eco8377, w_eco8378, w_eco8379, w_eco8380, w_eco8381, w_eco8382, w_eco8383, w_eco8384, w_eco8385, w_eco8386, w_eco8387, w_eco8388, w_eco8389, w_eco8390, w_eco8391, w_eco8392, w_eco8393, w_eco8394, w_eco8395, w_eco8396, w_eco8397, w_eco8398, w_eco8399, w_eco8400, w_eco8401, w_eco8402, w_eco8403, w_eco8404, w_eco8405, w_eco8406, w_eco8407, w_eco8408, w_eco8409, w_eco8410, w_eco8411, w_eco8412, w_eco8413, w_eco8414, w_eco8415, w_eco8416, w_eco8417, w_eco8418, w_eco8419, w_eco8420, w_eco8421, w_eco8422, w_eco8423, w_eco8424, w_eco8425, w_eco8426, w_eco8427, w_eco8428, w_eco8429, w_eco8430, w_eco8431, w_eco8432, w_eco8433, w_eco8434, w_eco8435, w_eco8436, w_eco8437, w_eco8438, w_eco8439, w_eco8440, w_eco8441, w_eco8442, w_eco8443, w_eco8444, w_eco8445, w_eco8446, w_eco8447, w_eco8448, w_eco8449, w_eco8450, w_eco8451, w_eco8452, w_eco8453, w_eco8454, w_eco8455, w_eco8456, w_eco8457, w_eco8458, w_eco8459, w_eco8460, w_eco8461, w_eco8462, w_eco8463, w_eco8464, w_eco8465, w_eco8466, w_eco8467, w_eco8468, w_eco8469, w_eco8470, w_eco8471, w_eco8472, w_eco8473, w_eco8474, w_eco8475, w_eco8476, w_eco8477, w_eco8478, w_eco8479, w_eco8480, w_eco8481, w_eco8482, w_eco8483, w_eco8484, w_eco8485, w_eco8486, w_eco8487, w_eco8488, w_eco8489, w_eco8490, w_eco8491, w_eco8492, w_eco8493, w_eco8494, w_eco8495, w_eco8496, w_eco8497, w_eco8498, w_eco8499, w_eco8500, w_eco8501, w_eco8502, w_eco8503, w_eco8504, w_eco8505, w_eco8506, w_eco8507, w_eco8508, w_eco8509, w_eco8510, w_eco8511, w_eco8512, w_eco8513, w_eco8514, w_eco8515, w_eco8516, w_eco8517, w_eco8518, w_eco8519, w_eco8520, w_eco8521, w_eco8522, w_eco8523, w_eco8524, w_eco8525, w_eco8526, w_eco8527, w_eco8528, w_eco8529, w_eco8530, w_eco8531, w_eco8532, w_eco8533, w_eco8534, w_eco8535, w_eco8536, w_eco8537, w_eco8538, w_eco8539, w_eco8540, w_eco8541, w_eco8542, w_eco8543, w_eco8544, w_eco8545, w_eco8546, w_eco8547, w_eco8548, w_eco8549, w_eco8550, w_eco8551, w_eco8552, w_eco8553, w_eco8554, w_eco8555, w_eco8556, w_eco8557, w_eco8558, w_eco8559, w_eco8560, w_eco8561, w_eco8562, w_eco8563, w_eco8564, w_eco8565, w_eco8566, w_eco8567, w_eco8568, w_eco8569, w_eco8570, w_eco8571, w_eco8572, w_eco8573, w_eco8574, w_eco8575, w_eco8576, w_eco8577, w_eco8578, w_eco8579, w_eco8580, w_eco8581, w_eco8582, w_eco8583, w_eco8584, w_eco8585, w_eco8586, w_eco8587, w_eco8588, w_eco8589, w_eco8590, w_eco8591, w_eco8592, w_eco8593, w_eco8594, w_eco8595, w_eco8596, w_eco8597, w_eco8598, w_eco8599, w_eco8600, w_eco8601, w_eco8602, w_eco8603, w_eco8604, w_eco8605, w_eco8606, w_eco8607, w_eco8608, w_eco8609, w_eco8610, w_eco8611, w_eco8612, w_eco8613, w_eco8614, w_eco8615, w_eco8616, w_eco8617, w_eco8618, w_eco8619, w_eco8620, w_eco8621, w_eco8622, w_eco8623, w_eco8624, w_eco8625, w_eco8626, w_eco8627, w_eco8628, w_eco8629, w_eco8630, w_eco8631, w_eco8632, w_eco8633, w_eco8634, w_eco8635, w_eco8636, w_eco8637, w_eco8638, w_eco8639, w_eco8640, w_eco8641, w_eco8642, w_eco8643, w_eco8644, w_eco8645, w_eco8646, w_eco8647, w_eco8648, w_eco8649, w_eco8650, w_eco8651, w_eco8652, w_eco8653, w_eco8654, w_eco8655, w_eco8656, w_eco8657, w_eco8658, w_eco8659, w_eco8660, w_eco8661, w_eco8662, w_eco8663, w_eco8664, w_eco8665, w_eco8666, w_eco8667, w_eco8668, w_eco8669, w_eco8670, w_eco8671, w_eco8672, w_eco8673, w_eco8674, w_eco8675, w_eco8676, w_eco8677, w_eco8678, w_eco8679, w_eco8680, w_eco8681, w_eco8682, w_eco8683, w_eco8684, w_eco8685, w_eco8686, w_eco8687, w_eco8688, w_eco8689, w_eco8690, w_eco8691, w_eco8692, w_eco8693, w_eco8694, w_eco8695, w_eco8696, w_eco8697, w_eco8698, w_eco8699, w_eco8700, w_eco8701, w_eco8702, w_eco8703, w_eco8704, w_eco8705, w_eco8706, w_eco8707, w_eco8708, w_eco8709, w_eco8710, w_eco8711, w_eco8712, w_eco8713, w_eco8714, w_eco8715, w_eco8716, w_eco8717, w_eco8718, w_eco8719, w_eco8720, w_eco8721, w_eco8722, w_eco8723, w_eco8724, w_eco8725, w_eco8726, w_eco8727, w_eco8728, w_eco8729, w_eco8730, w_eco8731, w_eco8732, w_eco8733, w_eco8734, w_eco8735, w_eco8736, w_eco8737, w_eco8738, w_eco8739, w_eco8740, w_eco8741, w_eco8742, w_eco8743, w_eco8744, w_eco8745, w_eco8746, w_eco8747, w_eco8748, w_eco8749, w_eco8750, w_eco8751, w_eco8752, w_eco8753, w_eco8754, w_eco8755, w_eco8756, w_eco8757, w_eco8758, w_eco8759, w_eco8760, w_eco8761, w_eco8762, w_eco8763, w_eco8764, w_eco8765, w_eco8766, w_eco8767, w_eco8768, w_eco8769, w_eco8770, w_eco8771, w_eco8772, w_eco8773, w_eco8774, w_eco8775, w_eco8776, w_eco8777, w_eco8778, w_eco8779, w_eco8780, w_eco8781, w_eco8782, w_eco8783, w_eco8784, w_eco8785, w_eco8786, w_eco8787, w_eco8788, w_eco8789, w_eco8790, w_eco8791, w_eco8792, w_eco8793, w_eco8794, w_eco8795, w_eco8796, w_eco8797, w_eco8798, w_eco8799, w_eco8800, w_eco8801, w_eco8802, w_eco8803, w_eco8804, w_eco8805, w_eco8806, w_eco8807, w_eco8808, w_eco8809, w_eco8810, w_eco8811, w_eco8812, w_eco8813, w_eco8814, w_eco8815, w_eco8816, w_eco8817, w_eco8818, w_eco8819, w_eco8820, w_eco8821, w_eco8822, w_eco8823, w_eco8824, w_eco8825, w_eco8826, w_eco8827, w_eco8828, w_eco8829, w_eco8830, w_eco8831, w_eco8832, w_eco8833, w_eco8834, w_eco8835, w_eco8836, w_eco8837, w_eco8838, w_eco8839, w_eco8840, w_eco8841, w_eco8842, w_eco8843, w_eco8844, w_eco8845, w_eco8846, w_eco8847, w_eco8848, w_eco8849, w_eco8850, w_eco8851, w_eco8852, w_eco8853, w_eco8854, w_eco8855, w_eco8856, w_eco8857, w_eco8858, w_eco8859, w_eco8860, w_eco8861, w_eco8862, w_eco8863, w_eco8864, w_eco8865, w_eco8866, w_eco8867, w_eco8868, w_eco8869, w_eco8870, w_eco8871, w_eco8872, w_eco8873, w_eco8874, w_eco8875, w_eco8876, w_eco8877, w_eco8878, w_eco8879, w_eco8880, w_eco8881, w_eco8882, w_eco8883, w_eco8884, w_eco8885, w_eco8886, w_eco8887, w_eco8888, w_eco8889, w_eco8890, w_eco8891, w_eco8892, w_eco8893, w_eco8894, w_eco8895, w_eco8896, w_eco8897, w_eco8898, w_eco8899, w_eco8900, w_eco8901, w_eco8902, w_eco8903, w_eco8904, w_eco8905, w_eco8906, w_eco8907, w_eco8908, w_eco8909, w_eco8910, w_eco8911, w_eco8912, w_eco8913, w_eco8914, w_eco8915, w_eco8916, w_eco8917, w_eco8918, w_eco8919, w_eco8920, w_eco8921, w_eco8922, w_eco8923, w_eco8924, w_eco8925, w_eco8926, w_eco8927, w_eco8928, w_eco8929, w_eco8930, w_eco8931, w_eco8932, w_eco8933, w_eco8934, w_eco8935, w_eco8936, w_eco8937, w_eco8938, w_eco8939, w_eco8940, w_eco8941, w_eco8942, w_eco8943, w_eco8944, w_eco8945, w_eco8946, w_eco8947, w_eco8948, w_eco8949, w_eco8950, w_eco8951, w_eco8952, w_eco8953, w_eco8954, w_eco8955, w_eco8956, w_eco8957, w_eco8958, w_eco8959, w_eco8960, w_eco8961, w_eco8962, w_eco8963, w_eco8964, w_eco8965, w_eco8966, w_eco8967, w_eco8968, w_eco8969, w_eco8970, w_eco8971, w_eco8972, w_eco8973, w_eco8974, w_eco8975, w_eco8976, w_eco8977, w_eco8978, w_eco8979, w_eco8980, w_eco8981, w_eco8982, w_eco8983, w_eco8984, w_eco8985, w_eco8986, w_eco8987, w_eco8988, w_eco8989, w_eco8990, w_eco8991, w_eco8992, w_eco8993, w_eco8994, w_eco8995, w_eco8996, w_eco8997, w_eco8998, w_eco8999, w_eco9000, w_eco9001, w_eco9002, w_eco9003, w_eco9004, w_eco9005, w_eco9006, w_eco9007, w_eco9008, w_eco9009, w_eco9010, w_eco9011, w_eco9012, w_eco9013, w_eco9014, w_eco9015, w_eco9016, w_eco9017, w_eco9018, w_eco9019, w_eco9020, w_eco9021, w_eco9022, w_eco9023, w_eco9024, w_eco9025, w_eco9026, w_eco9027, w_eco9028, w_eco9029, w_eco9030, w_eco9031, w_eco9032, w_eco9033, w_eco9034, w_eco9035, w_eco9036, w_eco9037, w_eco9038, w_eco9039, w_eco9040, w_eco9041, w_eco9042, w_eco9043, w_eco9044, w_eco9045, w_eco9046, w_eco9047, w_eco9048, w_eco9049, w_eco9050, w_eco9051, w_eco9052, w_eco9053, w_eco9054, w_eco9055, w_eco9056, w_eco9057, w_eco9058, w_eco9059, w_eco9060, w_eco9061, w_eco9062, w_eco9063, w_eco9064, w_eco9065, w_eco9066, w_eco9067, w_eco9068, w_eco9069, w_eco9070, w_eco9071, w_eco9072, w_eco9073, w_eco9074, w_eco9075, w_eco9076, w_eco9077, w_eco9078, w_eco9079, w_eco9080, w_eco9081, w_eco9082, w_eco9083, w_eco9084, w_eco9085, w_eco9086, w_eco9087, w_eco9088, w_eco9089, w_eco9090, w_eco9091, w_eco9092, w_eco9093, w_eco9094, w_eco9095, w_eco9096, w_eco9097, w_eco9098, w_eco9099, w_eco9100, w_eco9101, w_eco9102, w_eco9103, w_eco9104, w_eco9105, w_eco9106, w_eco9107, w_eco9108, w_eco9109, w_eco9110, w_eco9111, w_eco9112, w_eco9113, w_eco9114, w_eco9115, w_eco9116, w_eco9117, w_eco9118, w_eco9119, w_eco9120, w_eco9121, w_eco9122, w_eco9123, w_eco9124, w_eco9125, w_eco9126, w_eco9127, w_eco9128, w_eco9129, w_eco9130, w_eco9131, w_eco9132, w_eco9133, w_eco9134, w_eco9135, w_eco9136, w_eco9137, w_eco9138, w_eco9139, w_eco9140, w_eco9141, w_eco9142, w_eco9143, w_eco9144, w_eco9145, w_eco9146, w_eco9147, w_eco9148, w_eco9149, w_eco9150, w_eco9151, w_eco9152, w_eco9153, w_eco9154, w_eco9155, w_eco9156, w_eco9157, w_eco9158, w_eco9159, w_eco9160, w_eco9161, w_eco9162, w_eco9163, w_eco9164, w_eco9165, w_eco9166, w_eco9167, w_eco9168, w_eco9169, w_eco9170, w_eco9171, w_eco9172, w_eco9173, w_eco9174, w_eco9175, w_eco9176, w_eco9177, w_eco9178, w_eco9179, w_eco9180, w_eco9181, w_eco9182, w_eco9183, w_eco9184, w_eco9185, w_eco9186, w_eco9187, w_eco9188, w_eco9189, w_eco9190, w_eco9191, w_eco9192, w_eco9193, w_eco9194, w_eco9195, w_eco9196, w_eco9197, w_eco9198, w_eco9199, w_eco9200, w_eco9201, w_eco9202, w_eco9203, w_eco9204, w_eco9205, w_eco9206, w_eco9207, w_eco9208, w_eco9209, w_eco9210, w_eco9211, w_eco9212, w_eco9213, w_eco9214, w_eco9215, w_eco9216, w_eco9217, w_eco9218, w_eco9219, w_eco9220, w_eco9221, w_eco9222, w_eco9223, w_eco9224, w_eco9225, w_eco9226, w_eco9227, w_eco9228, w_eco9229, w_eco9230, w_eco9231, w_eco9232, w_eco9233, w_eco9234, w_eco9235, w_eco9236, w_eco9237, w_eco9238, w_eco9239, w_eco9240, w_eco9241, w_eco9242, w_eco9243, w_eco9244, w_eco9245, w_eco9246, w_eco9247, w_eco9248, w_eco9249, w_eco9250, w_eco9251, w_eco9252, w_eco9253, w_eco9254, w_eco9255, w_eco9256, w_eco9257, w_eco9258, w_eco9259, w_eco9260, w_eco9261, w_eco9262, w_eco9263, w_eco9264, w_eco9265, w_eco9266, w_eco9267, w_eco9268, w_eco9269, w_eco9270, w_eco9271, w_eco9272, w_eco9273, w_eco9274, w_eco9275, w_eco9276, w_eco9277, w_eco9278, w_eco9279, w_eco9280, w_eco9281, w_eco9282, w_eco9283, w_eco9284, w_eco9285, w_eco9286, w_eco9287, w_eco9288, w_eco9289, w_eco9290, w_eco9291, w_eco9292, w_eco9293, w_eco9294, w_eco9295, w_eco9296, w_eco9297, w_eco9298, w_eco9299, w_eco9300, w_eco9301, w_eco9302, w_eco9303, w_eco9304, w_eco9305, w_eco9306, w_eco9307, w_eco9308, w_eco9309, w_eco9310, w_eco9311, w_eco9312, w_eco9313, w_eco9314, w_eco9315, w_eco9316, w_eco9317, w_eco9318, w_eco9319, w_eco9320, w_eco9321, w_eco9322, w_eco9323, w_eco9324, w_eco9325, w_eco9326, w_eco9327, w_eco9328, w_eco9329, w_eco9330, w_eco9331, w_eco9332, w_eco9333, w_eco9334, w_eco9335, w_eco9336, w_eco9337, w_eco9338, w_eco9339, w_eco9340, w_eco9341, w_eco9342, w_eco9343, w_eco9344, w_eco9345, w_eco9346, w_eco9347, w_eco9348, w_eco9349, w_eco9350, w_eco9351, w_eco9352, w_eco9353, w_eco9354, w_eco9355, w_eco9356, w_eco9357, w_eco9358, w_eco9359, w_eco9360, w_eco9361, w_eco9362, w_eco9363, w_eco9364, w_eco9365, w_eco9366, w_eco9367, w_eco9368, w_eco9369, w_eco9370, w_eco9371, w_eco9372, w_eco9373, w_eco9374, w_eco9375, w_eco9376, w_eco9377, w_eco9378, w_eco9379, w_eco9380, w_eco9381, w_eco9382, w_eco9383, w_eco9384, w_eco9385, w_eco9386, w_eco9387, w_eco9388, w_eco9389, w_eco9390, w_eco9391, w_eco9392, w_eco9393, w_eco9394, w_eco9395, w_eco9396, w_eco9397, w_eco9398, w_eco9399, w_eco9400, w_eco9401, w_eco9402, w_eco9403, w_eco9404, w_eco9405, w_eco9406, w_eco9407, w_eco9408, w_eco9409, w_eco9410, w_eco9411, w_eco9412, w_eco9413, w_eco9414, w_eco9415, w_eco9416, w_eco9417, w_eco9418, w_eco9419, w_eco9420, w_eco9421, w_eco9422, w_eco9423, w_eco9424, w_eco9425, w_eco9426, w_eco9427, w_eco9428, w_eco9429, w_eco9430, w_eco9431, w_eco9432, w_eco9433, w_eco9434, w_eco9435, w_eco9436, w_eco9437, w_eco9438, w_eco9439, w_eco9440, w_eco9441, w_eco9442, w_eco9443, w_eco9444, w_eco9445, w_eco9446, w_eco9447, w_eco9448, w_eco9449, w_eco9450, w_eco9451, w_eco9452, w_eco9453, w_eco9454, w_eco9455, w_eco9456, w_eco9457, w_eco9458, w_eco9459, w_eco9460, w_eco9461, w_eco9462, w_eco9463, w_eco9464, w_eco9465, w_eco9466, w_eco9467, w_eco9468, w_eco9469, w_eco9470, w_eco9471, w_eco9472, w_eco9473, w_eco9474, w_eco9475, w_eco9476, w_eco9477, w_eco9478, w_eco9479, w_eco9480, w_eco9481, w_eco9482, w_eco9483, w_eco9484, w_eco9485, w_eco9486, w_eco9487, w_eco9488, w_eco9489, w_eco9490, w_eco9491, w_eco9492, w_eco9493, w_eco9494, w_eco9495, w_eco9496, w_eco9497, w_eco9498, w_eco9499, w_eco9500, w_eco9501, w_eco9502, w_eco9503, w_eco9504, w_eco9505, w_eco9506, w_eco9507, w_eco9508, w_eco9509, w_eco9510, w_eco9511, w_eco9512, w_eco9513, w_eco9514, w_eco9515, w_eco9516, w_eco9517, w_eco9518, w_eco9519, w_eco9520, w_eco9521, w_eco9522, w_eco9523, w_eco9524, w_eco9525, w_eco9526, w_eco9527, w_eco9528, w_eco9529, w_eco9530, w_eco9531, w_eco9532, w_eco9533, w_eco9534, w_eco9535, w_eco9536, w_eco9537, w_eco9538, w_eco9539, w_eco9540, w_eco9541, w_eco9542, w_eco9543, w_eco9544, w_eco9545, w_eco9546, w_eco9547, w_eco9548, w_eco9549, w_eco9550, w_eco9551, w_eco9552, w_eco9553, w_eco9554, w_eco9555, w_eco9556, w_eco9557, w_eco9558, w_eco9559, w_eco9560, w_eco9561, w_eco9562, w_eco9563, w_eco9564, w_eco9565, w_eco9566, w_eco9567, w_eco9568, w_eco9569, w_eco9570, w_eco9571, w_eco9572, w_eco9573, w_eco9574, w_eco9575, w_eco9576, w_eco9577, w_eco9578, w_eco9579, w_eco9580, w_eco9581, w_eco9582, w_eco9583, w_eco9584, w_eco9585, sub_wire7, w_eco9586, w_eco9587, w_eco9588, w_eco9589, w_eco9590, w_eco9591, w_eco9592, w_eco9593, w_eco9594, w_eco9595, w_eco9596, w_eco9597, w_eco9598, w_eco9599, w_eco9600, w_eco9601, w_eco9602, w_eco9603, w_eco9604, w_eco9605, w_eco9606, w_eco9607, w_eco9608, w_eco9609, w_eco9610, w_eco9611, w_eco9612, w_eco9613, w_eco9614, w_eco9615, w_eco9616, w_eco9617, w_eco9618, w_eco9619, w_eco9620, w_eco9621, w_eco9622, w_eco9623, w_eco9624, w_eco9625, w_eco9626, w_eco9627, w_eco9628, w_eco9629, w_eco9630, w_eco9631, w_eco9632, w_eco9633, w_eco9634, w_eco9635, w_eco9636, w_eco9637, w_eco9638, w_eco9639, w_eco9640, w_eco9641, w_eco9642, w_eco9643, w_eco9644, w_eco9645, w_eco9646, w_eco9647, w_eco9648, w_eco9649, w_eco9650, w_eco9651, w_eco9652, w_eco9653, w_eco9654, w_eco9655, w_eco9656, w_eco9657, w_eco9658, w_eco9659, w_eco9660, w_eco9661, w_eco9662, w_eco9663, w_eco9664, w_eco9665, w_eco9666, w_eco9667, w_eco9668, w_eco9669, w_eco9670, w_eco9671, w_eco9672, w_eco9673, w_eco9674, w_eco9675, w_eco9676, w_eco9677, w_eco9678, w_eco9679, w_eco9680, w_eco9681, w_eco9682, w_eco9683, w_eco9684, w_eco9685, w_eco9686, w_eco9687, w_eco9688, w_eco9689, w_eco9690, w_eco9691, w_eco9692, w_eco9693, w_eco9694, w_eco9695, w_eco9696, w_eco9697, w_eco9698, w_eco9699, w_eco9700, w_eco9701, w_eco9702, w_eco9703, w_eco9704, w_eco9705, w_eco9706, w_eco9707, w_eco9708, w_eco9709, w_eco9710, w_eco9711, w_eco9712, w_eco9713, w_eco9714, w_eco9715, w_eco9716, w_eco9717, w_eco9718, w_eco9719, w_eco9720, w_eco9721, w_eco9722, w_eco9723, w_eco9724, w_eco9725, w_eco9726, w_eco9727, w_eco9728, w_eco9729, w_eco9730, w_eco9731, w_eco9732, w_eco9733, w_eco9734, w_eco9735, w_eco9736, w_eco9737, w_eco9738, w_eco9739, w_eco9740, w_eco9741, w_eco9742, w_eco9743, w_eco9744, w_eco9745, w_eco9746, w_eco9747, w_eco9748, w_eco9749, w_eco9750, w_eco9751, w_eco9752, w_eco9753, w_eco9754, w_eco9755, w_eco9756, w_eco9757, w_eco9758, w_eco9759, w_eco9760, w_eco9761, w_eco9762, w_eco9763, w_eco9764, w_eco9765, w_eco9766, w_eco9767, w_eco9768, w_eco9769, w_eco9770, w_eco9771, w_eco9772, w_eco9773, w_eco9774, w_eco9775, w_eco9776, w_eco9777, w_eco9778, w_eco9779, w_eco9780, w_eco9781, w_eco9782, w_eco9783, w_eco9784, w_eco9785, w_eco9786, w_eco9787, w_eco9788, w_eco9789, w_eco9790, w_eco9791, w_eco9792, w_eco9793, w_eco9794, w_eco9795, w_eco9796, w_eco9797, w_eco9798, w_eco9799, w_eco9800, w_eco9801, w_eco9802, w_eco9803, w_eco9804, w_eco9805, w_eco9806, w_eco9807, w_eco9808, w_eco9809, w_eco9810, w_eco9811, w_eco9812, w_eco9813, w_eco9814, w_eco9815, w_eco9816, w_eco9817, w_eco9818, w_eco9819, w_eco9820, w_eco9821, w_eco9822, w_eco9823, w_eco9824, w_eco9825, w_eco9826, w_eco9827, w_eco9828, w_eco9829, w_eco9830, w_eco9831, w_eco9832, w_eco9833, w_eco9834, w_eco9835, w_eco9836, w_eco9837, w_eco9838, w_eco9839, w_eco9840, w_eco9841, w_eco9842, w_eco9843, w_eco9844, w_eco9845, w_eco9846, w_eco9847, w_eco9848, w_eco9849, w_eco9850, w_eco9851, w_eco9852, w_eco9853, w_eco9854, w_eco9855, w_eco9856, w_eco9857, w_eco9858, w_eco9859, w_eco9860, w_eco9861, w_eco9862, w_eco9863, w_eco9864, w_eco9865, w_eco9866, w_eco9867, w_eco9868, w_eco9869, w_eco9870, w_eco9871, w_eco9872, w_eco9873, w_eco9874, w_eco9875, w_eco9876, w_eco9877, w_eco9878, w_eco9879, w_eco9880, w_eco9881, w_eco9882, w_eco9883, w_eco9884, w_eco9885, w_eco9886, w_eco9887, w_eco9888, w_eco9889, w_eco9890, w_eco9891, w_eco9892, w_eco9893, w_eco9894, w_eco9895, w_eco9896, w_eco9897, w_eco9898, w_eco9899, w_eco9900, w_eco9901, w_eco9902, w_eco9903, w_eco9904, w_eco9905, w_eco9906, w_eco9907, w_eco9908, w_eco9909, w_eco9910, w_eco9911, w_eco9912, w_eco9913, w_eco9914, w_eco9915, w_eco9916, w_eco9917, w_eco9918, w_eco9919, w_eco9920, w_eco9921, w_eco9922, w_eco9923, w_eco9924, w_eco9925, w_eco9926, w_eco9927, w_eco9928, w_eco9929, w_eco9930, w_eco9931, w_eco9932, w_eco9933, w_eco9934, w_eco9935, w_eco9936, w_eco9937, w_eco9938, w_eco9939, w_eco9940, w_eco9941, w_eco9942, w_eco9943, w_eco9944, w_eco9945, w_eco9946, w_eco9947, w_eco9948, w_eco9949, w_eco9950, w_eco9951, w_eco9952, w_eco9953, w_eco9954, w_eco9955, w_eco9956, w_eco9957, w_eco9958, w_eco9959, w_eco9960, w_eco9961, w_eco9962, w_eco9963, w_eco9964, w_eco9965, w_eco9966, w_eco9967, w_eco9968, w_eco9969, w_eco9970, w_eco9971, w_eco9972, w_eco9973, w_eco9974, w_eco9975, w_eco9976, w_eco9977, w_eco9978, w_eco9979, w_eco9980, w_eco9981, w_eco9982, w_eco9983, w_eco9984, w_eco9985, w_eco9986, w_eco9987, w_eco9988, w_eco9989, w_eco9990, w_eco9991, w_eco9992, w_eco9993, w_eco9994, w_eco9995, w_eco9996, w_eco9997, w_eco9998, w_eco9999, w_eco10000, w_eco10001, w_eco10002, w_eco10003, w_eco10004, w_eco10005, w_eco10006, w_eco10007, w_eco10008, w_eco10009, w_eco10010, w_eco10011, w_eco10012, w_eco10013, w_eco10014, w_eco10015, w_eco10016, w_eco10017, w_eco10018, w_eco10019, w_eco10020, w_eco10021, w_eco10022, w_eco10023, w_eco10024, w_eco10025, w_eco10026, w_eco10027, w_eco10028, w_eco10029, w_eco10030, w_eco10031, w_eco10032, w_eco10033, w_eco10034, w_eco10035, w_eco10036, w_eco10037, w_eco10038, w_eco10039, w_eco10040, w_eco10041, w_eco10042, w_eco10043, w_eco10044, w_eco10045, w_eco10046, w_eco10047, w_eco10048, w_eco10049, w_eco10050, w_eco10051, w_eco10052, w_eco10053, w_eco10054, w_eco10055, w_eco10056, w_eco10057, w_eco10058, w_eco10059, w_eco10060, w_eco10061, w_eco10062, w_eco10063, w_eco10064, w_eco10065, w_eco10066, w_eco10067, w_eco10068, w_eco10069, w_eco10070, w_eco10071, w_eco10072, w_eco10073, w_eco10074, w_eco10075, w_eco10076, w_eco10077, w_eco10078, w_eco10079, w_eco10080, w_eco10081, w_eco10082, w_eco10083, w_eco10084, w_eco10085, w_eco10086, w_eco10087, w_eco10088, w_eco10089, w_eco10090, w_eco10091, w_eco10092, w_eco10093, w_eco10094, w_eco10095, w_eco10096, w_eco10097, w_eco10098, w_eco10099, w_eco10100, w_eco10101, w_eco10102, w_eco10103, w_eco10104, w_eco10105, w_eco10106, w_eco10107, w_eco10108, w_eco10109, w_eco10110, w_eco10111, w_eco10112, w_eco10113, w_eco10114, w_eco10115, w_eco10116, w_eco10117, w_eco10118, w_eco10119, w_eco10120, w_eco10121, w_eco10122, w_eco10123, w_eco10124, w_eco10125, w_eco10126, w_eco10127, w_eco10128, w_eco10129, w_eco10130, w_eco10131, w_eco10132, w_eco10133, w_eco10134, w_eco10135, w_eco10136, w_eco10137, w_eco10138, w_eco10139, w_eco10140, w_eco10141, w_eco10142, w_eco10143, w_eco10144, w_eco10145, w_eco10146, w_eco10147, w_eco10148, w_eco10149, w_eco10150, w_eco10151, w_eco10152, w_eco10153, w_eco10154, w_eco10155, w_eco10156, w_eco10157, w_eco10158, w_eco10159, w_eco10160, w_eco10161, w_eco10162, w_eco10163, w_eco10164, w_eco10165, w_eco10166, w_eco10167, w_eco10168, w_eco10169, w_eco10170, w_eco10171, w_eco10172, w_eco10173, w_eco10174, w_eco10175, w_eco10176, w_eco10177, w_eco10178, w_eco10179, w_eco10180, w_eco10181, w_eco10182, w_eco10183, w_eco10184, w_eco10185, w_eco10186, w_eco10187, w_eco10188, w_eco10189, w_eco10190, w_eco10191, w_eco10192, w_eco10193, w_eco10194, w_eco10195, w_eco10196, w_eco10197, w_eco10198, w_eco10199, w_eco10200, w_eco10201, w_eco10202, w_eco10203, w_eco10204, w_eco10205, sub_wire8, w_eco10206, w_eco10207, w_eco10208, w_eco10209, w_eco10210, w_eco10211, w_eco10212, w_eco10213, w_eco10214, w_eco10215, w_eco10216, w_eco10217, w_eco10218, w_eco10219, w_eco10220, w_eco10221, w_eco10222, w_eco10223, w_eco10224, w_eco10225, w_eco10226, w_eco10227, w_eco10228, w_eco10229, w_eco10230, w_eco10231, w_eco10232, w_eco10233, w_eco10234, w_eco10235, w_eco10236, w_eco10237, w_eco10238, w_eco10239, w_eco10240, w_eco10241, w_eco10242, w_eco10243, w_eco10244, w_eco10245, w_eco10246, w_eco10247, w_eco10248, w_eco10249, w_eco10250, w_eco10251, w_eco10252, w_eco10253, w_eco10254, w_eco10255, w_eco10256, w_eco10257, w_eco10258, w_eco10259, w_eco10260, w_eco10261, w_eco10262, w_eco10263, w_eco10264, w_eco10265, w_eco10266, w_eco10267, w_eco10268, w_eco10269, w_eco10270, w_eco10271, w_eco10272, w_eco10273, w_eco10274, w_eco10275, w_eco10276, w_eco10277, w_eco10278, w_eco10279, w_eco10280, w_eco10281, w_eco10282, w_eco10283, w_eco10284, w_eco10285, w_eco10286, w_eco10287, w_eco10288, w_eco10289, w_eco10290, w_eco10291, w_eco10292, w_eco10293, w_eco10294, w_eco10295, w_eco10296, w_eco10297, w_eco10298, w_eco10299, w_eco10300, w_eco10301, w_eco10302, w_eco10303, w_eco10304, w_eco10305, w_eco10306, w_eco10307, w_eco10308, w_eco10309, w_eco10310, w_eco10311, w_eco10312, w_eco10313, w_eco10314, w_eco10315, w_eco10316, w_eco10317, w_eco10318, w_eco10319, w_eco10320, w_eco10321, w_eco10322, w_eco10323, w_eco10324, w_eco10325, w_eco10326, w_eco10327, w_eco10328, w_eco10329, w_eco10330, w_eco10331, w_eco10332, w_eco10333, w_eco10334, w_eco10335, w_eco10336, w_eco10337, w_eco10338, w_eco10339, w_eco10340, w_eco10341, w_eco10342, w_eco10343, w_eco10344, w_eco10345, w_eco10346, w_eco10347, w_eco10348, w_eco10349, w_eco10350, w_eco10351, w_eco10352, w_eco10353, w_eco10354, w_eco10355, w_eco10356, w_eco10357, w_eco10358, w_eco10359, w_eco10360, w_eco10361, w_eco10362, w_eco10363, w_eco10364, w_eco10365, w_eco10366, w_eco10367, w_eco10368, w_eco10369, w_eco10370, w_eco10371, w_eco10372, w_eco10373, w_eco10374, w_eco10375, w_eco10376, w_eco10377, w_eco10378, w_eco10379, w_eco10380, w_eco10381, w_eco10382, w_eco10383, w_eco10384, w_eco10385, w_eco10386, w_eco10387, w_eco10388, w_eco10389, w_eco10390, w_eco10391, w_eco10392, w_eco10393, w_eco10394, w_eco10395, w_eco10396, w_eco10397, w_eco10398, w_eco10399, w_eco10400, w_eco10401, w_eco10402, w_eco10403, w_eco10404, w_eco10405, w_eco10406, w_eco10407, w_eco10408, w_eco10409, w_eco10410, w_eco10411, w_eco10412, w_eco10413, w_eco10414, w_eco10415, w_eco10416, w_eco10417, w_eco10418, w_eco10419, w_eco10420, w_eco10421, w_eco10422, w_eco10423, w_eco10424, w_eco10425, w_eco10426, w_eco10427, w_eco10428, w_eco10429, w_eco10430, w_eco10431, w_eco10432, w_eco10433, w_eco10434, w_eco10435, w_eco10436, w_eco10437, w_eco10438, w_eco10439, w_eco10440, w_eco10441, w_eco10442, w_eco10443, w_eco10444, w_eco10445, w_eco10446, w_eco10447, w_eco10448, w_eco10449, w_eco10450, w_eco10451, w_eco10452, w_eco10453, w_eco10454, w_eco10455, w_eco10456, w_eco10457, w_eco10458, w_eco10459, w_eco10460, w_eco10461, w_eco10462, w_eco10463, w_eco10464, w_eco10465, w_eco10466, w_eco10467, w_eco10468, w_eco10469, w_eco10470, w_eco10471, w_eco10472, w_eco10473, w_eco10474, w_eco10475, w_eco10476, w_eco10477, w_eco10478, w_eco10479, w_eco10480, w_eco10481, w_eco10482, w_eco10483, w_eco10484, w_eco10485, w_eco10486, w_eco10487, w_eco10488, w_eco10489, w_eco10490, w_eco10491, w_eco10492, w_eco10493, w_eco10494, w_eco10495, w_eco10496, w_eco10497, w_eco10498, w_eco10499, w_eco10500, w_eco10501, w_eco10502, w_eco10503, w_eco10504, w_eco10505, w_eco10506, w_eco10507, w_eco10508, w_eco10509, w_eco10510, w_eco10511, w_eco10512, w_eco10513, w_eco10514, w_eco10515, w_eco10516, w_eco10517, w_eco10518, w_eco10519, w_eco10520, w_eco10521, w_eco10522, w_eco10523, w_eco10524, w_eco10525, w_eco10526, w_eco10527, w_eco10528, w_eco10529, w_eco10530, w_eco10531, w_eco10532, w_eco10533, w_eco10534, w_eco10535, w_eco10536, w_eco10537, w_eco10538, w_eco10539, w_eco10540, w_eco10541, w_eco10542, w_eco10543, w_eco10544, w_eco10545, w_eco10546, w_eco10547, w_eco10548, w_eco10549, w_eco10550, w_eco10551, w_eco10552, w_eco10553, w_eco10554, w_eco10555, w_eco10556, w_eco10557, w_eco10558, w_eco10559, w_eco10560, w_eco10561, w_eco10562, w_eco10563, w_eco10564, w_eco10565, w_eco10566, w_eco10567, w_eco10568, w_eco10569, w_eco10570, w_eco10571, w_eco10572, w_eco10573, w_eco10574, w_eco10575, w_eco10576, w_eco10577, w_eco10578, w_eco10579, w_eco10580, w_eco10581, w_eco10582, w_eco10583, w_eco10584, w_eco10585, w_eco10586, w_eco10587, w_eco10588, w_eco10589, w_eco10590, w_eco10591, w_eco10592, w_eco10593, w_eco10594, w_eco10595, w_eco10596, w_eco10597, w_eco10598, w_eco10599, w_eco10600, w_eco10601, w_eco10602, w_eco10603, w_eco10604, w_eco10605, w_eco10606, w_eco10607, w_eco10608, w_eco10609, w_eco10610, w_eco10611, w_eco10612, w_eco10613, w_eco10614, w_eco10615, w_eco10616, w_eco10617, w_eco10618, w_eco10619, w_eco10620, w_eco10621, w_eco10622, w_eco10623, w_eco10624, w_eco10625, w_eco10626, w_eco10627, w_eco10628, w_eco10629, w_eco10630, w_eco10631, w_eco10632, w_eco10633, w_eco10634, w_eco10635, w_eco10636, w_eco10637, w_eco10638, w_eco10639, w_eco10640, w_eco10641, w_eco10642, w_eco10643, w_eco10644, w_eco10645, w_eco10646, w_eco10647, w_eco10648, w_eco10649, w_eco10650, w_eco10651, w_eco10652, w_eco10653, w_eco10654, w_eco10655, w_eco10656, w_eco10657, w_eco10658, w_eco10659, w_eco10660, w_eco10661, w_eco10662, w_eco10663, w_eco10664, w_eco10665, w_eco10666, w_eco10667, w_eco10668, w_eco10669, w_eco10670, w_eco10671, w_eco10672, w_eco10673, w_eco10674, w_eco10675, w_eco10676, w_eco10677, w_eco10678, w_eco10679, w_eco10680, w_eco10681, w_eco10682, w_eco10683, w_eco10684, w_eco10685, w_eco10686, w_eco10687, w_eco10688, w_eco10689, w_eco10690, w_eco10691, w_eco10692, w_eco10693, w_eco10694, w_eco10695, w_eco10696, w_eco10697, w_eco10698, w_eco10699, w_eco10700, w_eco10701, w_eco10702, w_eco10703, w_eco10704, w_eco10705, w_eco10706, w_eco10707, w_eco10708, w_eco10709, w_eco10710, w_eco10711, w_eco10712, w_eco10713, w_eco10714, w_eco10715, w_eco10716, w_eco10717, w_eco10718, w_eco10719, w_eco10720, w_eco10721, w_eco10722, w_eco10723, w_eco10724, w_eco10725, w_eco10726, w_eco10727, w_eco10728, w_eco10729, w_eco10730, w_eco10731, w_eco10732, w_eco10733, w_eco10734, w_eco10735, w_eco10736, w_eco10737, w_eco10738, w_eco10739, w_eco10740, w_eco10741, w_eco10742, w_eco10743, w_eco10744, w_eco10745, w_eco10746, w_eco10747, w_eco10748, w_eco10749, w_eco10750, w_eco10751, w_eco10752, w_eco10753, w_eco10754, w_eco10755, w_eco10756, w_eco10757, w_eco10758, w_eco10759, w_eco10760, w_eco10761, w_eco10762, w_eco10763, w_eco10764, w_eco10765, w_eco10766, w_eco10767, w_eco10768, w_eco10769, w_eco10770, w_eco10771, w_eco10772, w_eco10773, w_eco10774, w_eco10775, w_eco10776, w_eco10777, w_eco10778, w_eco10779, w_eco10780, w_eco10781, w_eco10782, w_eco10783, w_eco10784, w_eco10785, w_eco10786, w_eco10787, w_eco10788, w_eco10789, w_eco10790, w_eco10791, w_eco10792, w_eco10793, w_eco10794, w_eco10795, w_eco10796, w_eco10797, w_eco10798, w_eco10799, w_eco10800, w_eco10801, w_eco10802, w_eco10803, w_eco10804, w_eco10805, w_eco10806, w_eco10807, w_eco10808, w_eco10809, w_eco10810, w_eco10811, w_eco10812, w_eco10813, w_eco10814, w_eco10815, w_eco10816, w_eco10817, w_eco10818, w_eco10819, w_eco10820, w_eco10821, w_eco10822, w_eco10823, w_eco10824, w_eco10825, w_eco10826, w_eco10827, w_eco10828, w_eco10829, w_eco10830, w_eco10831, w_eco10832, w_eco10833, w_eco10834, w_eco10835, w_eco10836, w_eco10837, w_eco10838, w_eco10839, w_eco10840, w_eco10841, w_eco10842, w_eco10843, w_eco10844, w_eco10845, w_eco10846, w_eco10847, w_eco10848, w_eco10849, w_eco10850, w_eco10851, w_eco10852, w_eco10853, w_eco10854, w_eco10855, w_eco10856, w_eco10857, w_eco10858, w_eco10859, w_eco10860, w_eco10861, w_eco10862, w_eco10863, w_eco10864, w_eco10865, w_eco10866, w_eco10867, w_eco10868, w_eco10869, w_eco10870, w_eco10871, w_eco10872, w_eco10873, w_eco10874, w_eco10875, w_eco10876, w_eco10877, w_eco10878, w_eco10879, w_eco10880, w_eco10881, w_eco10882, w_eco10883, w_eco10884, w_eco10885, w_eco10886, w_eco10887, w_eco10888, w_eco10889, w_eco10890, w_eco10891, w_eco10892, w_eco10893, w_eco10894, w_eco10895, w_eco10896, w_eco10897, w_eco10898, w_eco10899, w_eco10900, w_eco10901, w_eco10902, w_eco10903, w_eco10904, w_eco10905, w_eco10906, w_eco10907, w_eco10908, w_eco10909, w_eco10910, w_eco10911, w_eco10912, w_eco10913, w_eco10914, w_eco10915, w_eco10916, w_eco10917, w_eco10918, w_eco10919, w_eco10920, w_eco10921, w_eco10922, w_eco10923, w_eco10924, w_eco10925, sub_wire9, w_eco10926, w_eco10927, w_eco10928, w_eco10929, w_eco10930, w_eco10931, w_eco10932, w_eco10933, w_eco10934, w_eco10935, w_eco10936, w_eco10937, w_eco10938, w_eco10939, w_eco10940, w_eco10941, w_eco10942, w_eco10943, w_eco10944, w_eco10945, w_eco10946, w_eco10947, w_eco10948, w_eco10949, w_eco10950, w_eco10951, w_eco10952, w_eco10953, w_eco10954, w_eco10955, w_eco10956, w_eco10957, w_eco10958, w_eco10959, w_eco10960, w_eco10961, w_eco10962, w_eco10963, w_eco10964, w_eco10965, w_eco10966, w_eco10967, w_eco10968, w_eco10969, w_eco10970, w_eco10971, w_eco10972, w_eco10973, w_eco10974, w_eco10975, w_eco10976, w_eco10977, w_eco10978, w_eco10979, w_eco10980, w_eco10981, w_eco10982, w_eco10983, w_eco10984, w_eco10985, w_eco10986, w_eco10987, w_eco10988, w_eco10989, w_eco10990, w_eco10991, w_eco10992, w_eco10993, w_eco10994, w_eco10995, w_eco10996, w_eco10997, w_eco10998, w_eco10999, w_eco11000, w_eco11001, w_eco11002, w_eco11003, w_eco11004, w_eco11005, w_eco11006, w_eco11007, w_eco11008, w_eco11009, w_eco11010, w_eco11011, w_eco11012, w_eco11013, w_eco11014, w_eco11015, w_eco11016, w_eco11017, w_eco11018, w_eco11019, w_eco11020, w_eco11021, w_eco11022, w_eco11023, w_eco11024, w_eco11025, w_eco11026, w_eco11027, w_eco11028, w_eco11029, w_eco11030, w_eco11031, w_eco11032, w_eco11033, w_eco11034, w_eco11035, w_eco11036, w_eco11037, w_eco11038, w_eco11039, w_eco11040, w_eco11041, w_eco11042, w_eco11043, w_eco11044, w_eco11045, w_eco11046, w_eco11047, w_eco11048, w_eco11049, w_eco11050, w_eco11051, w_eco11052, w_eco11053, w_eco11054, w_eco11055, w_eco11056, w_eco11057, w_eco11058, w_eco11059, w_eco11060, w_eco11061, w_eco11062, w_eco11063, w_eco11064, w_eco11065, w_eco11066, w_eco11067, w_eco11068, w_eco11069, w_eco11070, w_eco11071, w_eco11072, w_eco11073, w_eco11074, w_eco11075, w_eco11076, w_eco11077, w_eco11078, w_eco11079, w_eco11080, w_eco11081, w_eco11082, w_eco11083, w_eco11084, w_eco11085, w_eco11086, w_eco11087, w_eco11088, w_eco11089, w_eco11090, w_eco11091, w_eco11092, w_eco11093, w_eco11094, w_eco11095, w_eco11096, w_eco11097, w_eco11098, w_eco11099, w_eco11100, w_eco11101, w_eco11102, w_eco11103, w_eco11104, w_eco11105, w_eco11106, w_eco11107, w_eco11108, w_eco11109, w_eco11110, w_eco11111, w_eco11112, w_eco11113, w_eco11114, w_eco11115, w_eco11116, w_eco11117, w_eco11118, w_eco11119, w_eco11120, w_eco11121, w_eco11122, w_eco11123, w_eco11124, w_eco11125, w_eco11126, w_eco11127, w_eco11128, w_eco11129, w_eco11130, w_eco11131, w_eco11132, w_eco11133, w_eco11134, w_eco11135, w_eco11136, w_eco11137, w_eco11138, w_eco11139, w_eco11140, w_eco11141, w_eco11142, w_eco11143, w_eco11144, w_eco11145, w_eco11146, w_eco11147, w_eco11148, w_eco11149, w_eco11150, w_eco11151, w_eco11152, w_eco11153, w_eco11154, w_eco11155, w_eco11156, w_eco11157, w_eco11158, w_eco11159, w_eco11160, w_eco11161, w_eco11162, w_eco11163, w_eco11164, w_eco11165, w_eco11166, w_eco11167, w_eco11168, w_eco11169, w_eco11170, w_eco11171, w_eco11172, w_eco11173, w_eco11174, w_eco11175, w_eco11176, w_eco11177, w_eco11178, w_eco11179, w_eco11180, w_eco11181, w_eco11182, w_eco11183, w_eco11184, w_eco11185, w_eco11186, w_eco11187, w_eco11188, w_eco11189, w_eco11190, w_eco11191, w_eco11192, w_eco11193, w_eco11194, w_eco11195, w_eco11196, w_eco11197, w_eco11198, w_eco11199, w_eco11200, w_eco11201, w_eco11202, w_eco11203, w_eco11204, w_eco11205, w_eco11206, w_eco11207, w_eco11208, w_eco11209, w_eco11210, w_eco11211, w_eco11212, w_eco11213, w_eco11214, w_eco11215, w_eco11216, w_eco11217, w_eco11218, w_eco11219, w_eco11220, w_eco11221, w_eco11222, w_eco11223, w_eco11224, w_eco11225, w_eco11226, w_eco11227, w_eco11228, w_eco11229, w_eco11230, w_eco11231, w_eco11232, w_eco11233, w_eco11234, w_eco11235, w_eco11236, w_eco11237, w_eco11238, w_eco11239, w_eco11240, w_eco11241, w_eco11242, w_eco11243, w_eco11244, w_eco11245, w_eco11246, w_eco11247, w_eco11248, w_eco11249, w_eco11250, w_eco11251, w_eco11252, w_eco11253, w_eco11254, w_eco11255, w_eco11256, w_eco11257, w_eco11258, w_eco11259, w_eco11260, w_eco11261, w_eco11262, w_eco11263, w_eco11264, w_eco11265, w_eco11266, w_eco11267, w_eco11268, w_eco11269, w_eco11270, w_eco11271, w_eco11272, w_eco11273, w_eco11274, w_eco11275, w_eco11276, w_eco11277, w_eco11278, w_eco11279, w_eco11280, w_eco11281, w_eco11282, w_eco11283, w_eco11284, w_eco11285, w_eco11286, w_eco11287, w_eco11288, w_eco11289, w_eco11290, w_eco11291, w_eco11292, w_eco11293, w_eco11294, w_eco11295, w_eco11296, w_eco11297, w_eco11298, w_eco11299, w_eco11300, w_eco11301, w_eco11302, w_eco11303, w_eco11304, w_eco11305, w_eco11306, w_eco11307, w_eco11308, w_eco11309, w_eco11310, w_eco11311, w_eco11312, w_eco11313, w_eco11314, w_eco11315, w_eco11316, w_eco11317, w_eco11318, w_eco11319, w_eco11320, w_eco11321, w_eco11322, w_eco11323, w_eco11324, w_eco11325, w_eco11326, w_eco11327, w_eco11328, w_eco11329, w_eco11330, w_eco11331, w_eco11332, w_eco11333, w_eco11334, w_eco11335, w_eco11336, w_eco11337, w_eco11338, w_eco11339, w_eco11340, w_eco11341, w_eco11342, w_eco11343, w_eco11344, w_eco11345, w_eco11346, w_eco11347, w_eco11348, w_eco11349, w_eco11350, w_eco11351, w_eco11352, w_eco11353, w_eco11354, w_eco11355, w_eco11356, w_eco11357, w_eco11358, w_eco11359, w_eco11360, w_eco11361, w_eco11362, w_eco11363, w_eco11364, w_eco11365, w_eco11366, w_eco11367, w_eco11368, w_eco11369, w_eco11370, w_eco11371, w_eco11372, w_eco11373, w_eco11374, w_eco11375, w_eco11376, w_eco11377, w_eco11378, w_eco11379, w_eco11380, w_eco11381, w_eco11382, w_eco11383, w_eco11384, w_eco11385, w_eco11386, w_eco11387, w_eco11388, w_eco11389, w_eco11390, w_eco11391, w_eco11392, w_eco11393, w_eco11394, w_eco11395, w_eco11396, w_eco11397, w_eco11398, w_eco11399, w_eco11400, w_eco11401, w_eco11402, w_eco11403, w_eco11404, w_eco11405, w_eco11406, w_eco11407, w_eco11408, w_eco11409, w_eco11410, w_eco11411, w_eco11412, w_eco11413, w_eco11414, w_eco11415, w_eco11416, w_eco11417, w_eco11418, w_eco11419, w_eco11420, w_eco11421, w_eco11422, w_eco11423, w_eco11424, w_eco11425, w_eco11426, w_eco11427, w_eco11428, w_eco11429, w_eco11430, w_eco11431, w_eco11432, w_eco11433, w_eco11434, w_eco11435, w_eco11436, w_eco11437, w_eco11438, w_eco11439, w_eco11440, w_eco11441, w_eco11442, w_eco11443, w_eco11444, w_eco11445, w_eco11446, w_eco11447, w_eco11448, w_eco11449, w_eco11450, w_eco11451, w_eco11452, w_eco11453, w_eco11454, w_eco11455, w_eco11456, w_eco11457, w_eco11458, w_eco11459, w_eco11460, w_eco11461, w_eco11462, w_eco11463, w_eco11464, w_eco11465, w_eco11466, w_eco11467, w_eco11468, w_eco11469, w_eco11470, w_eco11471, w_eco11472, w_eco11473, w_eco11474, w_eco11475, w_eco11476, w_eco11477, w_eco11478, w_eco11479, w_eco11480, w_eco11481, w_eco11482, w_eco11483, w_eco11484, w_eco11485, w_eco11486, w_eco11487, w_eco11488, w_eco11489, w_eco11490, w_eco11491, w_eco11492, w_eco11493, w_eco11494, w_eco11495, w_eco11496, w_eco11497, w_eco11498, w_eco11499, w_eco11500, w_eco11501, w_eco11502, w_eco11503, w_eco11504, w_eco11505, w_eco11506, w_eco11507, w_eco11508, w_eco11509, w_eco11510, w_eco11511, w_eco11512, w_eco11513, w_eco11514, w_eco11515, w_eco11516, w_eco11517, w_eco11518, w_eco11519, w_eco11520, w_eco11521, w_eco11522, w_eco11523, w_eco11524, w_eco11525, w_eco11526, w_eco11527, w_eco11528, w_eco11529, w_eco11530, w_eco11531, w_eco11532, w_eco11533, w_eco11534, w_eco11535, w_eco11536, w_eco11537, w_eco11538, w_eco11539, w_eco11540, w_eco11541, w_eco11542, w_eco11543, w_eco11544, w_eco11545, w_eco11546, w_eco11547, w_eco11548, w_eco11549, w_eco11550, w_eco11551, w_eco11552, w_eco11553, w_eco11554, w_eco11555, w_eco11556, w_eco11557, w_eco11558, w_eco11559, w_eco11560, w_eco11561, w_eco11562, w_eco11563, w_eco11564, w_eco11565, w_eco11566, w_eco11567, w_eco11568, w_eco11569, w_eco11570, w_eco11571, w_eco11572, w_eco11573, w_eco11574, w_eco11575, w_eco11576, w_eco11577, w_eco11578, w_eco11579, w_eco11580, w_eco11581, w_eco11582, w_eco11583, w_eco11584, w_eco11585, w_eco11586, w_eco11587, w_eco11588, w_eco11589, w_eco11590, w_eco11591, w_eco11592, w_eco11593, w_eco11594, w_eco11595, w_eco11596, w_eco11597, w_eco11598, w_eco11599, w_eco11600, w_eco11601, w_eco11602, w_eco11603, w_eco11604, w_eco11605, w_eco11606, w_eco11607, w_eco11608, w_eco11609, w_eco11610, w_eco11611, w_eco11612, w_eco11613, w_eco11614, w_eco11615, w_eco11616, w_eco11617, w_eco11618, w_eco11619, w_eco11620, w_eco11621, w_eco11622, w_eco11623, w_eco11624, w_eco11625, w_eco11626, w_eco11627, w_eco11628, w_eco11629, w_eco11630, w_eco11631, w_eco11632, w_eco11633, w_eco11634, w_eco11635, w_eco11636, w_eco11637, w_eco11638, w_eco11639, w_eco11640, w_eco11641, w_eco11642, w_eco11643, w_eco11644, w_eco11645, w_eco11646, w_eco11647, w_eco11648, w_eco11649, w_eco11650, w_eco11651, w_eco11652, w_eco11653, w_eco11654, w_eco11655, w_eco11656, w_eco11657, w_eco11658, w_eco11659, w_eco11660, w_eco11661, w_eco11662, w_eco11663, w_eco11664, w_eco11665, w_eco11666, w_eco11667, w_eco11668, w_eco11669, w_eco11670, w_eco11671, w_eco11672, w_eco11673, w_eco11674, w_eco11675, w_eco11676, w_eco11677, w_eco11678, w_eco11679, w_eco11680, w_eco11681, w_eco11682, w_eco11683, w_eco11684, w_eco11685, w_eco11686, w_eco11687, w_eco11688, w_eco11689, w_eco11690, w_eco11691, w_eco11692, w_eco11693, w_eco11694, w_eco11695, w_eco11696, w_eco11697, w_eco11698, w_eco11699, w_eco11700, w_eco11701, w_eco11702, w_eco11703, w_eco11704, w_eco11705, w_eco11706, w_eco11707, w_eco11708, w_eco11709, w_eco11710, w_eco11711, w_eco11712, w_eco11713, w_eco11714, w_eco11715, w_eco11716, w_eco11717, w_eco11718, w_eco11719, w_eco11720, w_eco11721, w_eco11722, w_eco11723, w_eco11724, w_eco11725, w_eco11726, w_eco11727, w_eco11728, w_eco11729, w_eco11730, w_eco11731, w_eco11732, w_eco11733, w_eco11734, w_eco11735, w_eco11736, w_eco11737, w_eco11738, w_eco11739, w_eco11740, w_eco11741, w_eco11742, w_eco11743, w_eco11744, w_eco11745, w_eco11746, w_eco11747, w_eco11748, w_eco11749, w_eco11750, w_eco11751, w_eco11752, w_eco11753, w_eco11754, w_eco11755, w_eco11756, w_eco11757, w_eco11758, w_eco11759, w_eco11760, w_eco11761, w_eco11762, w_eco11763, w_eco11764, w_eco11765, w_eco11766, w_eco11767, w_eco11768, w_eco11769, w_eco11770, w_eco11771, w_eco11772, w_eco11773, w_eco11774, w_eco11775, w_eco11776, w_eco11777, w_eco11778, w_eco11779, w_eco11780, w_eco11781, w_eco11782, w_eco11783, w_eco11784, w_eco11785, w_eco11786, w_eco11787, w_eco11788, w_eco11789, w_eco11790, w_eco11791, w_eco11792, w_eco11793, w_eco11794, w_eco11795, w_eco11796, w_eco11797, w_eco11798, w_eco11799, w_eco11800, w_eco11801, w_eco11802, w_eco11803, w_eco11804, w_eco11805, w_eco11806, w_eco11807, w_eco11808, w_eco11809, w_eco11810, w_eco11811, w_eco11812, w_eco11813, w_eco11814, w_eco11815, w_eco11816, w_eco11817, w_eco11818, w_eco11819, w_eco11820, w_eco11821, w_eco11822, w_eco11823, w_eco11824, w_eco11825, w_eco11826, w_eco11827, w_eco11828, w_eco11829, w_eco11830, w_eco11831, w_eco11832, w_eco11833, w_eco11834, w_eco11835, w_eco11836, w_eco11837, w_eco11838, w_eco11839, w_eco11840, w_eco11841, w_eco11842, w_eco11843, w_eco11844, w_eco11845, w_eco11846, w_eco11847, w_eco11848, w_eco11849, w_eco11850, w_eco11851, w_eco11852, w_eco11853, w_eco11854, w_eco11855, w_eco11856, w_eco11857, w_eco11858, w_eco11859, w_eco11860, w_eco11861, w_eco11862, w_eco11863, w_eco11864, w_eco11865, w_eco11866, w_eco11867, w_eco11868, w_eco11869, w_eco11870, w_eco11871, w_eco11872, w_eco11873, w_eco11874, w_eco11875, w_eco11876, w_eco11877, w_eco11878, w_eco11879, w_eco11880, w_eco11881, w_eco11882, w_eco11883, w_eco11884, w_eco11885, w_eco11886, w_eco11887, w_eco11888, w_eco11889, w_eco11890, w_eco11891, w_eco11892, w_eco11893, w_eco11894, w_eco11895, w_eco11896, w_eco11897, w_eco11898, w_eco11899, w_eco11900, w_eco11901, w_eco11902, w_eco11903, w_eco11904, w_eco11905, w_eco11906, w_eco11907, w_eco11908, w_eco11909, w_eco11910, w_eco11911, w_eco11912, w_eco11913, w_eco11914, w_eco11915, w_eco11916, w_eco11917, w_eco11918, w_eco11919, w_eco11920, w_eco11921, w_eco11922, w_eco11923, w_eco11924, w_eco11925, w_eco11926, w_eco11927, w_eco11928, w_eco11929, w_eco11930, w_eco11931, w_eco11932, w_eco11933, w_eco11934, w_eco11935, w_eco11936, w_eco11937, w_eco11938, w_eco11939, w_eco11940, w_eco11941, w_eco11942, w_eco11943, w_eco11944, w_eco11945, w_eco11946, w_eco11947, w_eco11948, w_eco11949, w_eco11950, w_eco11951, w_eco11952, w_eco11953, w_eco11954, w_eco11955, w_eco11956, w_eco11957, w_eco11958, w_eco11959, w_eco11960, w_eco11961, w_eco11962, w_eco11963, w_eco11964, w_eco11965, w_eco11966, w_eco11967, w_eco11968, w_eco11969, w_eco11970, w_eco11971, w_eco11972, w_eco11973, w_eco11974, w_eco11975, w_eco11976, w_eco11977, w_eco11978, w_eco11979, w_eco11980, w_eco11981, w_eco11982, w_eco11983, w_eco11984, w_eco11985, w_eco11986, w_eco11987, w_eco11988, w_eco11989, w_eco11990, w_eco11991, w_eco11992, w_eco11993, w_eco11994, w_eco11995, w_eco11996, w_eco11997, w_eco11998, w_eco11999, w_eco12000, w_eco12001, w_eco12002, w_eco12003, w_eco12004, w_eco12005, w_eco12006, w_eco12007, w_eco12008, w_eco12009, w_eco12010, w_eco12011, w_eco12012, w_eco12013, w_eco12014, w_eco12015, w_eco12016, w_eco12017, w_eco12018, w_eco12019, w_eco12020, w_eco12021, w_eco12022, w_eco12023, w_eco12024, w_eco12025, w_eco12026, w_eco12027, w_eco12028, w_eco12029, w_eco12030, w_eco12031, w_eco12032, w_eco12033, w_eco12034, w_eco12035, w_eco12036, w_eco12037, w_eco12038, w_eco12039, w_eco12040, w_eco12041, w_eco12042, w_eco12043, w_eco12044, w_eco12045, w_eco12046, w_eco12047, w_eco12048, w_eco12049, w_eco12050, w_eco12051, w_eco12052, w_eco12053, w_eco12054, w_eco12055, w_eco12056, w_eco12057, w_eco12058, w_eco12059, w_eco12060, w_eco12061, w_eco12062, w_eco12063, w_eco12064, w_eco12065, w_eco12066, w_eco12067, w_eco12068, w_eco12069, w_eco12070, w_eco12071, w_eco12072, w_eco12073, w_eco12074, w_eco12075, w_eco12076, w_eco12077, w_eco12078, w_eco12079, w_eco12080, w_eco12081, w_eco12082, w_eco12083, w_eco12084, w_eco12085, w_eco12086, w_eco12087, w_eco12088, w_eco12089, w_eco12090, w_eco12091, w_eco12092, w_eco12093, w_eco12094, w_eco12095, w_eco12096, w_eco12097, w_eco12098, w_eco12099, w_eco12100, w_eco12101, w_eco12102, w_eco12103, w_eco12104, w_eco12105, w_eco12106, w_eco12107, w_eco12108, w_eco12109, w_eco12110, w_eco12111, w_eco12112, w_eco12113, w_eco12114, w_eco12115, w_eco12116, w_eco12117, w_eco12118, w_eco12119, w_eco12120, w_eco12121, w_eco12122, w_eco12123, w_eco12124, w_eco12125, w_eco12126, w_eco12127, w_eco12128, w_eco12129, w_eco12130, w_eco12131, w_eco12132, w_eco12133, w_eco12134, w_eco12135, w_eco12136, w_eco12137, w_eco12138, w_eco12139, w_eco12140, w_eco12141, w_eco12142, w_eco12143, w_eco12144, w_eco12145, w_eco12146, w_eco12147, w_eco12148, w_eco12149, w_eco12150, w_eco12151, w_eco12152, w_eco12153, w_eco12154, w_eco12155, w_eco12156, w_eco12157, w_eco12158, w_eco12159, w_eco12160, w_eco12161, w_eco12162, w_eco12163, w_eco12164, w_eco12165, w_eco12166, w_eco12167, w_eco12168, w_eco12169, w_eco12170, w_eco12171, w_eco12172, w_eco12173, w_eco12174, w_eco12175, w_eco12176, w_eco12177, w_eco12178, w_eco12179, w_eco12180, w_eco12181, w_eco12182, w_eco12183, w_eco12184, w_eco12185, w_eco12186, w_eco12187, w_eco12188, w_eco12189, w_eco12190, w_eco12191, w_eco12192, w_eco12193, w_eco12194, w_eco12195, w_eco12196, w_eco12197, w_eco12198, w_eco12199, w_eco12200, w_eco12201, w_eco12202, w_eco12203, w_eco12204, w_eco12205, w_eco12206, w_eco12207, w_eco12208, w_eco12209, w_eco12210, w_eco12211, w_eco12212, w_eco12213, w_eco12214, w_eco12215, w_eco12216, w_eco12217, w_eco12218, w_eco12219, w_eco12220, w_eco12221, w_eco12222, w_eco12223, w_eco12224, w_eco12225, w_eco12226, w_eco12227, w_eco12228, w_eco12229, w_eco12230, w_eco12231, w_eco12232, w_eco12233, w_eco12234, w_eco12235, w_eco12236, w_eco12237, w_eco12238, w_eco12239, w_eco12240, w_eco12241, w_eco12242, w_eco12243, w_eco12244, w_eco12245, w_eco12246, w_eco12247, w_eco12248, w_eco12249, w_eco12250, w_eco12251, w_eco12252, w_eco12253, w_eco12254, w_eco12255, w_eco12256, w_eco12257, w_eco12258, w_eco12259, w_eco12260, w_eco12261, w_eco12262, w_eco12263, w_eco12264, w_eco12265, w_eco12266, w_eco12267, w_eco12268, w_eco12269, w_eco12270, w_eco12271, w_eco12272, w_eco12273, w_eco12274, w_eco12275, w_eco12276, w_eco12277, w_eco12278, w_eco12279, w_eco12280, w_eco12281, w_eco12282, w_eco12283, w_eco12284, w_eco12285, w_eco12286, w_eco12287, w_eco12288, w_eco12289, w_eco12290, w_eco12291, w_eco12292, w_eco12293, w_eco12294, w_eco12295, w_eco12296, w_eco12297, w_eco12298, w_eco12299, w_eco12300, w_eco12301, w_eco12302, w_eco12303, w_eco12304, w_eco12305, w_eco12306, w_eco12307, w_eco12308, w_eco12309, w_eco12310, w_eco12311, w_eco12312, w_eco12313, w_eco12314, w_eco12315, w_eco12316, w_eco12317, w_eco12318, w_eco12319, w_eco12320, w_eco12321, w_eco12322, w_eco12323, w_eco12324, w_eco12325, w_eco12326, w_eco12327, w_eco12328, w_eco12329, w_eco12330, w_eco12331, w_eco12332, w_eco12333, w_eco12334, w_eco12335, w_eco12336, w_eco12337, w_eco12338, w_eco12339, w_eco12340, w_eco12341, w_eco12342, w_eco12343, w_eco12344, w_eco12345, w_eco12346, w_eco12347, w_eco12348, w_eco12349, w_eco12350, w_eco12351, w_eco12352, w_eco12353, w_eco12354, w_eco12355, w_eco12356, w_eco12357, w_eco12358, w_eco12359, w_eco12360, w_eco12361, w_eco12362, w_eco12363, w_eco12364, w_eco12365, w_eco12366, w_eco12367, w_eco12368, w_eco12369, w_eco12370, w_eco12371, w_eco12372, w_eco12373, w_eco12374, w_eco12375, w_eco12376, w_eco12377, w_eco12378, w_eco12379, w_eco12380, w_eco12381, w_eco12382, w_eco12383, w_eco12384, w_eco12385, w_eco12386, w_eco12387, w_eco12388, w_eco12389, w_eco12390, w_eco12391, w_eco12392, w_eco12393, w_eco12394, w_eco12395, w_eco12396, w_eco12397, w_eco12398, w_eco12399, w_eco12400, w_eco12401, w_eco12402, w_eco12403, w_eco12404, w_eco12405, w_eco12406, w_eco12407, w_eco12408, w_eco12409, w_eco12410, w_eco12411, w_eco12412, w_eco12413, w_eco12414, w_eco12415, w_eco12416, w_eco12417, w_eco12418, w_eco12419, w_eco12420, w_eco12421, w_eco12422, w_eco12423, w_eco12424, w_eco12425, w_eco12426, w_eco12427, w_eco12428, w_eco12429, w_eco12430, w_eco12431, w_eco12432, w_eco12433, w_eco12434, w_eco12435, w_eco12436, w_eco12437, w_eco12438, w_eco12439, w_eco12440, w_eco12441, w_eco12442, w_eco12443, w_eco12444, w_eco12445, w_eco12446, w_eco12447, w_eco12448, w_eco12449, w_eco12450, w_eco12451, w_eco12452, w_eco12453, w_eco12454, w_eco12455, w_eco12456, w_eco12457, w_eco12458, w_eco12459, w_eco12460, w_eco12461, w_eco12462, w_eco12463, w_eco12464, w_eco12465, w_eco12466, w_eco12467, w_eco12468, w_eco12469, w_eco12470, w_eco12471, w_eco12472, w_eco12473, w_eco12474, w_eco12475, w_eco12476, w_eco12477, w_eco12478, w_eco12479, w_eco12480, w_eco12481, w_eco12482, w_eco12483, w_eco12484, w_eco12485, w_eco12486, w_eco12487, w_eco12488, w_eco12489, w_eco12490, w_eco12491, w_eco12492, w_eco12493, w_eco12494, w_eco12495, w_eco12496, w_eco12497, w_eco12498, w_eco12499, w_eco12500, w_eco12501, w_eco12502, w_eco12503, w_eco12504, w_eco12505, w_eco12506, w_eco12507, w_eco12508, w_eco12509, w_eco12510, w_eco12511, w_eco12512, w_eco12513, w_eco12514, w_eco12515, w_eco12516, w_eco12517, w_eco12518, w_eco12519, w_eco12520, w_eco12521, w_eco12522, w_eco12523, w_eco12524, w_eco12525, w_eco12526, w_eco12527, w_eco12528, w_eco12529, w_eco12530, w_eco12531, w_eco12532, w_eco12533, w_eco12534, w_eco12535, w_eco12536, w_eco12537, w_eco12538, w_eco12539, w_eco12540, w_eco12541, w_eco12542, w_eco12543, w_eco12544, w_eco12545, w_eco12546, w_eco12547, w_eco12548, w_eco12549, w_eco12550, w_eco12551, w_eco12552, w_eco12553, w_eco12554, w_eco12555, w_eco12556, w_eco12557, w_eco12558, w_eco12559, w_eco12560, w_eco12561, w_eco12562, w_eco12563, w_eco12564, w_eco12565, w_eco12566, w_eco12567, w_eco12568, w_eco12569, w_eco12570, w_eco12571, w_eco12572, w_eco12573, w_eco12574, w_eco12575, w_eco12576, w_eco12577, w_eco12578, w_eco12579, w_eco12580, w_eco12581, w_eco12582, w_eco12583, w_eco12584, w_eco12585, w_eco12586, w_eco12587, w_eco12588, w_eco12589, w_eco12590, w_eco12591, w_eco12592, w_eco12593, w_eco12594, w_eco12595, w_eco12596, w_eco12597, w_eco12598, w_eco12599, w_eco12600, w_eco12601, w_eco12602, w_eco12603, w_eco12604, w_eco12605, w_eco12606, w_eco12607, w_eco12608, w_eco12609, w_eco12610, w_eco12611, w_eco12612, w_eco12613, w_eco12614, w_eco12615, w_eco12616, w_eco12617, w_eco12618, w_eco12619, w_eco12620, w_eco12621, w_eco12622, w_eco12623, w_eco12624, w_eco12625, w_eco12626, w_eco12627, w_eco12628, w_eco12629, w_eco12630, w_eco12631, w_eco12632, w_eco12633, w_eco12634, w_eco12635, w_eco12636, w_eco12637, w_eco12638, w_eco12639, w_eco12640, w_eco12641, w_eco12642, w_eco12643, w_eco12644, w_eco12645, w_eco12646, w_eco12647, w_eco12648, w_eco12649, w_eco12650, w_eco12651, w_eco12652, w_eco12653, w_eco12654, w_eco12655, w_eco12656, w_eco12657, w_eco12658, w_eco12659, w_eco12660, w_eco12661, w_eco12662, w_eco12663, w_eco12664, w_eco12665, w_eco12666, w_eco12667, w_eco12668, w_eco12669, w_eco12670, w_eco12671, w_eco12672, w_eco12673, w_eco12674, w_eco12675, w_eco12676, w_eco12677, w_eco12678, w_eco12679, w_eco12680, w_eco12681, w_eco12682, w_eco12683, w_eco12684, w_eco12685, w_eco12686, w_eco12687, w_eco12688, w_eco12689, w_eco12690, w_eco12691, w_eco12692, w_eco12693, w_eco12694, w_eco12695, w_eco12696, w_eco12697, w_eco12698, w_eco12699, w_eco12700, w_eco12701, w_eco12702, w_eco12703, w_eco12704, w_eco12705, w_eco12706, w_eco12707, w_eco12708, w_eco12709, w_eco12710, w_eco12711, w_eco12712, w_eco12713, w_eco12714, w_eco12715, w_eco12716, w_eco12717, w_eco12718, w_eco12719, w_eco12720, w_eco12721, w_eco12722, w_eco12723, w_eco12724, w_eco12725, w_eco12726, w_eco12727, w_eco12728, w_eco12729, w_eco12730, w_eco12731, w_eco12732, w_eco12733, w_eco12734, w_eco12735, w_eco12736, w_eco12737, w_eco12738, w_eco12739, w_eco12740, w_eco12741, w_eco12742, w_eco12743, w_eco12744, w_eco12745, w_eco12746, w_eco12747, w_eco12748, w_eco12749, w_eco12750, w_eco12751, w_eco12752, w_eco12753, w_eco12754, w_eco12755, w_eco12756, w_eco12757, w_eco12758, w_eco12759, w_eco12760, w_eco12761, w_eco12762, w_eco12763, w_eco12764, w_eco12765, w_eco12766, w_eco12767, w_eco12768, w_eco12769, w_eco12770, w_eco12771, w_eco12772, w_eco12773, w_eco12774, w_eco12775, w_eco12776, w_eco12777, w_eco12778, w_eco12779, w_eco12780, w_eco12781, w_eco12782, w_eco12783, w_eco12784, w_eco12785, w_eco12786, w_eco12787, w_eco12788, w_eco12789, w_eco12790, w_eco12791, w_eco12792, w_eco12793, w_eco12794, w_eco12795, w_eco12796, sub_wire10, w_eco12797, w_eco12798, w_eco12799, w_eco12800, w_eco12801, w_eco12802, w_eco12803, w_eco12804, w_eco12805, w_eco12806, w_eco12807, w_eco12808, w_eco12809, w_eco12810, w_eco12811, w_eco12812, w_eco12813, w_eco12814, w_eco12815, w_eco12816, w_eco12817, w_eco12818, w_eco12819, w_eco12820, w_eco12821, w_eco12822, w_eco12823, w_eco12824, w_eco12825, w_eco12826, w_eco12827, w_eco12828, w_eco12829, w_eco12830, w_eco12831, w_eco12832, w_eco12833, w_eco12834, w_eco12835, w_eco12836, w_eco12837, w_eco12838, w_eco12839, w_eco12840, w_eco12841, w_eco12842, w_eco12843, w_eco12844, w_eco12845, w_eco12846, w_eco12847, w_eco12848, w_eco12849, w_eco12850, w_eco12851, w_eco12852, w_eco12853, w_eco12854, w_eco12855, w_eco12856, w_eco12857, w_eco12858, w_eco12859, w_eco12860, w_eco12861, w_eco12862, w_eco12863, w_eco12864, w_eco12865, w_eco12866, w_eco12867, w_eco12868, w_eco12869, w_eco12870, w_eco12871, w_eco12872, w_eco12873, w_eco12874, w_eco12875, w_eco12876, w_eco12877, w_eco12878, w_eco12879, w_eco12880, w_eco12881, w_eco12882, w_eco12883, w_eco12884, w_eco12885, w_eco12886, w_eco12887, w_eco12888, w_eco12889, w_eco12890, w_eco12891, w_eco12892, w_eco12893, w_eco12894, w_eco12895, w_eco12896, w_eco12897, w_eco12898, w_eco12899, w_eco12900, w_eco12901, w_eco12902, w_eco12903, w_eco12904, w_eco12905, w_eco12906, w_eco12907, w_eco12908, w_eco12909, w_eco12910, w_eco12911, w_eco12912, w_eco12913, w_eco12914, w_eco12915, w_eco12916, w_eco12917, w_eco12918, w_eco12919, w_eco12920, w_eco12921, w_eco12922, w_eco12923, w_eco12924, w_eco12925, w_eco12926, w_eco12927, w_eco12928, w_eco12929, w_eco12930, w_eco12931, w_eco12932, w_eco12933, w_eco12934, w_eco12935, w_eco12936, w_eco12937, w_eco12938, w_eco12939, w_eco12940, w_eco12941, w_eco12942, w_eco12943, w_eco12944, w_eco12945, w_eco12946, w_eco12947, w_eco12948, w_eco12949, w_eco12950, w_eco12951, w_eco12952, w_eco12953, w_eco12954, w_eco12955, w_eco12956, w_eco12957, w_eco12958, w_eco12959, w_eco12960, w_eco12961, w_eco12962, w_eco12963, w_eco12964, w_eco12965, w_eco12966, w_eco12967, w_eco12968, w_eco12969, w_eco12970, w_eco12971, w_eco12972, w_eco12973, w_eco12974, w_eco12975, w_eco12976, w_eco12977, w_eco12978, w_eco12979, w_eco12980, w_eco12981, w_eco12982, w_eco12983, w_eco12984, w_eco12985, w_eco12986, w_eco12987, w_eco12988, w_eco12989, w_eco12990, w_eco12991, w_eco12992, w_eco12993, w_eco12994, w_eco12995, w_eco12996, w_eco12997, w_eco12998, w_eco12999, w_eco13000, w_eco13001, w_eco13002, w_eco13003, w_eco13004, w_eco13005, w_eco13006, w_eco13007, w_eco13008, w_eco13009, w_eco13010, w_eco13011, w_eco13012, w_eco13013, w_eco13014, w_eco13015, w_eco13016, w_eco13017, w_eco13018, w_eco13019, w_eco13020, w_eco13021, w_eco13022, w_eco13023, w_eco13024, w_eco13025, w_eco13026, w_eco13027, w_eco13028, w_eco13029, w_eco13030, w_eco13031, w_eco13032, w_eco13033, w_eco13034, w_eco13035, w_eco13036, w_eco13037, w_eco13038, w_eco13039, w_eco13040, w_eco13041, w_eco13042, w_eco13043, w_eco13044, w_eco13045, w_eco13046, w_eco13047, w_eco13048, w_eco13049, w_eco13050, w_eco13051, w_eco13052, w_eco13053, w_eco13054, w_eco13055, w_eco13056, w_eco13057, w_eco13058, w_eco13059, w_eco13060, w_eco13061, w_eco13062, w_eco13063, w_eco13064, w_eco13065, w_eco13066, w_eco13067, w_eco13068, w_eco13069, w_eco13070, w_eco13071, w_eco13072, w_eco13073, w_eco13074, w_eco13075, w_eco13076, w_eco13077, w_eco13078, w_eco13079, w_eco13080, w_eco13081, w_eco13082, w_eco13083, w_eco13084, w_eco13085, w_eco13086, w_eco13087, w_eco13088, w_eco13089, w_eco13090, w_eco13091, w_eco13092, w_eco13093, w_eco13094, w_eco13095, w_eco13096, w_eco13097, w_eco13098, w_eco13099, w_eco13100, w_eco13101, w_eco13102, w_eco13103, w_eco13104, w_eco13105, w_eco13106, w_eco13107, w_eco13108, w_eco13109, w_eco13110, w_eco13111, w_eco13112, w_eco13113, w_eco13114, w_eco13115, w_eco13116, w_eco13117, w_eco13118, w_eco13119, w_eco13120, w_eco13121, w_eco13122, w_eco13123, w_eco13124, w_eco13125, w_eco13126, w_eco13127, w_eco13128, w_eco13129, w_eco13130, w_eco13131, w_eco13132, w_eco13133, w_eco13134, w_eco13135, w_eco13136, w_eco13137, w_eco13138, w_eco13139, w_eco13140, w_eco13141, w_eco13142, w_eco13143, w_eco13144, w_eco13145, w_eco13146, w_eco13147, w_eco13148, w_eco13149, w_eco13150, w_eco13151, w_eco13152, w_eco13153, w_eco13154, w_eco13155, w_eco13156, w_eco13157, w_eco13158, w_eco13159, w_eco13160, w_eco13161, w_eco13162, w_eco13163, w_eco13164, w_eco13165, w_eco13166, w_eco13167, w_eco13168, w_eco13169, w_eco13170, w_eco13171, w_eco13172, w_eco13173, w_eco13174, w_eco13175, w_eco13176, w_eco13177, w_eco13178, w_eco13179, w_eco13180, w_eco13181, w_eco13182, w_eco13183, w_eco13184, w_eco13185, w_eco13186, w_eco13187, w_eco13188, w_eco13189, w_eco13190, w_eco13191, w_eco13192, w_eco13193, w_eco13194, w_eco13195, w_eco13196, w_eco13197, w_eco13198, w_eco13199, w_eco13200, w_eco13201, w_eco13202, w_eco13203, w_eco13204, w_eco13205, w_eco13206, w_eco13207, w_eco13208, w_eco13209, w_eco13210, sub_wire11, w_eco13211, w_eco13212, w_eco13213, w_eco13214, w_eco13215, w_eco13216, w_eco13217, w_eco13218, w_eco13219, w_eco13220, w_eco13221, w_eco13222, w_eco13223, w_eco13224, w_eco13225, w_eco13226, w_eco13227, w_eco13228, w_eco13229, w_eco13230, w_eco13231, w_eco13232, w_eco13233, w_eco13234, w_eco13235, w_eco13236, w_eco13237, w_eco13238, w_eco13239, w_eco13240, w_eco13241, w_eco13242, w_eco13243, w_eco13244, w_eco13245, w_eco13246, w_eco13247, w_eco13248, w_eco13249, w_eco13250, w_eco13251, w_eco13252, w_eco13253, w_eco13254, w_eco13255, w_eco13256, w_eco13257, w_eco13258, w_eco13259, w_eco13260, w_eco13261, w_eco13262, w_eco13263, w_eco13264, w_eco13265, w_eco13266, w_eco13267, w_eco13268, w_eco13269, w_eco13270, w_eco13271, w_eco13272, w_eco13273, w_eco13274, w_eco13275, w_eco13276, w_eco13277, w_eco13278, w_eco13279, w_eco13280, w_eco13281, w_eco13282, w_eco13283, w_eco13284, w_eco13285, w_eco13286, w_eco13287, w_eco13288, w_eco13289, w_eco13290, w_eco13291, w_eco13292, w_eco13293, w_eco13294, w_eco13295, w_eco13296, w_eco13297, w_eco13298, w_eco13299, w_eco13300, w_eco13301, w_eco13302, w_eco13303, w_eco13304, w_eco13305, w_eco13306, w_eco13307, w_eco13308, w_eco13309, w_eco13310, w_eco13311, w_eco13312, w_eco13313, w_eco13314, w_eco13315, w_eco13316, w_eco13317, w_eco13318, w_eco13319, w_eco13320, w_eco13321, w_eco13322, w_eco13323, w_eco13324, w_eco13325, w_eco13326, w_eco13327, w_eco13328, w_eco13329, w_eco13330, w_eco13331, w_eco13332, w_eco13333, w_eco13334, w_eco13335, w_eco13336, w_eco13337, w_eco13338, w_eco13339, w_eco13340, w_eco13341, w_eco13342, w_eco13343, w_eco13344, w_eco13345, w_eco13346, w_eco13347, w_eco13348, w_eco13349, w_eco13350, w_eco13351, w_eco13352, w_eco13353, w_eco13354, w_eco13355, w_eco13356, w_eco13357, w_eco13358, w_eco13359, w_eco13360, w_eco13361, w_eco13362, w_eco13363, w_eco13364, w_eco13365, w_eco13366, w_eco13367, w_eco13368, w_eco13369, w_eco13370, w_eco13371, w_eco13372, w_eco13373, w_eco13374, w_eco13375, w_eco13376, w_eco13377, w_eco13378, w_eco13379, w_eco13380, w_eco13381, w_eco13382, w_eco13383, w_eco13384, w_eco13385, w_eco13386, w_eco13387, w_eco13388, w_eco13389, w_eco13390, w_eco13391, w_eco13392, w_eco13393, w_eco13394, w_eco13395, w_eco13396, w_eco13397, w_eco13398, w_eco13399, w_eco13400, w_eco13401, w_eco13402, w_eco13403, w_eco13404, w_eco13405, w_eco13406, w_eco13407, w_eco13408, w_eco13409, w_eco13410, w_eco13411, w_eco13412, w_eco13413, w_eco13414, w_eco13415, w_eco13416, w_eco13417, w_eco13418, w_eco13419, w_eco13420, w_eco13421, w_eco13422, w_eco13423, w_eco13424, w_eco13425, w_eco13426, w_eco13427, w_eco13428, w_eco13429, w_eco13430, w_eco13431, w_eco13432, w_eco13433, w_eco13434, w_eco13435, w_eco13436, w_eco13437, w_eco13438, w_eco13439, w_eco13440, w_eco13441, w_eco13442, w_eco13443, w_eco13444, w_eco13445, w_eco13446, w_eco13447, w_eco13448, w_eco13449, w_eco13450, w_eco13451, w_eco13452, w_eco13453, w_eco13454, w_eco13455, w_eco13456, w_eco13457, w_eco13458, w_eco13459, w_eco13460, w_eco13461, w_eco13462, w_eco13463, w_eco13464, w_eco13465, w_eco13466, w_eco13467, w_eco13468, w_eco13469, w_eco13470, w_eco13471, w_eco13472, w_eco13473, w_eco13474, w_eco13475, w_eco13476, w_eco13477, w_eco13478, w_eco13479, w_eco13480, w_eco13481, w_eco13482, w_eco13483, w_eco13484, w_eco13485, w_eco13486, w_eco13487, w_eco13488, w_eco13489, w_eco13490, w_eco13491, w_eco13492, w_eco13493, w_eco13494, w_eco13495, w_eco13496, w_eco13497, w_eco13498, w_eco13499, w_eco13500, w_eco13501, w_eco13502, w_eco13503, w_eco13504, w_eco13505, w_eco13506, w_eco13507, w_eco13508, w_eco13509, w_eco13510, w_eco13511, w_eco13512, w_eco13513, w_eco13514, w_eco13515, w_eco13516, w_eco13517, w_eco13518, w_eco13519, w_eco13520, w_eco13521, w_eco13522, w_eco13523, w_eco13524, w_eco13525, w_eco13526, w_eco13527, w_eco13528, w_eco13529, w_eco13530, w_eco13531, w_eco13532, w_eco13533, w_eco13534, w_eco13535, w_eco13536, w_eco13537, w_eco13538, w_eco13539, w_eco13540, w_eco13541, w_eco13542, w_eco13543, w_eco13544, w_eco13545, w_eco13546, w_eco13547, w_eco13548, w_eco13549, w_eco13550, w_eco13551, w_eco13552, w_eco13553, w_eco13554, w_eco13555, w_eco13556, w_eco13557, w_eco13558, w_eco13559, w_eco13560, w_eco13561, w_eco13562, w_eco13563, w_eco13564, w_eco13565, w_eco13566, w_eco13567, w_eco13568, w_eco13569, w_eco13570, w_eco13571, w_eco13572, w_eco13573, w_eco13574, w_eco13575, w_eco13576, w_eco13577, w_eco13578, w_eco13579, w_eco13580, w_eco13581, w_eco13582, w_eco13583, w_eco13584, w_eco13585, w_eco13586, w_eco13587, w_eco13588, w_eco13589, w_eco13590, w_eco13591, w_eco13592, w_eco13593, w_eco13594, w_eco13595, w_eco13596, w_eco13597, w_eco13598, w_eco13599, w_eco13600, w_eco13601, w_eco13602, w_eco13603, w_eco13604, w_eco13605, w_eco13606, w_eco13607, w_eco13608, w_eco13609, w_eco13610, w_eco13611, w_eco13612, w_eco13613, w_eco13614, w_eco13615, w_eco13616, w_eco13617, w_eco13618, w_eco13619, w_eco13620, w_eco13621, w_eco13622, w_eco13623, w_eco13624, w_eco13625, w_eco13626, w_eco13627, w_eco13628, w_eco13629, w_eco13630, w_eco13631, w_eco13632, w_eco13633, w_eco13634, w_eco13635, w_eco13636, w_eco13637, w_eco13638, w_eco13639, w_eco13640, w_eco13641, w_eco13642, w_eco13643, w_eco13644, w_eco13645, w_eco13646, w_eco13647, w_eco13648, w_eco13649, w_eco13650, w_eco13651, w_eco13652, w_eco13653, w_eco13654, w_eco13655, w_eco13656, w_eco13657, w_eco13658, w_eco13659, w_eco13660, w_eco13661, w_eco13662, w_eco13663, w_eco13664, w_eco13665, w_eco13666, w_eco13667, w_eco13668, w_eco13669, w_eco13670, w_eco13671, w_eco13672, w_eco13673, w_eco13674, w_eco13675, w_eco13676, w_eco13677, w_eco13678, w_eco13679, w_eco13680, w_eco13681, w_eco13682, w_eco13683, w_eco13684, w_eco13685, w_eco13686, w_eco13687, w_eco13688, w_eco13689, w_eco13690, w_eco13691, w_eco13692, w_eco13693, w_eco13694, w_eco13695, w_eco13696, sub_wire12, w_eco13697, w_eco13698, w_eco13699, w_eco13700, w_eco13701, w_eco13702, w_eco13703, w_eco13704, w_eco13705, w_eco13706, w_eco13707, w_eco13708, w_eco13709, w_eco13710, w_eco13711, w_eco13712, w_eco13713, w_eco13714, w_eco13715, w_eco13716, w_eco13717, w_eco13718, w_eco13719, w_eco13720, w_eco13721, w_eco13722, w_eco13723, w_eco13724, w_eco13725, w_eco13726, w_eco13727, w_eco13728, w_eco13729, w_eco13730, w_eco13731, w_eco13732, w_eco13733, w_eco13734, w_eco13735, w_eco13736, w_eco13737, w_eco13738, w_eco13739, w_eco13740, w_eco13741, w_eco13742, w_eco13743, w_eco13744, w_eco13745, w_eco13746, w_eco13747, w_eco13748, w_eco13749, w_eco13750, w_eco13751, w_eco13752, w_eco13753, w_eco13754, w_eco13755, w_eco13756, w_eco13757, w_eco13758, w_eco13759, w_eco13760, w_eco13761, w_eco13762, w_eco13763, w_eco13764, w_eco13765, w_eco13766, w_eco13767, w_eco13768, w_eco13769, w_eco13770, w_eco13771, w_eco13772, w_eco13773, w_eco13774, w_eco13775, w_eco13776, w_eco13777, w_eco13778, w_eco13779, w_eco13780, w_eco13781, w_eco13782, w_eco13783, w_eco13784, w_eco13785, w_eco13786, w_eco13787, w_eco13788, w_eco13789, w_eco13790, w_eco13791, w_eco13792, w_eco13793, w_eco13794, w_eco13795, w_eco13796, w_eco13797, w_eco13798, w_eco13799, w_eco13800, w_eco13801, w_eco13802, w_eco13803, w_eco13804, w_eco13805, w_eco13806, w_eco13807, w_eco13808, w_eco13809, w_eco13810, w_eco13811, w_eco13812, w_eco13813, w_eco13814, w_eco13815, w_eco13816, w_eco13817, w_eco13818, w_eco13819, w_eco13820, w_eco13821, w_eco13822, w_eco13823, w_eco13824, w_eco13825, w_eco13826, w_eco13827, w_eco13828, w_eco13829, w_eco13830, w_eco13831, w_eco13832, w_eco13833, w_eco13834, w_eco13835, w_eco13836, w_eco13837, w_eco13838, w_eco13839, w_eco13840, w_eco13841, w_eco13842, w_eco13843, w_eco13844, w_eco13845, w_eco13846, w_eco13847, w_eco13848, w_eco13849, w_eco13850, w_eco13851, w_eco13852, w_eco13853, w_eco13854, w_eco13855, w_eco13856, w_eco13857, w_eco13858, w_eco13859, w_eco13860, w_eco13861, w_eco13862, w_eco13863, w_eco13864, w_eco13865, w_eco13866, w_eco13867, w_eco13868, w_eco13869, w_eco13870, w_eco13871, w_eco13872, w_eco13873, w_eco13874, w_eco13875, w_eco13876, w_eco13877, w_eco13878, w_eco13879, w_eco13880, w_eco13881, w_eco13882, w_eco13883, w_eco13884, w_eco13885, w_eco13886, w_eco13887, w_eco13888, w_eco13889, w_eco13890, w_eco13891, w_eco13892, w_eco13893, w_eco13894, w_eco13895, w_eco13896, w_eco13897, w_eco13898, w_eco13899, w_eco13900, w_eco13901, w_eco13902, w_eco13903, w_eco13904, w_eco13905, w_eco13906, w_eco13907, w_eco13908, w_eco13909, w_eco13910, w_eco13911, w_eco13912, w_eco13913, w_eco13914, w_eco13915, w_eco13916, w_eco13917, w_eco13918, w_eco13919, w_eco13920, w_eco13921, w_eco13922, w_eco13923, w_eco13924, w_eco13925, w_eco13926, w_eco13927, w_eco13928, w_eco13929, w_eco13930, w_eco13931, w_eco13932, w_eco13933, w_eco13934, w_eco13935, w_eco13936, w_eco13937, w_eco13938, w_eco13939, w_eco13940, w_eco13941, w_eco13942, w_eco13943, w_eco13944, w_eco13945, w_eco13946, w_eco13947, w_eco13948, w_eco13949, w_eco13950, w_eco13951, w_eco13952, w_eco13953, w_eco13954, w_eco13955, w_eco13956, w_eco13957, w_eco13958, w_eco13959, w_eco13960, w_eco13961, w_eco13962, w_eco13963, w_eco13964, w_eco13965, w_eco13966, w_eco13967, w_eco13968, w_eco13969, w_eco13970, w_eco13971, w_eco13972, w_eco13973, w_eco13974, w_eco13975, w_eco13976, w_eco13977, w_eco13978, w_eco13979, w_eco13980, w_eco13981, w_eco13982, w_eco13983, w_eco13984, w_eco13985, w_eco13986, w_eco13987, w_eco13988, w_eco13989, w_eco13990, w_eco13991, w_eco13992, w_eco13993, w_eco13994, w_eco13995, w_eco13996, w_eco13997, w_eco13998, w_eco13999, w_eco14000, w_eco14001, w_eco14002, w_eco14003, w_eco14004, w_eco14005, w_eco14006, w_eco14007, w_eco14008, w_eco14009, w_eco14010, w_eco14011, w_eco14012, w_eco14013, w_eco14014, w_eco14015, w_eco14016, w_eco14017, w_eco14018, w_eco14019, w_eco14020, w_eco14021, w_eco14022, w_eco14023, w_eco14024, w_eco14025, w_eco14026, w_eco14027, w_eco14028, w_eco14029, w_eco14030, w_eco14031, w_eco14032, w_eco14033, w_eco14034, w_eco14035, w_eco14036, w_eco14037, w_eco14038, w_eco14039, w_eco14040, w_eco14041, w_eco14042, w_eco14043, w_eco14044, w_eco14045, w_eco14046, w_eco14047, w_eco14048, w_eco14049, w_eco14050, w_eco14051, w_eco14052, w_eco14053, w_eco14054, w_eco14055, w_eco14056, w_eco14057, w_eco14058, w_eco14059, w_eco14060, w_eco14061, w_eco14062, w_eco14063, w_eco14064, w_eco14065, w_eco14066, w_eco14067, w_eco14068, w_eco14069, w_eco14070, w_eco14071, w_eco14072, w_eco14073, w_eco14074, w_eco14075, w_eco14076, w_eco14077, w_eco14078, w_eco14079, w_eco14080, w_eco14081, w_eco14082, w_eco14083, w_eco14084, w_eco14085, w_eco14086, w_eco14087, w_eco14088, w_eco14089, w_eco14090, w_eco14091, w_eco14092, w_eco14093, w_eco14094, w_eco14095, w_eco14096, w_eco14097, w_eco14098, w_eco14099, w_eco14100, w_eco14101, w_eco14102, w_eco14103, w_eco14104, w_eco14105, w_eco14106, w_eco14107, w_eco14108, w_eco14109, w_eco14110, w_eco14111, w_eco14112, w_eco14113, w_eco14114, w_eco14115, w_eco14116, w_eco14117, w_eco14118, w_eco14119, w_eco14120, w_eco14121, w_eco14122, w_eco14123, w_eco14124, w_eco14125, w_eco14126, w_eco14127, w_eco14128, w_eco14129, w_eco14130, w_eco14131, w_eco14132, w_eco14133, w_eco14134, w_eco14135, w_eco14136, w_eco14137, w_eco14138, w_eco14139, w_eco14140, w_eco14141, w_eco14142, w_eco14143, w_eco14144, w_eco14145, w_eco14146, w_eco14147, w_eco14148, w_eco14149, w_eco14150, w_eco14151, w_eco14152, w_eco14153, w_eco14154, w_eco14155, w_eco14156, w_eco14157, w_eco14158, w_eco14159, w_eco14160, w_eco14161, w_eco14162, w_eco14163, w_eco14164, w_eco14165, w_eco14166, w_eco14167, w_eco14168, w_eco14169, w_eco14170, w_eco14171, w_eco14172, w_eco14173, w_eco14174, w_eco14175, w_eco14176, w_eco14177, w_eco14178, w_eco14179, w_eco14180, w_eco14181, w_eco14182, w_eco14183, w_eco14184, w_eco14185, w_eco14186, w_eco14187, w_eco14188, w_eco14189, w_eco14190, w_eco14191, w_eco14192, w_eco14193, w_eco14194, w_eco14195, w_eco14196, w_eco14197, w_eco14198, w_eco14199, w_eco14200, w_eco14201, w_eco14202, w_eco14203, w_eco14204, w_eco14205, w_eco14206, w_eco14207, w_eco14208, w_eco14209, w_eco14210, w_eco14211, w_eco14212, w_eco14213, w_eco14214, w_eco14215, w_eco14216, w_eco14217, w_eco14218, w_eco14219, w_eco14220, w_eco14221, w_eco14222, w_eco14223, w_eco14224, w_eco14225, w_eco14226, w_eco14227, w_eco14228, w_eco14229, w_eco14230, sub_wire13, w_eco14231, w_eco14232, w_eco14233, w_eco14234, w_eco14235, w_eco14236, w_eco14237, w_eco14238, w_eco14239, w_eco14240, w_eco14241, w_eco14242, w_eco14243, w_eco14244, w_eco14245, w_eco14246, w_eco14247, w_eco14248, w_eco14249, w_eco14250, w_eco14251, w_eco14252, w_eco14253, w_eco14254, w_eco14255, w_eco14256, w_eco14257, w_eco14258, w_eco14259, w_eco14260, w_eco14261, w_eco14262, w_eco14263, w_eco14264, w_eco14265, w_eco14266, w_eco14267, w_eco14268, w_eco14269, w_eco14270, w_eco14271, w_eco14272, w_eco14273, w_eco14274, w_eco14275, w_eco14276, w_eco14277, w_eco14278, w_eco14279, w_eco14280, w_eco14281, w_eco14282, w_eco14283, w_eco14284, w_eco14285, w_eco14286, w_eco14287, w_eco14288, w_eco14289, w_eco14290, w_eco14291, w_eco14292, w_eco14293, w_eco14294, w_eco14295, w_eco14296, w_eco14297, w_eco14298, w_eco14299, w_eco14300, w_eco14301, w_eco14302, w_eco14303, w_eco14304, w_eco14305, w_eco14306, w_eco14307, w_eco14308, w_eco14309, w_eco14310, w_eco14311, w_eco14312, w_eco14313, w_eco14314, w_eco14315, w_eco14316, w_eco14317, w_eco14318, w_eco14319, w_eco14320, w_eco14321, w_eco14322, w_eco14323, w_eco14324, w_eco14325, w_eco14326, w_eco14327, w_eco14328, w_eco14329, w_eco14330, w_eco14331, w_eco14332, w_eco14333, w_eco14334, w_eco14335, w_eco14336, w_eco14337, w_eco14338, w_eco14339, w_eco14340, w_eco14341, w_eco14342, w_eco14343, w_eco14344, w_eco14345, w_eco14346, w_eco14347, w_eco14348, w_eco14349, w_eco14350, w_eco14351, w_eco14352, w_eco14353, w_eco14354, w_eco14355, w_eco14356, w_eco14357, w_eco14358, w_eco14359, w_eco14360, w_eco14361, w_eco14362, w_eco14363, w_eco14364, w_eco14365, w_eco14366, w_eco14367, w_eco14368, w_eco14369, w_eco14370, w_eco14371, w_eco14372, w_eco14373, w_eco14374, w_eco14375, w_eco14376, w_eco14377, w_eco14378, w_eco14379, w_eco14380, w_eco14381, w_eco14382, w_eco14383, w_eco14384, w_eco14385, w_eco14386, w_eco14387, w_eco14388, w_eco14389, w_eco14390, w_eco14391, w_eco14392, w_eco14393, w_eco14394, w_eco14395, w_eco14396, w_eco14397, w_eco14398, w_eco14399, w_eco14400, w_eco14401, w_eco14402, w_eco14403, w_eco14404, w_eco14405, w_eco14406, w_eco14407, w_eco14408, w_eco14409, w_eco14410, w_eco14411, w_eco14412, w_eco14413, w_eco14414, w_eco14415, w_eco14416, w_eco14417, w_eco14418, w_eco14419, w_eco14420, w_eco14421, w_eco14422, w_eco14423, w_eco14424, w_eco14425, w_eco14426, w_eco14427, w_eco14428, w_eco14429, w_eco14430, w_eco14431, w_eco14432, w_eco14433, w_eco14434, w_eco14435, w_eco14436, w_eco14437, w_eco14438, w_eco14439, w_eco14440, w_eco14441, w_eco14442, w_eco14443, w_eco14444, w_eco14445, w_eco14446, w_eco14447, w_eco14448, w_eco14449, w_eco14450, w_eco14451, w_eco14452, w_eco14453, w_eco14454, w_eco14455, w_eco14456, w_eco14457, w_eco14458, w_eco14459, w_eco14460, w_eco14461, w_eco14462, w_eco14463, w_eco14464, w_eco14465, w_eco14466, w_eco14467, w_eco14468, w_eco14469, w_eco14470, w_eco14471, w_eco14472, w_eco14473, w_eco14474, w_eco14475, w_eco14476, w_eco14477, w_eco14478, w_eco14479, w_eco14480, w_eco14481, w_eco14482, w_eco14483, w_eco14484, w_eco14485, w_eco14486, w_eco14487, w_eco14488, w_eco14489, w_eco14490, w_eco14491, w_eco14492, w_eco14493, w_eco14494, w_eco14495, w_eco14496, w_eco14497, w_eco14498, w_eco14499, w_eco14500, w_eco14501, w_eco14502, w_eco14503, w_eco14504, w_eco14505, w_eco14506, w_eco14507, w_eco14508, w_eco14509, w_eco14510, w_eco14511, w_eco14512, w_eco14513, w_eco14514, w_eco14515, w_eco14516, w_eco14517, w_eco14518, w_eco14519, w_eco14520, w_eco14521, w_eco14522, w_eco14523, w_eco14524, w_eco14525, w_eco14526, w_eco14527, w_eco14528, w_eco14529, w_eco14530, w_eco14531, w_eco14532, w_eco14533, w_eco14534, w_eco14535, w_eco14536, w_eco14537, w_eco14538, w_eco14539, w_eco14540, w_eco14541, w_eco14542, w_eco14543, w_eco14544, w_eco14545, w_eco14546, w_eco14547, w_eco14548, w_eco14549, w_eco14550, w_eco14551, w_eco14552, w_eco14553, w_eco14554, w_eco14555, w_eco14556, w_eco14557, w_eco14558, w_eco14559, w_eco14560, w_eco14561, w_eco14562, w_eco14563, sub_wire14, w_eco14564, w_eco14565, w_eco14566, w_eco14567, w_eco14568, w_eco14569, w_eco14570, w_eco14571, w_eco14572, w_eco14573, w_eco14574, w_eco14575, w_eco14576, w_eco14577, w_eco14578, w_eco14579, w_eco14580, w_eco14581, w_eco14582, w_eco14583, w_eco14584, w_eco14585, w_eco14586, w_eco14587, w_eco14588, w_eco14589, w_eco14590, w_eco14591, w_eco14592, w_eco14593, w_eco14594, w_eco14595, w_eco14596, w_eco14597, w_eco14598, w_eco14599, w_eco14600, w_eco14601, w_eco14602, w_eco14603, w_eco14604, w_eco14605, w_eco14606, w_eco14607, w_eco14608, w_eco14609, w_eco14610, w_eco14611, w_eco14612, w_eco14613, w_eco14614, w_eco14615, w_eco14616, w_eco14617, w_eco14618, w_eco14619, w_eco14620, w_eco14621, w_eco14622, w_eco14623, w_eco14624, w_eco14625, w_eco14626, w_eco14627, w_eco14628, w_eco14629, w_eco14630, w_eco14631, w_eco14632, w_eco14633, w_eco14634, w_eco14635, w_eco14636, w_eco14637, w_eco14638, w_eco14639, w_eco14640, w_eco14641, w_eco14642, w_eco14643, w_eco14644, w_eco14645, w_eco14646, w_eco14647, w_eco14648, w_eco14649, w_eco14650, w_eco14651, w_eco14652, w_eco14653, w_eco14654, w_eco14655, w_eco14656, w_eco14657, w_eco14658, w_eco14659, w_eco14660, w_eco14661, w_eco14662, w_eco14663, w_eco14664, w_eco14665, w_eco14666, w_eco14667, w_eco14668, w_eco14669, w_eco14670, w_eco14671, w_eco14672, w_eco14673, w_eco14674, w_eco14675, w_eco14676, w_eco14677, w_eco14678, w_eco14679, w_eco14680, w_eco14681, w_eco14682, w_eco14683, w_eco14684, w_eco14685, w_eco14686, w_eco14687, w_eco14688, w_eco14689, w_eco14690, w_eco14691, w_eco14692, w_eco14693, w_eco14694, w_eco14695, w_eco14696, w_eco14697, w_eco14698, w_eco14699, w_eco14700, w_eco14701, w_eco14702, w_eco14703, w_eco14704, w_eco14705, w_eco14706, w_eco14707, w_eco14708, w_eco14709, w_eco14710, w_eco14711, w_eco14712, w_eco14713, w_eco14714, w_eco14715, w_eco14716, w_eco14717, w_eco14718, w_eco14719, w_eco14720, w_eco14721, w_eco14722, w_eco14723, w_eco14724, w_eco14725, w_eco14726, w_eco14727, w_eco14728, w_eco14729, w_eco14730, w_eco14731, w_eco14732, w_eco14733, w_eco14734, w_eco14735, w_eco14736, w_eco14737, w_eco14738, w_eco14739, w_eco14740, w_eco14741, w_eco14742, w_eco14743, w_eco14744, w_eco14745, w_eco14746, w_eco14747, w_eco14748, w_eco14749, w_eco14750, w_eco14751, w_eco14752, w_eco14753, w_eco14754, w_eco14755, w_eco14756, w_eco14757, w_eco14758, w_eco14759, w_eco14760, w_eco14761, w_eco14762, w_eco14763, w_eco14764, w_eco14765, w_eco14766, w_eco14767, w_eco14768, w_eco14769, w_eco14770, w_eco14771, w_eco14772, w_eco14773, w_eco14774, w_eco14775, w_eco14776, w_eco14777, w_eco14778, w_eco14779, w_eco14780, w_eco14781, w_eco14782, w_eco14783, w_eco14784, w_eco14785, w_eco14786, w_eco14787, w_eco14788, w_eco14789, w_eco14790, w_eco14791, w_eco14792, w_eco14793, w_eco14794, w_eco14795, w_eco14796, w_eco14797, w_eco14798, w_eco14799, w_eco14800, w_eco14801, w_eco14802, w_eco14803, w_eco14804, w_eco14805, w_eco14806, w_eco14807, w_eco14808, w_eco14809, w_eco14810, w_eco14811, w_eco14812, w_eco14813, w_eco14814, w_eco14815, w_eco14816, w_eco14817, w_eco14818, w_eco14819, w_eco14820, w_eco14821, w_eco14822, w_eco14823, w_eco14824, w_eco14825, w_eco14826, w_eco14827, w_eco14828, w_eco14829, w_eco14830, w_eco14831, w_eco14832, w_eco14833, w_eco14834, w_eco14835, w_eco14836, w_eco14837, w_eco14838, w_eco14839, w_eco14840, w_eco14841, w_eco14842, w_eco14843, w_eco14844, w_eco14845, w_eco14846, w_eco14847, sub_wire15, w_eco14848, w_eco14849, w_eco14850, w_eco14851, w_eco14852, w_eco14853, w_eco14854, w_eco14855, w_eco14856, w_eco14857, w_eco14858, w_eco14859, w_eco14860, w_eco14861, w_eco14862, w_eco14863, w_eco14864, w_eco14865, w_eco14866, w_eco14867, w_eco14868, w_eco14869, w_eco14870, w_eco14871, w_eco14872, w_eco14873, w_eco14874, w_eco14875, w_eco14876, w_eco14877, w_eco14878, w_eco14879, w_eco14880, w_eco14881, w_eco14882, w_eco14883, w_eco14884, w_eco14885, w_eco14886, w_eco14887, w_eco14888, w_eco14889, w_eco14890, w_eco14891, w_eco14892, w_eco14893, w_eco14894, w_eco14895, w_eco14896, w_eco14897, w_eco14898, w_eco14899, w_eco14900, w_eco14901, w_eco14902, w_eco14903, w_eco14904, w_eco14905, w_eco14906, w_eco14907, w_eco14908, w_eco14909, w_eco14910, w_eco14911, w_eco14912, w_eco14913, w_eco14914, w_eco14915, w_eco14916, w_eco14917, w_eco14918, w_eco14919, w_eco14920, w_eco14921, w_eco14922, w_eco14923, w_eco14924, w_eco14925, w_eco14926, w_eco14927, w_eco14928, w_eco14929, w_eco14930, w_eco14931, w_eco14932, w_eco14933, w_eco14934, w_eco14935, w_eco14936, w_eco14937, w_eco14938, w_eco14939, w_eco14940, w_eco14941, w_eco14942, w_eco14943, w_eco14944, w_eco14945, w_eco14946, w_eco14947, w_eco14948, w_eco14949, w_eco14950, w_eco14951, w_eco14952, w_eco14953, w_eco14954, w_eco14955, w_eco14956, w_eco14957, w_eco14958, w_eco14959, w_eco14960, w_eco14961, w_eco14962, w_eco14963, w_eco14964, w_eco14965, w_eco14966, w_eco14967, w_eco14968, w_eco14969, w_eco14970, w_eco14971, w_eco14972, w_eco14973, w_eco14974, w_eco14975, w_eco14976, w_eco14977, w_eco14978, w_eco14979, w_eco14980, w_eco14981, w_eco14982, w_eco14983, w_eco14984, w_eco14985, w_eco14986, w_eco14987, w_eco14988, w_eco14989, w_eco14990, w_eco14991, w_eco14992, w_eco14993, w_eco14994, w_eco14995, w_eco14996, w_eco14997, w_eco14998, w_eco14999, w_eco15000, w_eco15001, w_eco15002, w_eco15003, w_eco15004, w_eco15005, w_eco15006, w_eco15007, w_eco15008, w_eco15009, w_eco15010, w_eco15011, w_eco15012, w_eco15013, w_eco15014, w_eco15015, w_eco15016, w_eco15017, w_eco15018, w_eco15019, w_eco15020, w_eco15021, w_eco15022, w_eco15023, w_eco15024, w_eco15025, w_eco15026, w_eco15027, w_eco15028, w_eco15029, w_eco15030, w_eco15031, w_eco15032, w_eco15033, w_eco15034, w_eco15035, w_eco15036, w_eco15037, w_eco15038, w_eco15039, w_eco15040, w_eco15041, w_eco15042, w_eco15043, w_eco15044, w_eco15045, w_eco15046, w_eco15047, w_eco15048, w_eco15049, w_eco15050, w_eco15051, w_eco15052, w_eco15053, w_eco15054, w_eco15055, w_eco15056, w_eco15057, w_eco15058, w_eco15059, w_eco15060, w_eco15061, w_eco15062, w_eco15063, w_eco15064, w_eco15065, w_eco15066, w_eco15067, w_eco15068, w_eco15069, w_eco15070, w_eco15071, w_eco15072, w_eco15073, w_eco15074, w_eco15075, w_eco15076, w_eco15077, w_eco15078, w_eco15079, w_eco15080, w_eco15081, w_eco15082, w_eco15083, w_eco15084, w_eco15085, w_eco15086, w_eco15087, w_eco15088, w_eco15089, w_eco15090, w_eco15091, w_eco15092, w_eco15093, w_eco15094, w_eco15095, w_eco15096, w_eco15097, w_eco15098, w_eco15099, w_eco15100, w_eco15101, w_eco15102, w_eco15103, w_eco15104, w_eco15105, w_eco15106, w_eco15107, w_eco15108, w_eco15109, w_eco15110, w_eco15111, w_eco15112, w_eco15113, w_eco15114, w_eco15115, w_eco15116, w_eco15117, w_eco15118, w_eco15119, w_eco15120, w_eco15121, w_eco15122, w_eco15123, w_eco15124, w_eco15125, w_eco15126, w_eco15127, w_eco15128, w_eco15129, w_eco15130, w_eco15131, w_eco15132, w_eco15133, w_eco15134, w_eco15135, w_eco15136, w_eco15137, w_eco15138, w_eco15139, w_eco15140, w_eco15141, w_eco15142, w_eco15143, w_eco15144, w_eco15145, w_eco15146, w_eco15147, w_eco15148, w_eco15149, w_eco15150, w_eco15151, w_eco15152, w_eco15153, w_eco15154, w_eco15155, w_eco15156, sub_wire16, w_eco15157, w_eco15158, w_eco15159, w_eco15160, w_eco15161, w_eco15162, w_eco15163, w_eco15164, w_eco15165, w_eco15166, w_eco15167, w_eco15168, w_eco15169, w_eco15170, w_eco15171, w_eco15172, w_eco15173, w_eco15174, w_eco15175, w_eco15176, w_eco15177, w_eco15178, w_eco15179, w_eco15180, w_eco15181, w_eco15182, w_eco15183, w_eco15184, w_eco15185, w_eco15186, w_eco15187, w_eco15188, w_eco15189, w_eco15190, w_eco15191, w_eco15192, w_eco15193, w_eco15194, w_eco15195, w_eco15196, w_eco15197, w_eco15198, w_eco15199, w_eco15200, w_eco15201, w_eco15202, w_eco15203, w_eco15204, w_eco15205, w_eco15206, w_eco15207, w_eco15208, w_eco15209, w_eco15210, w_eco15211, w_eco15212, w_eco15213, w_eco15214, w_eco15215, w_eco15216, w_eco15217, w_eco15218, w_eco15219, w_eco15220, w_eco15221, w_eco15222, w_eco15223, w_eco15224, w_eco15225, w_eco15226, w_eco15227, w_eco15228, w_eco15229, w_eco15230, w_eco15231, w_eco15232, w_eco15233, w_eco15234, w_eco15235, w_eco15236, w_eco15237, w_eco15238, w_eco15239, w_eco15240, w_eco15241, w_eco15242, w_eco15243, w_eco15244, w_eco15245, w_eco15246, w_eco15247, w_eco15248, w_eco15249, w_eco15250, w_eco15251, w_eco15252, w_eco15253, w_eco15254, w_eco15255, w_eco15256, w_eco15257, w_eco15258, w_eco15259, w_eco15260, w_eco15261, w_eco15262, w_eco15263, w_eco15264, w_eco15265, w_eco15266, w_eco15267, w_eco15268, w_eco15269, w_eco15270, w_eco15271, w_eco15272, w_eco15273, w_eco15274, w_eco15275, w_eco15276, w_eco15277, w_eco15278, w_eco15279, w_eco15280, w_eco15281, w_eco15282, w_eco15283, w_eco15284, w_eco15285, w_eco15286, w_eco15287, w_eco15288, w_eco15289, w_eco15290, w_eco15291, w_eco15292, w_eco15293, w_eco15294, w_eco15295, w_eco15296, w_eco15297, w_eco15298, w_eco15299, w_eco15300, w_eco15301, w_eco15302, w_eco15303, w_eco15304, w_eco15305, w_eco15306, w_eco15307, w_eco15308, w_eco15309, w_eco15310, w_eco15311, w_eco15312, w_eco15313, w_eco15314, w_eco15315, w_eco15316, w_eco15317, w_eco15318, w_eco15319, w_eco15320, w_eco15321, w_eco15322, w_eco15323, w_eco15324, w_eco15325, w_eco15326, w_eco15327, w_eco15328, w_eco15329, w_eco15330, w_eco15331, w_eco15332, w_eco15333, w_eco15334, w_eco15335, w_eco15336, w_eco15337, w_eco15338, w_eco15339, w_eco15340, w_eco15341, w_eco15342, w_eco15343, w_eco15344, w_eco15345, w_eco15346, w_eco15347, w_eco15348, w_eco15349, w_eco15350, w_eco15351, w_eco15352, w_eco15353, w_eco15354, w_eco15355, w_eco15356, w_eco15357, w_eco15358, w_eco15359, w_eco15360, w_eco15361, w_eco15362, w_eco15363, w_eco15364, w_eco15365, w_eco15366, w_eco15367, w_eco15368, w_eco15369, w_eco15370, w_eco15371, w_eco15372, w_eco15373, w_eco15374, w_eco15375, w_eco15376, w_eco15377, w_eco15378, w_eco15379, w_eco15380, w_eco15381, w_eco15382, w_eco15383, w_eco15384, w_eco15385, w_eco15386, w_eco15387, w_eco15388, w_eco15389, w_eco15390, w_eco15391, w_eco15392, w_eco15393, w_eco15394, w_eco15395, w_eco15396, w_eco15397, w_eco15398, w_eco15399, w_eco15400, w_eco15401, w_eco15402, w_eco15403, w_eco15404, w_eco15405, w_eco15406, w_eco15407, w_eco15408, w_eco15409, w_eco15410, w_eco15411, w_eco15412, w_eco15413, w_eco15414, w_eco15415, w_eco15416, w_eco15417, w_eco15418, w_eco15419, w_eco15420, w_eco15421, w_eco15422, w_eco15423, w_eco15424, w_eco15425, w_eco15426, w_eco15427, w_eco15428, w_eco15429, w_eco15430, w_eco15431, w_eco15432, w_eco15433, w_eco15434, w_eco15435, w_eco15436, w_eco15437, w_eco15438, w_eco15439, w_eco15440, w_eco15441, w_eco15442, w_eco15443, w_eco15444, w_eco15445, w_eco15446, w_eco15447, w_eco15448, w_eco15449, w_eco15450, w_eco15451, w_eco15452, w_eco15453, w_eco15454, w_eco15455, w_eco15456, w_eco15457, w_eco15458, w_eco15459, w_eco15460, w_eco15461, w_eco15462, w_eco15463, w_eco15464, w_eco15465, w_eco15466, w_eco15467, w_eco15468, w_eco15469, w_eco15470, w_eco15471, w_eco15472, w_eco15473, w_eco15474, w_eco15475, w_eco15476, w_eco15477, w_eco15478, w_eco15479, w_eco15480, w_eco15481, w_eco15482, w_eco15483, sub_wire17, w_eco15484, w_eco15485, w_eco15486, w_eco15487, w_eco15488, w_eco15489, w_eco15490, w_eco15491, w_eco15492, w_eco15493, w_eco15494, w_eco15495, w_eco15496, w_eco15497, w_eco15498, w_eco15499, w_eco15500, w_eco15501, w_eco15502, w_eco15503, w_eco15504, w_eco15505, w_eco15506, w_eco15507, w_eco15508, w_eco15509, w_eco15510, w_eco15511, w_eco15512, w_eco15513, w_eco15514, w_eco15515, w_eco15516, w_eco15517, w_eco15518, w_eco15519, w_eco15520, w_eco15521, w_eco15522, w_eco15523, w_eco15524, w_eco15525, w_eco15526, w_eco15527, w_eco15528, w_eco15529, w_eco15530, w_eco15531, w_eco15532, w_eco15533, w_eco15534, w_eco15535, w_eco15536, w_eco15537, w_eco15538, w_eco15539, w_eco15540, w_eco15541, w_eco15542, w_eco15543, w_eco15544, w_eco15545, w_eco15546, w_eco15547, w_eco15548, w_eco15549, w_eco15550, w_eco15551, w_eco15552, w_eco15553, w_eco15554, w_eco15555, w_eco15556, w_eco15557, w_eco15558, w_eco15559, w_eco15560, w_eco15561, w_eco15562, w_eco15563, w_eco15564, w_eco15565, w_eco15566, w_eco15567, w_eco15568, w_eco15569, w_eco15570, w_eco15571, w_eco15572, w_eco15573, w_eco15574, w_eco15575, w_eco15576, w_eco15577, w_eco15578, w_eco15579, w_eco15580, w_eco15581, w_eco15582, w_eco15583, w_eco15584, w_eco15585, w_eco15586, w_eco15587, w_eco15588, w_eco15589, w_eco15590, w_eco15591, w_eco15592, w_eco15593, w_eco15594, w_eco15595, w_eco15596, w_eco15597, w_eco15598, w_eco15599, w_eco15600, w_eco15601, w_eco15602, w_eco15603, w_eco15604, w_eco15605, w_eco15606, w_eco15607, w_eco15608, w_eco15609, w_eco15610, w_eco15611, w_eco15612, w_eco15613, w_eco15614, w_eco15615, w_eco15616, w_eco15617, w_eco15618, w_eco15619, w_eco15620, w_eco15621, w_eco15622, w_eco15623, w_eco15624, w_eco15625, w_eco15626, w_eco15627, w_eco15628, w_eco15629, w_eco15630, w_eco15631, w_eco15632, w_eco15633, w_eco15634, w_eco15635, w_eco15636, w_eco15637, w_eco15638, w_eco15639, w_eco15640, w_eco15641, w_eco15642, w_eco15643, w_eco15644, w_eco15645, w_eco15646, w_eco15647, w_eco15648, w_eco15649, w_eco15650, w_eco15651, w_eco15652, w_eco15653, w_eco15654, w_eco15655, w_eco15656, w_eco15657, w_eco15658, w_eco15659, w_eco15660, w_eco15661, w_eco15662, w_eco15663, w_eco15664, w_eco15665, w_eco15666, w_eco15667, w_eco15668, w_eco15669, w_eco15670, w_eco15671, w_eco15672, w_eco15673, w_eco15674, w_eco15675, w_eco15676, w_eco15677, w_eco15678, w_eco15679, w_eco15680, w_eco15681, w_eco15682, w_eco15683, w_eco15684, w_eco15685, w_eco15686, w_eco15687, w_eco15688, w_eco15689, w_eco15690, w_eco15691, w_eco15692, w_eco15693, w_eco15694, w_eco15695, w_eco15696, w_eco15697, w_eco15698, w_eco15699, w_eco15700, w_eco15701, w_eco15702, w_eco15703, w_eco15704, w_eco15705, w_eco15706, w_eco15707, w_eco15708, w_eco15709, w_eco15710, w_eco15711, w_eco15712, w_eco15713, w_eco15714, w_eco15715, w_eco15716, w_eco15717, w_eco15718, w_eco15719, w_eco15720, w_eco15721, w_eco15722, w_eco15723, w_eco15724, w_eco15725, w_eco15726, w_eco15727, w_eco15728, w_eco15729, w_eco15730, w_eco15731, w_eco15732, w_eco15733, w_eco15734, w_eco15735, w_eco15736, w_eco15737, w_eco15738, w_eco15739, w_eco15740, w_eco15741, w_eco15742, w_eco15743, w_eco15744, w_eco15745, w_eco15746, w_eco15747, w_eco15748, w_eco15749, w_eco15750, w_eco15751, w_eco15752, w_eco15753, w_eco15754, w_eco15755, w_eco15756, w_eco15757, w_eco15758, w_eco15759, w_eco15760, w_eco15761, w_eco15762, w_eco15763, w_eco15764, w_eco15765, w_eco15766, w_eco15767, w_eco15768, w_eco15769, w_eco15770, w_eco15771, w_eco15772, w_eco15773, w_eco15774, w_eco15775, w_eco15776, w_eco15777, w_eco15778, w_eco15779, w_eco15780, w_eco15781, w_eco15782, w_eco15783, w_eco15784, w_eco15785, w_eco15786, w_eco15787, w_eco15788, w_eco15789, w_eco15790, w_eco15791, w_eco15792, w_eco15793, w_eco15794, w_eco15795, w_eco15796, w_eco15797, w_eco15798, w_eco15799, w_eco15800, w_eco15801, w_eco15802, w_eco15803, w_eco15804, w_eco15805, w_eco15806, w_eco15807, w_eco15808, w_eco15809, w_eco15810, w_eco15811, w_eco15812, w_eco15813, w_eco15814, w_eco15815, w_eco15816, w_eco15817, w_eco15818, w_eco15819, w_eco15820, w_eco15821, w_eco15822, w_eco15823, w_eco15824, w_eco15825, w_eco15826, w_eco15827, w_eco15828, sub_wire18, w_eco15829, w_eco15830, w_eco15831, w_eco15832, w_eco15833, w_eco15834, w_eco15835, w_eco15836, w_eco15837, w_eco15838, w_eco15839, w_eco15840, w_eco15841, w_eco15842, w_eco15843, w_eco15844, w_eco15845, w_eco15846, w_eco15847, w_eco15848, w_eco15849, w_eco15850, w_eco15851, w_eco15852, w_eco15853, w_eco15854, w_eco15855, w_eco15856, w_eco15857, w_eco15858, w_eco15859, w_eco15860, w_eco15861, w_eco15862, w_eco15863, w_eco15864, w_eco15865, w_eco15866, w_eco15867, w_eco15868, w_eco15869, w_eco15870, w_eco15871, w_eco15872, w_eco15873, w_eco15874, w_eco15875, w_eco15876, w_eco15877, w_eco15878, w_eco15879, w_eco15880, w_eco15881, w_eco15882, w_eco15883, w_eco15884, w_eco15885, w_eco15886, w_eco15887, w_eco15888, w_eco15889, w_eco15890, w_eco15891, w_eco15892, w_eco15893, w_eco15894, w_eco15895, w_eco15896, w_eco15897, w_eco15898, w_eco15899, w_eco15900, w_eco15901, w_eco15902, w_eco15903, w_eco15904, w_eco15905, w_eco15906, w_eco15907, w_eco15908, w_eco15909, w_eco15910, w_eco15911, w_eco15912, w_eco15913, w_eco15914, w_eco15915, w_eco15916, w_eco15917, w_eco15918, w_eco15919, w_eco15920, w_eco15921, w_eco15922, w_eco15923, w_eco15924, w_eco15925, w_eco15926, w_eco15927, w_eco15928, w_eco15929, w_eco15930, w_eco15931, w_eco15932, w_eco15933, w_eco15934, w_eco15935, w_eco15936, w_eco15937, w_eco15938, w_eco15939, w_eco15940, w_eco15941, w_eco15942, w_eco15943, w_eco15944, w_eco15945, w_eco15946, w_eco15947, w_eco15948, w_eco15949, w_eco15950, w_eco15951, w_eco15952, w_eco15953, w_eco15954, w_eco15955, w_eco15956, w_eco15957, w_eco15958, w_eco15959, w_eco15960, w_eco15961, w_eco15962, w_eco15963, w_eco15964, w_eco15965, w_eco15966, w_eco15967, w_eco15968, w_eco15969, w_eco15970, w_eco15971, w_eco15972, w_eco15973, w_eco15974;

	assign \mux_cnt_122_11_g657/data0 = 0;
	assign \mux_cnt_122_11_g661/data0 = 0;
	assign \mux_cnt_122_11_g665/data0 = 0;
	assign \mux_cnt_122_11_g669/data0 = 0;
	assign \mux_cnt_122_11_g673/data0 = 0;
	assign \mux_cnt_122_11_g677/data0 = 0;
	assign \mux_cnt_122_11_g681/data0 = 0;
	assign \mux_cnt_122_11_g713/data0 = 0;
	assign \mux_cnt_122_11_g653/data0 = 0;
	assign \mux_cnt_122_11_g685/data0 = 0;
	assign \mux_cnt_122_11_g689/data0 = 0;
	assign \mux_cnt_122_11_g693/data0 = 0;
	assign \mux_cnt_122_11_g697/data0 = 0;
	assign \mux_cnt_122_11_g701/data0 = 0;
	assign \mux_cnt_122_11_g705/data0 = 0;
	assign \mux_cnt_122_11_g709/data0 = 0;
	or \mux_cnt_122_11_g657/org(sub_wire0, \mux_cnt_122_11_g657/w_0, \mux_cnt_122_11_g657/w_1, \mux_cnt_122_11_g657/w_2, \mux_cnt_122_11_g657/w_3, \mux_cnt_122_11_g657/w_4);
	and \mux_cnt_122_11_g657/a_4(\mux_cnt_122_11_g657/w_4, Gate, Tgate[6]);
	and \mux_cnt_122_11_g657/a_3(\mux_cnt_122_11_g657/w_3, n_326, Tgdel[6]);
	and \mux_cnt_122_11_g657/a_2(\mux_cnt_122_11_g657/w_2, n_746, cnt_nxt[6]);
	and \mux_cnt_122_11_g657/a_1(\mux_cnt_122_11_g657/w_1, Sync, Tsync[6]);
	and \mux_cnt_122_11_g657/a_0(\mux_cnt_122_11_g657/w_0, n_744, \mux_cnt_122_11_g657/data0);
	or \mux_cnt_122_11_g661/org(sub_wire3, \mux_cnt_122_11_g661/w_0, \mux_cnt_122_11_g661/w_1, \mux_cnt_122_11_g661/w_2, \mux_cnt_122_11_g661/w_3, \mux_cnt_122_11_g661/w_4);
	and \mux_cnt_122_11_g661/a_4(\mux_cnt_122_11_g661/w_4, Gate, Tgate[5]);
	and \mux_cnt_122_11_g661/a_3(\mux_cnt_122_11_g661/w_3, n_326, Tgdel[5]);
	and \mux_cnt_122_11_g661/a_2(\mux_cnt_122_11_g661/w_2, n_746, cnt_nxt[5]);
	and \mux_cnt_122_11_g661/a_1(\mux_cnt_122_11_g661/w_1, Sync, Tsync[5]);
	and \mux_cnt_122_11_g661/a_0(\mux_cnt_122_11_g661/w_0, n_744, \mux_cnt_122_11_g661/data0);
	or \mux_cnt_122_11_g665/org(sub_wire4, \mux_cnt_122_11_g665/w_0, \mux_cnt_122_11_g665/w_1, \mux_cnt_122_11_g665/w_2, \mux_cnt_122_11_g665/w_3, \mux_cnt_122_11_g665/w_4);
	and \mux_cnt_122_11_g665/a_4(\mux_cnt_122_11_g665/w_4, Gate, Tgate[4]);
	and \mux_cnt_122_11_g665/a_3(\mux_cnt_122_11_g665/w_3, n_326, Tgdel[4]);
	and \mux_cnt_122_11_g665/a_2(\mux_cnt_122_11_g665/w_2, n_746, cnt_nxt[4]);
	and \mux_cnt_122_11_g665/a_1(\mux_cnt_122_11_g665/w_1, Sync, Tsync[4]);
	and \mux_cnt_122_11_g665/a_0(\mux_cnt_122_11_g665/w_0, n_744, \mux_cnt_122_11_g665/data0);
	or \mux_cnt_122_11_g669/org(sub_wire5, \mux_cnt_122_11_g669/w_0, \mux_cnt_122_11_g669/w_1, \mux_cnt_122_11_g669/w_2, \mux_cnt_122_11_g669/w_3, \mux_cnt_122_11_g669/w_4);
	and \mux_cnt_122_11_g669/a_4(\mux_cnt_122_11_g669/w_4, Gate, Tgate[3]);
	and \mux_cnt_122_11_g669/a_3(\mux_cnt_122_11_g669/w_3, n_326, Tgdel[3]);
	and \mux_cnt_122_11_g669/a_2(\mux_cnt_122_11_g669/w_2, n_746, cnt_nxt[3]);
	and \mux_cnt_122_11_g669/a_1(\mux_cnt_122_11_g669/w_1, Sync, Tsync[3]);
	and \mux_cnt_122_11_g669/a_0(\mux_cnt_122_11_g669/w_0, n_744, \mux_cnt_122_11_g669/data0);
	or \mux_cnt_122_11_g673/org(sub_wire6, \mux_cnt_122_11_g673/w_0, \mux_cnt_122_11_g673/w_1, \mux_cnt_122_11_g673/w_2, \mux_cnt_122_11_g673/w_3, \mux_cnt_122_11_g673/w_4);
	and \mux_cnt_122_11_g673/a_4(\mux_cnt_122_11_g673/w_4, Gate, Tgate[2]);
	and \mux_cnt_122_11_g673/a_3(\mux_cnt_122_11_g673/w_3, n_326, Tgdel[2]);
	and \mux_cnt_122_11_g673/a_2(\mux_cnt_122_11_g673/w_2, n_746, cnt_nxt[2]);
	and \mux_cnt_122_11_g673/a_1(\mux_cnt_122_11_g673/w_1, Sync, Tsync[2]);
	and \mux_cnt_122_11_g673/a_0(\mux_cnt_122_11_g673/w_0, n_744, \mux_cnt_122_11_g673/data0);
	or \mux_cnt_122_11_g677/org(sub_wire7, \mux_cnt_122_11_g677/w_0, \mux_cnt_122_11_g677/w_1, \mux_cnt_122_11_g677/w_2, \mux_cnt_122_11_g677/w_3, \mux_cnt_122_11_g677/w_4);
	and \mux_cnt_122_11_g677/a_4(\mux_cnt_122_11_g677/w_4, Gate, Tgate[1]);
	and \mux_cnt_122_11_g677/a_3(\mux_cnt_122_11_g677/w_3, n_326, Tgdel[1]);
	and \mux_cnt_122_11_g677/a_2(\mux_cnt_122_11_g677/w_2, n_746, cnt_nxt[1]);
	and \mux_cnt_122_11_g677/a_1(\mux_cnt_122_11_g677/w_1, Sync, Tsync[1]);
	and \mux_cnt_122_11_g677/a_0(\mux_cnt_122_11_g677/w_0, n_744, \mux_cnt_122_11_g677/data0);
	or \mux_cnt_122_11_g681/org(sub_wire8, \mux_cnt_122_11_g681/w_0, \mux_cnt_122_11_g681/w_1, \mux_cnt_122_11_g681/w_2, \mux_cnt_122_11_g681/w_3, \mux_cnt_122_11_g681/w_4);
	and \mux_cnt_122_11_g681/a_4(\mux_cnt_122_11_g681/w_4, Gate, Tgate[0]);
	and \mux_cnt_122_11_g681/a_3(\mux_cnt_122_11_g681/w_3, n_326, Tgdel[0]);
	and \mux_cnt_122_11_g681/a_2(\mux_cnt_122_11_g681/w_2, n_746, n_995);
	and \mux_cnt_122_11_g681/a_1(\mux_cnt_122_11_g681/w_1, Sync, Tsync[0]);
	and \mux_cnt_122_11_g681/a_0(\mux_cnt_122_11_g681/w_0, n_744, \mux_cnt_122_11_g681/data0);
	or \mux_cnt_122_11_g713/org(sub_wire9, \mux_cnt_122_11_g713/w_0, \mux_cnt_122_11_g713/w_1, \mux_cnt_122_11_g713/w_2, \mux_cnt_122_11_g713/w_3, \mux_cnt_122_11_g713/w_4);
	and \mux_cnt_122_11_g713/a_4(\mux_cnt_122_11_g713/w_4, Gate, Tgate[7]);
	and \mux_cnt_122_11_g713/a_3(\mux_cnt_122_11_g713/w_3, n_326, Tgdel[7]);
	and \mux_cnt_122_11_g713/a_2(\mux_cnt_122_11_g713/w_2, n_746, cnt_nxt[7]);
	and \mux_cnt_122_11_g713/a_1(\mux_cnt_122_11_g713/w_1, Sync, Tsync[7]);
	and \mux_cnt_122_11_g713/a_0(\mux_cnt_122_11_g713/w_0, n_744, \mux_cnt_122_11_g713/data0);
	or \mux_cnt_122_11_g653/org(sub_wire10, \mux_cnt_122_11_g653/w_0, \mux_cnt_122_11_g653/w_1, \mux_cnt_122_11_g653/w_2);
	and \mux_cnt_122_11_g653/a_2(\mux_cnt_122_11_g653/w_2, Gate, Tgate[15]);
	and \mux_cnt_122_11_g653/a_1(\mux_cnt_122_11_g653/w_1, n_746, cnt_nxt[15]);
	and \mux_cnt_122_11_g653/a_0(\mux_cnt_122_11_g653/w_0, n_741, \mux_cnt_122_11_g653/data0);
	or \mux_cnt_122_11_g685/org(sub_wire11, \mux_cnt_122_11_g685/w_0, \mux_cnt_122_11_g685/w_1, \mux_cnt_122_11_g685/w_2);
	and \mux_cnt_122_11_g685/a_2(\mux_cnt_122_11_g685/w_2, Gate, Tgate[14]);
	and \mux_cnt_122_11_g685/a_1(\mux_cnt_122_11_g685/w_1, n_746, cnt_nxt[14]);
	and \mux_cnt_122_11_g685/a_0(\mux_cnt_122_11_g685/w_0, n_741, \mux_cnt_122_11_g685/data0);
	or \mux_cnt_122_11_g689/org(sub_wire12, \mux_cnt_122_11_g689/w_0, \mux_cnt_122_11_g689/w_1, \mux_cnt_122_11_g689/w_2);
	and \mux_cnt_122_11_g689/a_2(\mux_cnt_122_11_g689/w_2, Gate, Tgate[13]);
	and \mux_cnt_122_11_g689/a_1(\mux_cnt_122_11_g689/w_1, n_746, cnt_nxt[13]);
	and \mux_cnt_122_11_g689/a_0(\mux_cnt_122_11_g689/w_0, n_741, \mux_cnt_122_11_g689/data0);
	or \mux_cnt_122_11_g693/org(sub_wire13, \mux_cnt_122_11_g693/w_0, \mux_cnt_122_11_g693/w_1, \mux_cnt_122_11_g693/w_2);
	and \mux_cnt_122_11_g693/a_2(\mux_cnt_122_11_g693/w_2, Gate, Tgate[12]);
	and \mux_cnt_122_11_g693/a_1(\mux_cnt_122_11_g693/w_1, n_746, cnt_nxt[12]);
	and \mux_cnt_122_11_g693/a_0(\mux_cnt_122_11_g693/w_0, n_741, \mux_cnt_122_11_g693/data0);
	or \mux_cnt_122_11_g697/org(sub_wire14, \mux_cnt_122_11_g697/w_0, \mux_cnt_122_11_g697/w_1, \mux_cnt_122_11_g697/w_2);
	and \mux_cnt_122_11_g697/a_2(\mux_cnt_122_11_g697/w_2, Gate, Tgate[11]);
	and \mux_cnt_122_11_g697/a_1(\mux_cnt_122_11_g697/w_1, n_746, cnt_nxt[11]);
	and \mux_cnt_122_11_g697/a_0(\mux_cnt_122_11_g697/w_0, n_741, \mux_cnt_122_11_g697/data0);
	or \mux_cnt_122_11_g701/org(sub_wire15, \mux_cnt_122_11_g701/w_0, \mux_cnt_122_11_g701/w_1, \mux_cnt_122_11_g701/w_2);
	and \mux_cnt_122_11_g701/a_2(\mux_cnt_122_11_g701/w_2, Gate, Tgate[10]);
	and \mux_cnt_122_11_g701/a_1(\mux_cnt_122_11_g701/w_1, n_746, cnt_nxt[10]);
	and \mux_cnt_122_11_g701/a_0(\mux_cnt_122_11_g701/w_0, n_741, \mux_cnt_122_11_g701/data0);
	or \mux_cnt_122_11_g705/org(sub_wire16, \mux_cnt_122_11_g705/w_0, \mux_cnt_122_11_g705/w_1, \mux_cnt_122_11_g705/w_2);
	and \mux_cnt_122_11_g705/a_2(\mux_cnt_122_11_g705/w_2, Gate, Tgate[9]);
	and \mux_cnt_122_11_g705/a_1(\mux_cnt_122_11_g705/w_1, n_746, cnt_nxt[9]);
	and \mux_cnt_122_11_g705/a_0(\mux_cnt_122_11_g705/w_0, n_741, \mux_cnt_122_11_g705/data0);
	or \mux_cnt_122_11_g709/org(sub_wire17, \mux_cnt_122_11_g709/w_0, \mux_cnt_122_11_g709/w_1, \mux_cnt_122_11_g709/w_2);
	and \mux_cnt_122_11_g709/a_2(\mux_cnt_122_11_g709/w_2, Gate, Tgate[8]);
	and \mux_cnt_122_11_g709/a_1(\mux_cnt_122_11_g709/w_1, n_746, cnt_nxt[8]);
	and \mux_cnt_122_11_g709/a_0(\mux_cnt_122_11_g709/w_0, n_741, \mux_cnt_122_11_g709/data0);
	nor sub_108_39_g111(sub_108_39_n_159, sub_108_39_n_949, prev_cnt[14]);
	xnor sub_108_39_g167(cnt_nxt[1], prev_cnt[0], prev_cnt[1]);
	xnor sub_108_39_g169(cnt_nxt[2], sub_108_39_n_103, prev_cnt[2]);
	xnor sub_108_39_g172(cnt_nxt[3], n_1052, prev_cnt[3]);
	xnor sub_108_39_g174(cnt_nxt[4], sub_108_39_n_139, prev_cnt[4]);
	xnor sub_108_39_g177(cnt_nxt[5], n_1241, prev_cnt[5]);
	xnor sub_108_39_g179(cnt_nxt[6], n_1062, prev_cnt[6]);
	xnor sub_108_39_g182(cnt_nxt[7], n_1242, prev_cnt[7]);
	xnor sub_108_39_g184(cnt_nxt[8], sub_108_39_n_166, prev_cnt[8]);
	xnor sub_108_39_g187(cnt_nxt[9], n_1245, prev_cnt[9]);
	xnor sub_108_39_g189(cnt_nxt[10], n_1246, prev_cnt[10]);
	xnor sub_108_39_g192(cnt_nxt[11], n_1247, prev_cnt[11]);
	xnor sub_108_39_g195(cnt_nxt[12], n_1069, prev_cnt[12]);
	xnor sub_108_39_g198(cnt_nxt[13], n_1248, prev_cnt[13]);
	xnor sub_108_39_g200(cnt_nxt[14], n_1249, prev_cnt[14]);
	xnor sub_108_39_g203(cnt_nxt[15], n_1250, prev_cnt[15]);
	not g1040(n_1184, prev_cnt[4]);
	not g1041(n_1185, prev_cnt[8]);
	not g1044(n_1188, prev_cnt[13]);
	not g1045(n_1189, prev_cnt[12]);
	nand g1059(sub_108_39_n_949, n_1188, n_1189);
	not g1060(n_1203, sub_108_39_n_159);
	not g1072(n_1212, sub_108_39_n_109);
	not g1079(n_1216, sub_108_39_n_151);
	nor g1104(n_1231, n_1212, prev_cnt[6]);
	nor g1110(n_1235, n_1216, prev_cnt[12]);
	nor g1111(n_1236, sub_108_39_n_949, n_1216);
	nor g1112(n_1237, n_1203, n_1216);
	nand g1116(n_1241, n_1382, n_1184);
	nand g1117(n_1242, n_1231, n_1382);
	nand g1120(n_1245, n_1387, n_1185);
	nand g1121(n_1246, sub_108_39_n_119, n_1387);
	nand g1122(n_1247, n_1049, n_1387);
	nand g1123(n_1248, n_1235, n_1387);
	nand g1124(n_1249, n_1236, n_1387);
	nand g1125(n_1250, n_1237, n_1387);
	nor g719(n_941, ena, rst);
	not g1097(n_1226, n_941);
	not g1054(n_1198, prev_state[4]);
	not g1053(n_1197, prev_state[3]);
	not g1052(n_1196, prev_state[2]);
	not g1051(n_1195, prev_state[1]);
	nand g1098(n_1227, n_1198, n_1197, n_1196, n_1195);
	not g1039(n_1183, prev_state[0]);
	nor g1099(n_1160, n_1227, n_1183);
	not g1100(n_1228, n_1160);
	not g1043(n_1187, ena);
	nor g1101(n_1229, n_1228, n_1187, rst);
	not g1102(n_1230, n_1229);
	nor g751(n_977, prev_cnt_len[14], prev_cnt_len[15], prev_cnt_len[12], prev_cnt_len[13]);
	nor g755(n_976, prev_cnt_len[4], prev_cnt_len[5], prev_cnt_len[6], prev_cnt_len[7]);
	nor g760(n_975, prev_cnt_len[10], prev_cnt_len[11], prev_cnt_len[8], prev_cnt_len[9]);
	not g1050(n_1194, prev_cnt_len[3]);
	not g1049(n_1193, prev_cnt_len[2]);
	not g1048(n_1192, prev_cnt_len[1]);
	not g1047(n_1191, prev_cnt_len[0]);
	nand g1063(n_1206, n_1194, n_1193, n_1192, n_1191);
	not g1064(n_1207, n_1206);
	nand g1065(sub_111_47_n_67, n_977, n_976, n_975, n_1207);
	nand g1061(n_1204, prev_state[4], n_1197, n_1196, n_1195);
	nor g22(n_45, n_1204, prev_state[0]);
	not g1062(n_1205, n_45);
	nor g1067(n_1161, n_1205, n_1187, rst);
	not g1068(n_1209, n_1161);
	nor g1069(sub_wire18, sub_111_47_n_67, n_1209);
	not g646(n_732, Done);
	nand g1103(sub_wire2, n_1230, n_732);
	not g843(n_1043, Sync);
	nand g1095(n_1224, n_1198, n_1197, n_1196, prev_state[1]);
	nor g16(n_43, n_1224, prev_state[0]);
	not g1096(n_1225, n_43);
	nor g1106(n_1164, n_1225, n_1187, rst);
	not g1107(n_1232, n_1164);
	nor g759(n_1078, prev_cnt[12], prev_cnt[13], prev_cnt[14], prev_cnt[15]);
	nor sub_108_39_g70(sub_108_39_n_119, prev_cnt[8], prev_cnt[9]);
	not g1073(n_1213, sub_108_39_n_119);
	nor g1076(n_1049, n_1213, prev_cnt[10]);
	not g1077(n_1215, n_1049);
	nor g1078(sub_108_39_n_151, n_1215, prev_cnt[11]);
	nor sub_108_39_g62(sub_108_39_n_109, prev_cnt[4], prev_cnt[5]);
	not g1046(n_1190, prev_cnt[1]);
	not g775(n_995, prev_cnt[0]);
	nand g1080(sub_108_39_n_103, n_1190, n_995);
	not g1081(n_1217, sub_108_39_n_103);
	not g1056(n_1200, prev_cnt[2]);
	nand g1082(n_1052, n_1217, n_1200);
	not g1083(n_1218, n_1052);
	not g1057(n_1201, prev_cnt[3]);
	nand g1084(sub_108_39_n_139, n_1218, n_1201);
	not g1085(n_1382, sub_108_39_n_139);
	nand g1086(n_1062, sub_108_39_n_109, n_1382);
	not g1087(n_1220, n_1062);
	not g1058(n_1202, prev_cnt[7]);
	not g1055(n_1199, prev_cnt[6]);
	nand g1088(sub_108_39_n_166, n_1220, n_1202, n_1199);
	not g1089(n_1387, sub_108_39_n_166);
	nand g1090(n_1069, sub_108_39_n_151, n_1387);
	not g1091(n_1222, n_1069);
	nand g1092(sub_108_39_n_67, n_1078, n_1222);
	nor g1126(n_326, n_1232, sub_108_39_n_67);
	not g1127(n_1251, n_326);
	nand g1132(n_1256, n_1226, n_1043, n_1251);
	not g1133(n_1257, n_1256);
	not g1042(n_1186, rst);
	nand g1135(n_741, n_1257, n_1186);
	not g1066(n_1208, sub_111_47_n_67);
	nor g1113(n_1238, n_1208, n_1209);
	not g1114(n_1239, n_1238);
	nand g1070(n_1210, n_1198, n_1197, prev_state[2], n_1195);
	nor g18(n_44, n_1210, prev_state[0]);
	not g1071(n_1211, n_44);
	nand g1108(n_1233, n_1205, n_1225, n_1228);
	not g1109(n_1234, n_1233);
	nand g1115(n_1240, n_1211, n_1234);
	nor g1118(n_1243, n_1240, n_1187, rst);
	not g1119(n_1244, n_1243);
	not g1093(n_1223, sub_108_39_n_67);
	nor g1128(n_1252, n_1232, n_1223);
	not g1129(n_1253, n_1252);
	nor g1074(n_1162, n_1211, n_1187, rst);
	not g1075(n_1214, n_1162);
	nor g1130(n_1254, n_1214, n_1223);
	not g1131(n_1255, n_1254);
	nand g1134(n_746, n_1239, n_1244, n_1253, n_1255);
	nor g1094(sub_wire1, n_1214, sub_108_39_n_67);
	nand g1105(n_744, n_1226, n_1186);
	assign w_eco0 = rst;
	and _ECO_1(w_eco1, !Tsync[6], prev_cnt[1], !prev_cnt[6], prev_cnt[9]);
	and _ECO_2(w_eco2, !Tsync[6], prev_cnt[2], !prev_cnt[6], prev_cnt[9]);
	and _ECO_3(w_eco3, !Tsync[6], prev_cnt[4], !prev_cnt[6], prev_cnt[9]);
	and _ECO_4(w_eco4, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[1], !prev_cnt[6]);
	and _ECO_5(w_eco5, !Tsync[6], prev_cnt[6], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6(w_eco6, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7(w_eco7, !Tsync[6], prev_cnt[0], !prev_cnt[6], prev_cnt[9]);
	and _ECO_8(w_eco8, !Tsync[6], prev_cnt[1], !prev_cnt[6], prev_cnt[15]);
	and _ECO_9(w_eco9, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[2], !prev_cnt[6]);
	and _ECO_10(w_eco10, !Tsync[6], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_11(w_eco11, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_12(w_eco12, !Tsync[6], prev_cnt[5], !prev_cnt[6], prev_cnt[9]);
	and _ECO_13(w_eco13, !Tsync[6], prev_cnt[1], !prev_cnt[6], prev_cnt[11]);
	and _ECO_14(w_eco14, !Tsync[6], prev_cnt[2], !prev_cnt[6], prev_cnt[15]);
	and _ECO_15(w_eco15, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[4], !prev_cnt[6]);
	and _ECO_16(w_eco16, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_17(w_eco17, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_18(w_eco18, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_19(w_eco19, !Tsync[6], prev_cnt[3], !prev_cnt[6], prev_cnt[9]);
	and _ECO_20(w_eco20, !Tsync[6], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6]);
	and _ECO_21(w_eco21, !Tsync[6], prev_cnt[1], !prev_cnt[6], prev_cnt[10]);
	and _ECO_22(w_eco22, !Tsync[6], prev_cnt[2], !prev_cnt[6], prev_cnt[11]);
	and _ECO_23(w_eco23, !Tsync[6], prev_cnt[4], !prev_cnt[6], prev_cnt[15]);
	and _ECO_24(w_eco24, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[0], !prev_cnt[6]);
	and _ECO_25(w_eco25, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_26(w_eco26, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_27(w_eco27, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_28(w_eco28, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_29(w_eco29, !Tsync[6], prev_cnt[1], !prev_cnt[6], prev_cnt[8]);
	and _ECO_30(w_eco30, !Tsync[6], prev_cnt[2], !prev_cnt[6], prev_cnt[10]);
	and _ECO_31(w_eco31, !Tsync[6], prev_cnt[4], !prev_cnt[6], prev_cnt[11]);
	and _ECO_32(w_eco32, !Tsync[6], prev_cnt[0], !prev_cnt[6], prev_cnt[15]);
	and _ECO_33(w_eco33, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[5], !prev_cnt[6]);
	and _ECO_34(w_eco34, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_35(w_eco35, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_36(w_eco36, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_37(w_eco37, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_38(w_eco38, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_39(w_eco39, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_40(w_eco40, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_41(w_eco41, !Tsync[6], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12]);
	and _ECO_42(w_eco42, !Tsync[6], prev_cnt[2], !prev_cnt[6], prev_cnt[8]);
	and _ECO_43(w_eco43, !Tsync[6], prev_cnt[4], !prev_cnt[6], prev_cnt[10]);
	and _ECO_44(w_eco44, !Tsync[6], prev_cnt[0], !prev_cnt[6], prev_cnt[11]);
	and _ECO_45(w_eco45, !Tsync[6], prev_cnt[5], !prev_cnt[6], prev_cnt[15]);
	and _ECO_46(w_eco46, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[3], !prev_cnt[6]);
	and _ECO_47(w_eco47, !Tsync[6], prev_cnt[9], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_48(w_eco48, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_49(w_eco49, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_50(w_eco50, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_51(w_eco51, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_52(w_eco52, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_53(w_eco53, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_54(w_eco54, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_55(w_eco55, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_56(w_eco56, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_57(w_eco57, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_58(w_eco58, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_59(w_eco59, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_60(w_eco60, !Tsync[6], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13]);
	and _ECO_61(w_eco61, !Tsync[6], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12]);
	and _ECO_62(w_eco62, !Tsync[6], prev_cnt[4], !prev_cnt[6], prev_cnt[8]);
	and _ECO_63(w_eco63, !Tsync[6], prev_cnt[0], !prev_cnt[6], prev_cnt[10]);
	and _ECO_64(w_eco64, !Tsync[6], prev_cnt[5], !prev_cnt[6], prev_cnt[11]);
	and _ECO_65(w_eco65, !Tsync[6], prev_cnt[3], !prev_cnt[6], prev_cnt[15]);
	and _ECO_66(w_eco66, !Tsync[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_67(w_eco67, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_68(w_eco68, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_69(w_eco69, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_70(w_eco70, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_71(w_eco71, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_72(w_eco72, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_73(w_eco73, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_74(w_eco74, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_75(w_eco75, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_76(w_eco76, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_77(w_eco77, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_78(w_eco78, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_79(w_eco79, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_80(w_eco80, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_81(w_eco81, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_82(w_eco82, !Tsync[6], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13]);
	and _ECO_83(w_eco83, !Tsync[6], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12]);
	and _ECO_84(w_eco84, !Tsync[6], prev_cnt[0], !prev_cnt[6], prev_cnt[8]);
	and _ECO_85(w_eco85, !Tsync[6], prev_cnt[5], !prev_cnt[6], prev_cnt[10]);
	and _ECO_86(w_eco86, !Tsync[6], prev_cnt[3], !prev_cnt[6], prev_cnt[11]);
	and _ECO_87(w_eco87, !Tgdel[6], !Tsync[6], prev_cnt[1], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_88(w_eco88, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_89(w_eco89, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_90(w_eco90, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_91(w_eco91, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_92(w_eco92, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_93(w_eco93, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_94(w_eco94, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_95(w_eco95, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_96(w_eco96, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_97(w_eco97, !Tgate[6], !Tsync[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_98(w_eco98, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_99(w_eco99, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_100(w_eco100, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_101(w_eco101, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_102(w_eco102, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_103(w_eco103, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_104(w_eco104, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_105(w_eco105, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_106(w_eco106, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_107(w_eco107, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_108(w_eco108, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_109(w_eco109, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_110(w_eco110, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_111(w_eco111, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_112(w_eco112, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_113(w_eco113, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_114(w_eco114, !Tsync[6], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13]);
	and _ECO_115(w_eco115, !Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12]);
	and _ECO_116(w_eco116, !Tsync[6], prev_cnt[5], !prev_cnt[6], prev_cnt[8]);
	and _ECO_117(w_eco117, !Tsync[6], prev_cnt[3], !prev_cnt[6], prev_cnt[10]);
	and _ECO_118(w_eco118, !Tsync[6], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_119(w_eco119, !Tgdel[6], !Tsync[6], prev_cnt[2], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_120(w_eco120, !Tgdel[6], !Tsync[6], prev_cnt[1], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_121(w_eco121, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_122(w_eco122, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_123(w_eco123, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_124(w_eco124, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_125(w_eco125, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_126(w_eco126, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_127(w_eco127, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_128(w_eco128, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_129(w_eco129, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_130(w_eco130, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_131(w_eco131, !Tgate[6], !Tsync[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_132(w_eco132, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_133(w_eco133, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_134(w_eco134, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_135(w_eco135, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_136(w_eco136, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_137(w_eco137, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_138(w_eco138, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_139(w_eco139, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_140(w_eco140, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_141(w_eco141, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_142(w_eco142, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_143(w_eco143, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_144(w_eco144, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_145(w_eco145, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_146(w_eco146, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_147(w_eco147, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_148(w_eco148, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_149(w_eco149, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_150(w_eco150, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_151(w_eco151, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_152(w_eco152, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_153(w_eco153, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_154(w_eco154, !Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13]);
	and _ECO_155(w_eco155, !Tsync[6], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12]);
	and _ECO_156(w_eco156, !Tsync[6], prev_cnt[3], !prev_cnt[6], prev_cnt[8]);
	and _ECO_157(w_eco157, !Tgdel[6], !Tsync[6], prev_cnt[4], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_158(w_eco158, !Tsync[6], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_159(w_eco159, !Tgdel[6], !Tsync[6], prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_160(w_eco160, !Tgate[6], !Tsync[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_161(w_eco161, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_162(w_eco162, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_163(w_eco163, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_164(w_eco164, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_165(w_eco165, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_166(w_eco166, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_167(w_eco167, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_168(w_eco168, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_169(w_eco169, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_170(w_eco170, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_171(w_eco171, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_172(w_eco172, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_173(w_eco173, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_174(w_eco174, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_175(w_eco175, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_176(w_eco176, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_177(w_eco177, !Tgate[6], !Tsync[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_178(w_eco178, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_179(w_eco179, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_180(w_eco180, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_181(w_eco181, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_182(w_eco182, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_183(w_eco183, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_184(w_eco184, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_185(w_eco185, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_186(w_eco186, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_187(w_eco187, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_188(w_eco188, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_189(w_eco189, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_190(w_eco190, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_191(w_eco191, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_192(w_eco192, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_193(w_eco193, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_194(w_eco194, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_195(w_eco195, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_196(w_eco196, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_197(w_eco197, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_198(w_eco198, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_199(w_eco199, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_200(w_eco200, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_201(w_eco201, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_202(w_eco202, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_203(w_eco203, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_204(w_eco204, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_205(w_eco205, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_206(w_eco206, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_207(w_eco207, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_208(w_eco208, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_209(w_eco209, !Tsync[6], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13]);
	and _ECO_210(w_eco210, !Tsync[6], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12]);
	and _ECO_211(w_eco211, !Tsync[6], prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_212(w_eco212, !Tgdel[6], !Tsync[6], prev_cnt[0], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_213(w_eco213, !Tgdel[6], !Tsync[6], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_214(w_eco214, !Tgate[6], !Tsync[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_215(w_eco215, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_216(w_eco216, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_217(w_eco217, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_218(w_eco218, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_219(w_eco219, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_220(w_eco220, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_221(w_eco221, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_222(w_eco222, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_223(w_eco223, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_224(w_eco224, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_225(w_eco225, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_226(w_eco226, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_227(w_eco227, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_228(w_eco228, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_229(w_eco229, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_230(w_eco230, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_231(w_eco231, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_232(w_eco232, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_233(w_eco233, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_234(w_eco234, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_235(w_eco235, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_236(w_eco236, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_237(w_eco237, !Tgate[6], !Tsync[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_238(w_eco238, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_239(w_eco239, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_240(w_eco240, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_241(w_eco241, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_242(w_eco242, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_243(w_eco243, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_244(w_eco244, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_245(w_eco245, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_246(w_eco246, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_247(w_eco247, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_248(w_eco248, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_249(w_eco249, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_250(w_eco250, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_251(w_eco251, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_252(w_eco252, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_253(w_eco253, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_254(w_eco254, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_255(w_eco255, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_256(w_eco256, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_257(w_eco257, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_258(w_eco258, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_259(w_eco259, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_260(w_eco260, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_261(w_eco261, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_262(w_eco262, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_263(w_eco263, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_264(w_eco264, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_265(w_eco265, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_266(w_eco266, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_267(w_eco267, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_268(w_eco268, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_269(w_eco269, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_270(w_eco270, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_271(w_eco271, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_272(w_eco272, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_273(w_eco273, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_274(w_eco274, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_275(w_eco275, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_276(w_eco276, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_277(w_eco277, !Tsync[6], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13]);
	and _ECO_278(w_eco278, !Tsync[6], prev_cnt[11], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_279(w_eco279, !Tsync[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_280(w_eco280, !Tgdel[6], !Tsync[6], prev_cnt[5], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_281(w_eco281, !Tsync[6], prev_cnt[10], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_282(w_eco282, !Tgdel[6], !Tsync[6], prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_283(w_eco283, !Tsync[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_284(w_eco284, !Tgate[6], !Tsync[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_285(w_eco285, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_286(w_eco286, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_287(w_eco287, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_288(w_eco288, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_289(w_eco289, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_290(w_eco290, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_291(w_eco291, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_292(w_eco292, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_293(w_eco293, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_294(w_eco294, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_295(w_eco295, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_296(w_eco296, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_297(w_eco297, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_298(w_eco298, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_299(w_eco299, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_300(w_eco300, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_301(w_eco301, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_302(w_eco302, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_303(w_eco303, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_304(w_eco304, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_305(w_eco305, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_306(w_eco306, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_307(w_eco307, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_308(w_eco308, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_309(w_eco309, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_310(w_eco310, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_311(w_eco311, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_312(w_eco312, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_313(w_eco313, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_314(w_eco314, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_315(w_eco315, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_316(w_eco316, !Tgate[6], !Tsync[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_317(w_eco317, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_318(w_eco318, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_319(w_eco319, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_320(w_eco320, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_321(w_eco321, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_322(w_eco322, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_323(w_eco323, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_324(w_eco324, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_325(w_eco325, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_326(w_eco326, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_327(w_eco327, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_328(w_eco328, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_329(w_eco329, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_330(w_eco330, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_331(w_eco331, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_332(w_eco332, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_333(w_eco333, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_334(w_eco334, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_335(w_eco335, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_336(w_eco336, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_337(w_eco337, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_338(w_eco338, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_339(w_eco339, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_340(w_eco340, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_341(w_eco341, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_342(w_eco342, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_343(w_eco343, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_344(w_eco344, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_345(w_eco345, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_346(w_eco346, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_347(w_eco347, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_348(w_eco348, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_349(w_eco349, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_350(w_eco350, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_351(w_eco351, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_352(w_eco352, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_353(w_eco353, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_354(w_eco354, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_355(w_eco355, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_356(w_eco356, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_357(w_eco357, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_358(w_eco358, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_359(w_eco359, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_360(w_eco360, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_361(w_eco361, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_362(w_eco362, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_363(w_eco363, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_364(w_eco364, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_365(w_eco365, !Tsync[6], prev_cnt[8], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_366(w_eco366, !Tgdel[6], !Tsync[6], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_367(w_eco367, !Tsync[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_368(w_eco368, !Tgate[6], !Tsync[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_369(w_eco369, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_370(w_eco370, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_371(w_eco371, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_372(w_eco372, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_373(w_eco373, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_374(w_eco374, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_375(w_eco375, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_376(w_eco376, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_377(w_eco377, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_378(w_eco378, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_379(w_eco379, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_380(w_eco380, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_381(w_eco381, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_382(w_eco382, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_383(w_eco383, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_384(w_eco384, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_385(w_eco385, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_386(w_eco386, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_387(w_eco387, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_388(w_eco388, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_389(w_eco389, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_390(w_eco390, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_391(w_eco391, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_392(w_eco392, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_393(w_eco393, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_394(w_eco394, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_395(w_eco395, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_396(w_eco396, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_397(w_eco397, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_398(w_eco398, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_399(w_eco399, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_400(w_eco400, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_401(w_eco401, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_402(w_eco402, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_403(w_eco403, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_404(w_eco404, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_405(w_eco405, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_406(w_eco406, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_407(w_eco407, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_408(w_eco408, !Tgate[6], !Tsync[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_409(w_eco409, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_410(w_eco410, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_411(w_eco411, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_412(w_eco412, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_413(w_eco413, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_414(w_eco414, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_415(w_eco415, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_416(w_eco416, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_417(w_eco417, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_418(w_eco418, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_419(w_eco419, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_420(w_eco420, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_421(w_eco421, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_422(w_eco422, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_423(w_eco423, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_424(w_eco424, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_425(w_eco425, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_426(w_eco426, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_427(w_eco427, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_428(w_eco428, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_429(w_eco429, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_430(w_eco430, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_431(w_eco431, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_432(w_eco432, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_433(w_eco433, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_434(w_eco434, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_435(w_eco435, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_436(w_eco436, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_437(w_eco437, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_438(w_eco438, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_439(w_eco439, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_440(w_eco440, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_441(w_eco441, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_442(w_eco442, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_443(w_eco443, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_444(w_eco444, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_445(w_eco445, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_446(w_eco446, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_447(w_eco447, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_448(w_eco448, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_449(w_eco449, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_450(w_eco450, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_451(w_eco451, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_452(w_eco452, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_453(w_eco453, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_454(w_eco454, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_455(w_eco455, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_456(w_eco456, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_457(w_eco457, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_458(w_eco458, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_459(w_eco459, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_460(w_eco460, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_461(w_eco461, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_462(w_eco462, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_463(w_eco463, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_464(w_eco464, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_465(w_eco465, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_466(w_eco466, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_467(w_eco467, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_468(w_eco468, !Tgdel[6], !Tsync[6], prev_cnt[3], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_469(w_eco469, !Tsync[6], !prev_cnt[14], prev_cnt[12], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_470(w_eco470, !Tsync[6], !prev_cnt[14], prev_cnt[13], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_471(w_eco471, !Tsync[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_472(w_eco472, !Tgate[6], !Tsync[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_473(w_eco473, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_474(w_eco474, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_475(w_eco475, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_476(w_eco476, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_477(w_eco477, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_478(w_eco478, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_479(w_eco479, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_480(w_eco480, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_481(w_eco481, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_482(w_eco482, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_483(w_eco483, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_484(w_eco484, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_485(w_eco485, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_486(w_eco486, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_487(w_eco487, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_488(w_eco488, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_489(w_eco489, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_490(w_eco490, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_491(w_eco491, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_492(w_eco492, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_493(w_eco493, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_494(w_eco494, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_495(w_eco495, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_496(w_eco496, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_497(w_eco497, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_498(w_eco498, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_499(w_eco499, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_500(w_eco500, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_501(w_eco501, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_502(w_eco502, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_503(w_eco503, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_504(w_eco504, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_505(w_eco505, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_506(w_eco506, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_507(w_eco507, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_508(w_eco508, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_509(w_eco509, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_510(w_eco510, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_511(w_eco511, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_512(w_eco512, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_513(w_eco513, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_514(w_eco514, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_515(w_eco515, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_516(w_eco516, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_517(w_eco517, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_518(w_eco518, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_519(w_eco519, prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_520(w_eco520, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_521(w_eco521, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_522(w_eco522, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_523(w_eco523, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_524(w_eco524, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_525(w_eco525, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_526(w_eco526, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_527(w_eco527, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_528(w_eco528, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_529(w_eco529, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_530(w_eco530, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_531(w_eco531, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_532(w_eco532, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_533(w_eco533, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_534(w_eco534, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_535(w_eco535, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_536(w_eco536, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_537(w_eco537, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_538(w_eco538, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_539(w_eco539, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_540(w_eco540, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_541(w_eco541, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_542(w_eco542, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_543(w_eco543, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_544(w_eco544, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_545(w_eco545, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_546(w_eco546, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_547(w_eco547, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_548(w_eco548, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_549(w_eco549, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_550(w_eco550, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_551(w_eco551, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_552(w_eco552, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_553(w_eco553, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_554(w_eco554, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_555(w_eco555, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_556(w_eco556, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_557(w_eco557, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_558(w_eco558, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_559(w_eco559, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_560(w_eco560, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_561(w_eco561, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_562(w_eco562, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_563(w_eco563, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_564(w_eco564, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_565(w_eco565, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_566(w_eco566, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_567(w_eco567, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_568(w_eco568, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_569(w_eco569, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_570(w_eco570, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_571(w_eco571, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_572(w_eco572, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_573(w_eco573, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_574(w_eco574, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_575(w_eco575, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_576(w_eco576, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_577(w_eco577, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_578(w_eco578, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_579(w_eco579, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_580(w_eco580, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_581(w_eco581, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_582(w_eco582, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_583(w_eco583, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_584(w_eco584, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_585(w_eco585, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_586(w_eco586, !Tgate[6], !Tgdel[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_587(w_eco587, !Tgdel[6], !Tsync[6], prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_588(w_eco588, !Tsync[6], !prev_cnt[14], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_589(w_eco589, !Tsync[6], !prev_cnt[14], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_590(w_eco590, !Tgate[6], !Tsync[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_591(w_eco591, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_592(w_eco592, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_593(w_eco593, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_594(w_eco594, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_595(w_eco595, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_596(w_eco596, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_597(w_eco597, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_598(w_eco598, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_599(w_eco599, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_600(w_eco600, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_601(w_eco601, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_602(w_eco602, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_603(w_eco603, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_604(w_eco604, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_605(w_eco605, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_606(w_eco606, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_607(w_eco607, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_608(w_eco608, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_609(w_eco609, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_610(w_eco610, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_611(w_eco611, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_612(w_eco612, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_613(w_eco613, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_614(w_eco614, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_615(w_eco615, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_616(w_eco616, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_617(w_eco617, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_618(w_eco618, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_619(w_eco619, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_620(w_eco620, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_621(w_eco621, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_622(w_eco622, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_623(w_eco623, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_624(w_eco624, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_625(w_eco625, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_626(w_eco626, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_627(w_eco627, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_628(w_eco628, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_629(w_eco629, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_630(w_eco630, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_631(w_eco631, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_632(w_eco632, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_633(w_eco633, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_634(w_eco634, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_635(w_eco635, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_636(w_eco636, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_637(w_eco637, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_638(w_eco638, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_639(w_eco639, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_640(w_eco640, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_641(w_eco641, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_642(w_eco642, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_643(w_eco643, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_644(w_eco644, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_645(w_eco645, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_646(w_eco646, prev_cnt[2], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_647(w_eco647, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_648(w_eco648, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_649(w_eco649, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_650(w_eco650, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_651(w_eco651, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_652(w_eco652, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_653(w_eco653, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_654(w_eco654, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_655(w_eco655, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_656(w_eco656, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_657(w_eco657, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_658(w_eco658, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_659(w_eco659, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_660(w_eco660, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_661(w_eco661, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_662(w_eco662, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_663(w_eco663, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_664(w_eco664, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_665(w_eco665, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_666(w_eco666, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_667(w_eco667, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_668(w_eco668, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_669(w_eco669, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_670(w_eco670, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_671(w_eco671, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_672(w_eco672, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_673(w_eco673, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_674(w_eco674, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_675(w_eco675, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_676(w_eco676, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_677(w_eco677, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_678(w_eco678, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_679(w_eco679, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_680(w_eco680, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_681(w_eco681, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_682(w_eco682, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_683(w_eco683, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_684(w_eco684, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_685(w_eco685, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_686(w_eco686, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_687(w_eco687, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_688(w_eco688, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_689(w_eco689, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_690(w_eco690, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_691(w_eco691, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_692(w_eco692, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_693(w_eco693, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_694(w_eco694, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_695(w_eco695, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_696(w_eco696, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_697(w_eco697, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_698(w_eco698, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_699(w_eco699, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_700(w_eco700, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_701(w_eco701, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_702(w_eco702, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_703(w_eco703, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_704(w_eco704, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_705(w_eco705, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_706(w_eco706, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_707(w_eco707, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_708(w_eco708, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_709(w_eco709, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_710(w_eco710, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_711(w_eco711, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_712(w_eco712, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_713(w_eco713, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_714(w_eco714, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_715(w_eco715, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_716(w_eco716, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_717(w_eco717, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_718(w_eco718, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_719(w_eco719, !Tgate[6], !Tgdel[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_720(w_eco720, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_721(w_eco721, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_722(w_eco722, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_723(w_eco723, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_724(w_eco724, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_725(w_eco725, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_726(w_eco726, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_727(w_eco727, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_728(w_eco728, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_729(w_eco729, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_730(w_eco730, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_731(w_eco731, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_732(w_eco732, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_733(w_eco733, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_734(w_eco734, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_735(w_eco735, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_736(w_eco736, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_737(w_eco737, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_738(w_eco738, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_739(w_eco739, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_740(w_eco740, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_741(w_eco741, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_742(w_eco742, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_743(w_eco743, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_744(w_eco744, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_745(w_eco745, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_746(w_eco746, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_747(w_eco747, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_748(w_eco748, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_749(w_eco749, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_750(w_eco750, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_751(w_eco751, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_752(w_eco752, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_753(w_eco753, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_754(w_eco754, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_755(w_eco755, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_756(w_eco756, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_757(w_eco757, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_758(w_eco758, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_759(w_eco759, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_760(w_eco760, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_761(w_eco761, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_762(w_eco762, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_763(w_eco763, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_764(w_eco764, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_765(w_eco765, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_766(w_eco766, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_767(w_eco767, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_768(w_eco768, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_769(w_eco769, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_770(w_eco770, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_771(w_eco771, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_772(w_eco772, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_773(w_eco773, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_774(w_eco774, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_775(w_eco775, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_776(w_eco776, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_777(w_eco777, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_778(w_eco778, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_779(w_eco779, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_780(w_eco780, prev_cnt[4], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_781(w_eco781, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_782(w_eco782, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_783(w_eco783, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_784(w_eco784, !Tgate[6], !Tgdel[6], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_785(w_eco785, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_786(w_eco786, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_787(w_eco787, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_788(w_eco788, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_789(w_eco789, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_790(w_eco790, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_791(w_eco791, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_792(w_eco792, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_793(w_eco793, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_794(w_eco794, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_795(w_eco795, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_796(w_eco796, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_797(w_eco797, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_798(w_eco798, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_799(w_eco799, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_800(w_eco800, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_801(w_eco801, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_802(w_eco802, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_803(w_eco803, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_804(w_eco804, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_805(w_eco805, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_806(w_eco806, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_807(w_eco807, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_808(w_eco808, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_809(w_eco809, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_810(w_eco810, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_811(w_eco811, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_812(w_eco812, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_813(w_eco813, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_814(w_eco814, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_815(w_eco815, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_816(w_eco816, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_817(w_eco817, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_818(w_eco818, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_819(w_eco819, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_820(w_eco820, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_821(w_eco821, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_822(w_eco822, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_823(w_eco823, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_824(w_eco824, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_825(w_eco825, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_826(w_eco826, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_827(w_eco827, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_828(w_eco828, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_829(w_eco829, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_830(w_eco830, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_831(w_eco831, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_832(w_eco832, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_833(w_eco833, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_834(w_eco834, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_835(w_eco835, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_836(w_eco836, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_837(w_eco837, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_838(w_eco838, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_839(w_eco839, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_840(w_eco840, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_841(w_eco841, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_842(w_eco842, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_843(w_eco843, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_844(w_eco844, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_845(w_eco845, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_846(w_eco846, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_847(w_eco847, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_848(w_eco848, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_849(w_eco849, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_850(w_eco850, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_851(w_eco851, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_852(w_eco852, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_853(w_eco853, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_854(w_eco854, !Tgate[6], !Tgdel[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_855(w_eco855, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_856(w_eco856, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_857(w_eco857, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_858(w_eco858, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_859(w_eco859, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_860(w_eco860, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_861(w_eco861, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_862(w_eco862, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_863(w_eco863, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_864(w_eco864, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_865(w_eco865, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_866(w_eco866, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_867(w_eco867, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_868(w_eco868, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_869(w_eco869, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_870(w_eco870, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_871(w_eco871, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_872(w_eco872, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_873(w_eco873, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_874(w_eco874, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_875(w_eco875, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_876(w_eco876, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_877(w_eco877, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_878(w_eco878, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_879(w_eco879, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_880(w_eco880, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_881(w_eco881, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_882(w_eco882, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_883(w_eco883, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_884(w_eco884, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_885(w_eco885, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_886(w_eco886, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_887(w_eco887, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_888(w_eco888, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_889(w_eco889, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_890(w_eco890, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_891(w_eco891, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_892(w_eco892, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_893(w_eco893, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_894(w_eco894, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_895(w_eco895, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_896(w_eco896, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_897(w_eco897, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_898(w_eco898, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_899(w_eco899, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_900(w_eco900, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_901(w_eco901, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_902(w_eco902, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_903(w_eco903, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_904(w_eco904, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_905(w_eco905, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_906(w_eco906, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_907(w_eco907, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_908(w_eco908, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_909(w_eco909, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_910(w_eco910, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_911(w_eco911, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_912(w_eco912, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_913(w_eco913, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_914(w_eco914, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_915(w_eco915, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_916(w_eco916, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_917(w_eco917, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_918(w_eco918, prev_cnt[0], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_919(w_eco919, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_920(w_eco920, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_921(w_eco921, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_922(w_eco922, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_923(w_eco923, prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_924(w_eco924, !Tgate[6], !Tgdel[6], prev_cnt[2], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_925(w_eco925, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_926(w_eco926, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_927(w_eco927, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_928(w_eco928, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_929(w_eco929, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_930(w_eco930, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_931(w_eco931, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_932(w_eco932, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_933(w_eco933, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_934(w_eco934, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_935(w_eco935, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_936(w_eco936, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_937(w_eco937, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_938(w_eco938, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_939(w_eco939, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_940(w_eco940, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_941(w_eco941, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_942(w_eco942, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_943(w_eco943, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_944(w_eco944, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_945(w_eco945, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_946(w_eco946, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_947(w_eco947, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_948(w_eco948, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_949(w_eco949, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_950(w_eco950, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_951(w_eco951, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_952(w_eco952, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_953(w_eco953, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_954(w_eco954, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_955(w_eco955, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_956(w_eco956, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_957(w_eco957, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_958(w_eco958, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_959(w_eco959, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_960(w_eco960, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_961(w_eco961, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_962(w_eco962, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_963(w_eco963, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_964(w_eco964, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_965(w_eco965, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_966(w_eco966, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_967(w_eco967, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_968(w_eco968, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_969(w_eco969, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_970(w_eco970, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_971(w_eco971, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_972(w_eco972, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_973(w_eco973, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_974(w_eco974, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_975(w_eco975, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_976(w_eco976, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_977(w_eco977, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_978(w_eco978, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_979(w_eco979, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_980(w_eco980, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_981(w_eco981, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_982(w_eco982, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_983(w_eco983, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_984(w_eco984, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_985(w_eco985, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_986(w_eco986, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_987(w_eco987, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_988(w_eco988, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_989(w_eco989, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_990(w_eco990, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_991(w_eco991, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_992(w_eco992, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_993(w_eco993, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_994(w_eco994, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_995(w_eco995, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_996(w_eco996, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_997(w_eco997, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_998(w_eco998, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_999(w_eco999, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1000(w_eco1000, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1001(w_eco1001, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1002(w_eco1002, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1003(w_eco1003, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1004(w_eco1004, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1005(w_eco1005, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1006(w_eco1006, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1007(w_eco1007, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1008(w_eco1008, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1009(w_eco1009, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1010(w_eco1010, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1011(w_eco1011, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1012(w_eco1012, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1013(w_eco1013, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1014(w_eco1014, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1015(w_eco1015, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1016(w_eco1016, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1017(w_eco1017, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1018(w_eco1018, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1019(w_eco1019, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1020(w_eco1020, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1021(w_eco1021, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1022(w_eco1022, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1023(w_eco1023, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1024(w_eco1024, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1025(w_eco1025, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1026(w_eco1026, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1027(w_eco1027, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1028(w_eco1028, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1029(w_eco1029, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1030(w_eco1030, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1031(w_eco1031, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1032(w_eco1032, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1033(w_eco1033, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1034(w_eco1034, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1035(w_eco1035, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1036(w_eco1036, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1037(w_eco1037, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1038(w_eco1038, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1039(w_eco1039, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1040(w_eco1040, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1041(w_eco1041, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1042(w_eco1042, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1043(w_eco1043, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1044(w_eco1044, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1045(w_eco1045, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1046(w_eco1046, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1047(w_eco1047, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1048(w_eco1048, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1049(w_eco1049, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1050(w_eco1050, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1051(w_eco1051, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1052(w_eco1052, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1053(w_eco1053, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1054(w_eco1054, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1055(w_eco1055, prev_cnt[5], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1056(w_eco1056, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1057(w_eco1057, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1058(w_eco1058, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1059(w_eco1059, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1060(w_eco1060, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1061(w_eco1061, prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1062(w_eco1062, prev_cnt[2], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1063(w_eco1063, !Tgate[6], !Tgdel[6], prev_cnt[4], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1064(w_eco1064, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1065(w_eco1065, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1066(w_eco1066, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1067(w_eco1067, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1068(w_eco1068, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1069(w_eco1069, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1070(w_eco1070, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1071(w_eco1071, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1072(w_eco1072, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1073(w_eco1073, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1074(w_eco1074, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1075(w_eco1075, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1076(w_eco1076, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1077(w_eco1077, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1078(w_eco1078, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1079(w_eco1079, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1080(w_eco1080, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1081(w_eco1081, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1082(w_eco1082, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1083(w_eco1083, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1084(w_eco1084, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1085(w_eco1085, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1086(w_eco1086, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1087(w_eco1087, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1088(w_eco1088, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1089(w_eco1089, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1090(w_eco1090, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1091(w_eco1091, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1092(w_eco1092, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1093(w_eco1093, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1094(w_eco1094, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1095(w_eco1095, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1096(w_eco1096, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1097(w_eco1097, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1098(w_eco1098, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1099(w_eco1099, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1100(w_eco1100, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1101(w_eco1101, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1102(w_eco1102, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1103(w_eco1103, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1104(w_eco1104, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1105(w_eco1105, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1106(w_eco1106, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1107(w_eco1107, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1108(w_eco1108, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1109(w_eco1109, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1110(w_eco1110, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1111(w_eco1111, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1112(w_eco1112, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1113(w_eco1113, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1114(w_eco1114, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1115(w_eco1115, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1116(w_eco1116, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1117(w_eco1117, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1118(w_eco1118, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1119(w_eco1119, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1120(w_eco1120, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1121(w_eco1121, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1122(w_eco1122, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1123(w_eco1123, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1124(w_eco1124, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1125(w_eco1125, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1126(w_eco1126, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1127(w_eco1127, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1128(w_eco1128, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1129(w_eco1129, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1130(w_eco1130, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1131(w_eco1131, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1132(w_eco1132, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1133(w_eco1133, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1134(w_eco1134, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1135(w_eco1135, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1136(w_eco1136, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1137(w_eco1137, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1138(w_eco1138, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1139(w_eco1139, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1140(w_eco1140, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1141(w_eco1141, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1142(w_eco1142, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1143(w_eco1143, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1144(w_eco1144, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1145(w_eco1145, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1146(w_eco1146, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1147(w_eco1147, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1148(w_eco1148, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1149(w_eco1149, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1150(w_eco1150, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1151(w_eco1151, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1152(w_eco1152, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1153(w_eco1153, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1154(w_eco1154, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1155(w_eco1155, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1156(w_eco1156, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1157(w_eco1157, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1158(w_eco1158, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1159(w_eco1159, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1160(w_eco1160, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1161(w_eco1161, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1162(w_eco1162, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1163(w_eco1163, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1164(w_eco1164, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1165(w_eco1165, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1166(w_eco1166, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1167(w_eco1167, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1168(w_eco1168, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1169(w_eco1169, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1170(w_eco1170, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1171(w_eco1171, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1172(w_eco1172, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1173(w_eco1173, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1174(w_eco1174, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1175(w_eco1175, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1176(w_eco1176, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1177(w_eco1177, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1178(w_eco1178, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1179(w_eco1179, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1180(w_eco1180, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1181(w_eco1181, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1182(w_eco1182, prev_cnt[3], !prev_cnt[6], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1183(w_eco1183, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1184(w_eco1184, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1185(w_eco1185, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1186(w_eco1186, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1187(w_eco1187, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1188(w_eco1188, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1189(w_eco1189, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1190(w_eco1190, prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1191(w_eco1191, prev_cnt[2], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1192(w_eco1192, prev_cnt[4], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1193(w_eco1193, !Tgate[6], !Tgdel[6], prev_cnt[0], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1194(w_eco1194, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1195(w_eco1195, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1196(w_eco1196, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1197(w_eco1197, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1198(w_eco1198, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1199(w_eco1199, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1200(w_eco1200, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1201(w_eco1201, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1202(w_eco1202, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1203(w_eco1203, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1204(w_eco1204, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1205(w_eco1205, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1206(w_eco1206, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1207(w_eco1207, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1208(w_eco1208, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1209(w_eco1209, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1210(w_eco1210, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1211(w_eco1211, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1212(w_eco1212, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1213(w_eco1213, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1214(w_eco1214, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1215(w_eco1215, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1216(w_eco1216, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1217(w_eco1217, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1218(w_eco1218, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1219(w_eco1219, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1220(w_eco1220, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1221(w_eco1221, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1222(w_eco1222, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1223(w_eco1223, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1224(w_eco1224, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1225(w_eco1225, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1226(w_eco1226, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1227(w_eco1227, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1228(w_eco1228, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1229(w_eco1229, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1230(w_eco1230, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1231(w_eco1231, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1232(w_eco1232, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1233(w_eco1233, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1234(w_eco1234, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1235(w_eco1235, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1236(w_eco1236, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1237(w_eco1237, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1238(w_eco1238, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1239(w_eco1239, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1240(w_eco1240, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1241(w_eco1241, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1242(w_eco1242, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1243(w_eco1243, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1244(w_eco1244, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1245(w_eco1245, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1246(w_eco1246, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1247(w_eco1247, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1248(w_eco1248, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1249(w_eco1249, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1250(w_eco1250, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1251(w_eco1251, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1252(w_eco1252, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1253(w_eco1253, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1254(w_eco1254, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1255(w_eco1255, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1256(w_eco1256, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1257(w_eco1257, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1258(w_eco1258, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1259(w_eco1259, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1260(w_eco1260, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1261(w_eco1261, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1262(w_eco1262, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1263(w_eco1263, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1264(w_eco1264, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1265(w_eco1265, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1266(w_eco1266, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1267(w_eco1267, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1268(w_eco1268, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1269(w_eco1269, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1270(w_eco1270, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1271(w_eco1271, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1272(w_eco1272, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1273(w_eco1273, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1274(w_eco1274, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1275(w_eco1275, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1276(w_eco1276, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1277(w_eco1277, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1278(w_eco1278, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1279(w_eco1279, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1280(w_eco1280, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1281(w_eco1281, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1282(w_eco1282, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1283(w_eco1283, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1284(w_eco1284, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1285(w_eco1285, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1286(w_eco1286, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1287(w_eco1287, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1288(w_eco1288, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1289(w_eco1289, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1290(w_eco1290, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1291(w_eco1291, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1292(w_eco1292, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1293(w_eco1293, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1294(w_eco1294, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1295(w_eco1295, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1296(w_eco1296, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1297(w_eco1297, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1298(w_eco1298, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1299(w_eco1299, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1300(w_eco1300, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1301(w_eco1301, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1302(w_eco1302, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1303(w_eco1303, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1304(w_eco1304, prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1305(w_eco1305, prev_cnt[2], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1306(w_eco1306, prev_cnt[4], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1307(w_eco1307, prev_cnt[0], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1308(w_eco1308, !Tgate[6], !Tgdel[6], prev_cnt[5], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1309(w_eco1309, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1310(w_eco1310, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1311(w_eco1311, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1312(w_eco1312, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1313(w_eco1313, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1314(w_eco1314, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1315(w_eco1315, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1316(w_eco1316, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1317(w_eco1317, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1318(w_eco1318, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1319(w_eco1319, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1320(w_eco1320, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1321(w_eco1321, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1322(w_eco1322, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1323(w_eco1323, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1324(w_eco1324, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1325(w_eco1325, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1326(w_eco1326, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1327(w_eco1327, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1328(w_eco1328, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1329(w_eco1329, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1330(w_eco1330, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1331(w_eco1331, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1332(w_eco1332, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1333(w_eco1333, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1334(w_eco1334, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1335(w_eco1335, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1336(w_eco1336, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1337(w_eco1337, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1338(w_eco1338, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1339(w_eco1339, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1340(w_eco1340, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1341(w_eco1341, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1342(w_eco1342, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1343(w_eco1343, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1344(w_eco1344, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1345(w_eco1345, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1346(w_eco1346, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1347(w_eco1347, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1348(w_eco1348, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1349(w_eco1349, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1350(w_eco1350, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1351(w_eco1351, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1352(w_eco1352, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1353(w_eco1353, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1354(w_eco1354, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1355(w_eco1355, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1356(w_eco1356, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1357(w_eco1357, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1358(w_eco1358, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1359(w_eco1359, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1360(w_eco1360, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1361(w_eco1361, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1362(w_eco1362, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1363(w_eco1363, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1364(w_eco1364, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1365(w_eco1365, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1366(w_eco1366, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1367(w_eco1367, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1368(w_eco1368, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1369(w_eco1369, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1370(w_eco1370, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1371(w_eco1371, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1372(w_eco1372, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1373(w_eco1373, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1374(w_eco1374, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1375(w_eco1375, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1376(w_eco1376, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1377(w_eco1377, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1378(w_eco1378, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1379(w_eco1379, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1380(w_eco1380, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1381(w_eco1381, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1382(w_eco1382, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1383(w_eco1383, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1384(w_eco1384, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1385(w_eco1385, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1386(w_eco1386, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1387(w_eco1387, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1388(w_eco1388, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1389(w_eco1389, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1390(w_eco1390, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1391(w_eco1391, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1392(w_eco1392, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1393(w_eco1393, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1394(w_eco1394, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1395(w_eco1395, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1396(w_eco1396, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1397(w_eco1397, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1398(w_eco1398, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1399(w_eco1399, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1400(w_eco1400, prev_cnt[2], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1401(w_eco1401, prev_cnt[4], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1402(w_eco1402, prev_cnt[0], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1403(w_eco1403, prev_cnt[5], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1404(w_eco1404, !Tgate[6], !Tgdel[6], prev_cnt[3], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1405(w_eco1405, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1406(w_eco1406, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1407(w_eco1407, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1408(w_eco1408, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1409(w_eco1409, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1410(w_eco1410, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1411(w_eco1411, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1412(w_eco1412, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1413(w_eco1413, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1414(w_eco1414, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1415(w_eco1415, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1416(w_eco1416, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1417(w_eco1417, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1418(w_eco1418, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1419(w_eco1419, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1420(w_eco1420, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1421(w_eco1421, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1422(w_eco1422, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1423(w_eco1423, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1424(w_eco1424, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1425(w_eco1425, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1426(w_eco1426, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1427(w_eco1427, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1428(w_eco1428, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1429(w_eco1429, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1430(w_eco1430, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1431(w_eco1431, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1432(w_eco1432, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1433(w_eco1433, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1434(w_eco1434, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1435(w_eco1435, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1436(w_eco1436, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1437(w_eco1437, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1438(w_eco1438, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1439(w_eco1439, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1440(w_eco1440, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1441(w_eco1441, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1442(w_eco1442, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1443(w_eco1443, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1444(w_eco1444, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1445(w_eco1445, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1446(w_eco1446, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1447(w_eco1447, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1448(w_eco1448, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1449(w_eco1449, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1450(w_eco1450, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1451(w_eco1451, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1452(w_eco1452, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1453(w_eco1453, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1454(w_eco1454, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1455(w_eco1455, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1456(w_eco1456, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1457(w_eco1457, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1458(w_eco1458, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1459(w_eco1459, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1460(w_eco1460, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1461(w_eco1461, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1462(w_eco1462, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1463(w_eco1463, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1464(w_eco1464, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1465(w_eco1465, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1466(w_eco1466, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1467(w_eco1467, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1468(w_eco1468, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1469(w_eco1469, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1470(w_eco1470, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1471(w_eco1471, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1472(w_eco1472, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1473(w_eco1473, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1474(w_eco1474, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1475(w_eco1475, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1476(w_eco1476, prev_cnt[4], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1477(w_eco1477, prev_cnt[0], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1478(w_eco1478, prev_cnt[5], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1479(w_eco1479, prev_cnt[3], !prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1480(w_eco1480, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1481(w_eco1481, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1482(w_eco1482, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1483(w_eco1483, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1484(w_eco1484, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1485(w_eco1485, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1486(w_eco1486, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1487(w_eco1487, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1488(w_eco1488, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1489(w_eco1489, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1490(w_eco1490, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1491(w_eco1491, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1492(w_eco1492, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1493(w_eco1493, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1494(w_eco1494, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1495(w_eco1495, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1496(w_eco1496, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1497(w_eco1497, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1498(w_eco1498, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1499(w_eco1499, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1500(w_eco1500, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1501(w_eco1501, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1502(w_eco1502, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1503(w_eco1503, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1504(w_eco1504, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1505(w_eco1505, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1506(w_eco1506, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1507(w_eco1507, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1508(w_eco1508, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1509(w_eco1509, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1510(w_eco1510, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1511(w_eco1511, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1512(w_eco1512, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1513(w_eco1513, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1514(w_eco1514, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1515(w_eco1515, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1516(w_eco1516, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1517(w_eco1517, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1518(w_eco1518, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1519(w_eco1519, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1520(w_eco1520, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1521(w_eco1521, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1522(w_eco1522, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1523(w_eco1523, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1524(w_eco1524, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1525(w_eco1525, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1526(w_eco1526, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1527(w_eco1527, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1528(w_eco1528, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1529(w_eco1529, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1530(w_eco1530, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1531(w_eco1531, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1532(w_eco1532, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1533(w_eco1533, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1534(w_eco1534, prev_cnt[0], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1535(w_eco1535, prev_cnt[5], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1536(w_eco1536, prev_cnt[3], !prev_cnt[6], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1537(w_eco1537, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1538(w_eco1538, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1539(w_eco1539, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1540(w_eco1540, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1541(w_eco1541, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1542(w_eco1542, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1543(w_eco1543, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1544(w_eco1544, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1545(w_eco1545, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1546(w_eco1546, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1547(w_eco1547, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1548(w_eco1548, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1549(w_eco1549, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1550(w_eco1550, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1551(w_eco1551, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1552(w_eco1552, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1553(w_eco1553, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1554(w_eco1554, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1555(w_eco1555, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1556(w_eco1556, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1557(w_eco1557, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1558(w_eco1558, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1559(w_eco1559, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1560(w_eco1560, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1561(w_eco1561, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1562(w_eco1562, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1563(w_eco1563, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1564(w_eco1564, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1565(w_eco1565, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1566(w_eco1566, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1567(w_eco1567, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1568(w_eco1568, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1569(w_eco1569, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1570(w_eco1570, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1571(w_eco1571, prev_cnt[5], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1572(w_eco1572, prev_cnt[3], !prev_cnt[6], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1573(w_eco1573, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1574(w_eco1574, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1575(w_eco1575, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1576(w_eco1576, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1577(w_eco1577, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1578(w_eco1578, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1579(w_eco1579, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1580(w_eco1580, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1581(w_eco1581, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1582(w_eco1582, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1583(w_eco1583, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1584(w_eco1584, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1585(w_eco1585, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1586(w_eco1586, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1587(w_eco1587, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1588(w_eco1588, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1589(w_eco1589, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1590(w_eco1590, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1591(w_eco1591, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1592(w_eco1592, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1593(w_eco1593, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1594(w_eco1594, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1595(w_eco1595, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1596(w_eco1596, prev_cnt[3], !prev_cnt[6], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1597(w_eco1597, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1598(w_eco1598, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1599(w_eco1599, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1600(w_eco1600, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1601(w_eco1601, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1602(w_eco1602, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1603(w_eco1603, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1604(w_eco1604, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1605(w_eco1605, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1606(w_eco1606, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1607(w_eco1607, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1608(w_eco1608, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1609(w_eco1609, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1610(w_eco1610, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1611(w_eco1611, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1612(w_eco1612, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1613(w_eco1613, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1614(w_eco1614, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1615(w_eco1615, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1616(w_eco1616, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1617(w_eco1617, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1618(w_eco1618, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1619(w_eco1619, !Tgate[6], !Tsync[6], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1620(w_eco1620, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1621(w_eco1621, !Tgate[6], !Tsync[6], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_1622(w_eco1622, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621);
	xor _ECO_out0(cnt[6], sub_wire0, w_eco1622);
	assign w_eco1623 = rst;
	assign w_eco1624 = prev_cnt[9];
	assign w_eco1625 = prev_cnt[15];
	assign w_eco1626 = prev_cnt[11];
	assign w_eco1627 = prev_cnt[6];
	assign w_eco1628 = prev_cnt[10];
	assign w_eco1629 = prev_cnt[8];
	and _ECO_1630(w_eco1630, !prev_cnt[14], prev_cnt[12]);
	and _ECO_1631(w_eco1631, !prev_cnt[14], prev_cnt[13]);
	and _ECO_1632(w_eco1632, ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1633(w_eco1633, ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_1634(w_eco1634, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7]);
	or _ECO_1635(w_eco1635, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634);
	xor _ECO_out1(Gate, sub_wire1, w_eco1635);
	assign w_eco1636 = rst;
	and _ECO_1637(w_eco1637, ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1638(w_eco1638, ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_1639(w_eco1639, !prev_cnt[2], ena, !prev_state[0]);
	and _ECO_1640(w_eco1640, !Tsync[2], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_1641(w_eco1641, !Tsync[2], !prev_cnt[2], ena, prev_state[3], !prev_state[2]);
	and _ECO_1642(w_eco1642, !Tsync[2], !prev_cnt[2], ena, prev_state[1]);
	and _ECO_1643(w_eco1643, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_1644(w_eco1644, !prev_cnt[2], ena, !prev_state[3], prev_state[1]);
	and _ECO_1645(w_eco1645, !Tsync[2], !prev_cnt[2], ena, prev_state[4], !prev_state[2]);
	and _ECO_1646(w_eco1646, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1647(w_eco1647, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_1648(w_eco1648, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1649(w_eco1649, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1650(w_eco1650, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1651(w_eco1651, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1652(w_eco1652, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1653(w_eco1653, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1654(w_eco1654, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1655(w_eco1655, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1656(w_eco1656, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1657(w_eco1657, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1658(w_eco1658, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1659(w_eco1659, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1660(w_eco1660, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1661(w_eco1661, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1662(w_eco1662, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1663(w_eco1663, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1664(w_eco1664, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1665(w_eco1665, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1666(w_eco1666, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1667(w_eco1667, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1668(w_eco1668, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1669(w_eco1669, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1670(w_eco1670, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1671(w_eco1671, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1672(w_eco1672, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1673(w_eco1673, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1674(w_eco1674, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1675(w_eco1675, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1676(w_eco1676, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1677(w_eco1677, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1678(w_eco1678, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1679(w_eco1679, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1680(w_eco1680, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1681(w_eco1681, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1682(w_eco1682, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1683(w_eco1683, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1684(w_eco1684, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1685(w_eco1685, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1686(w_eco1686, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1687(w_eco1687, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1688(w_eco1688, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1689(w_eco1689, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1690(w_eco1690, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1691(w_eco1691, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1692(w_eco1692, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1693(w_eco1693, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1694(w_eco1694, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1695(w_eco1695, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1696(w_eco1696, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1697(w_eco1697, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1698(w_eco1698, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1699(w_eco1699, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1700(w_eco1700, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1701(w_eco1701, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1702(w_eco1702, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1703(w_eco1703, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1704(w_eco1704, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1705(w_eco1705, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1706(w_eco1706, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1707(w_eco1707, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1708(w_eco1708, Tsync[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1709(w_eco1709, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1710(w_eco1710, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1711(w_eco1711, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1712(w_eco1712, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1713(w_eco1713, !Tsync[2], !prev_cnt[2], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1714(w_eco1714, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1715(w_eco1715, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1716(w_eco1716, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1717(w_eco1717, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1718(w_eco1718, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1719(w_eco1719, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1720(w_eco1720, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1721(w_eco1721, prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1722(w_eco1722, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1723(w_eco1723, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1724(w_eco1724, !Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1725(w_eco1725, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1726(w_eco1726, !Tsync[2], !prev_cnt[2], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1727(w_eco1727, prev_cnt[2], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1728(w_eco1728, !Tsync[2], !prev_cnt[2], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1729(w_eco1729, !Tsync[2], !prev_cnt[2], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1730(w_eco1730, !prev_cnt[2], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_1731(w_eco1731, !Tsync[2], !prev_cnt[2], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_1732(w_eco1732, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731);
	xor _ECO_out2(Sync, sub_wire2, w_eco1732);
	and _ECO_1733(w_eco1733, rst, prev_state[3], prev_state[0]);
	and _ECO_1734(w_eco1734, prev_cnt[1], prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1735(w_eco1735, Tsync[5], !rst, !prev_state[0]);
	and _ECO_1736(w_eco1736, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1737(w_eco1737, prev_cnt[1], prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1738(w_eco1738, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1739(w_eco1739, prev_cnt[1], prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1740(w_eco1740, prev_cnt[2], prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1741(w_eco1741, prev_cnt[1], prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1742(w_eco1742, prev_cnt[1], prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1743(w_eco1743, Tsync[5], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1744(w_eco1744, prev_cnt[1], prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1745(w_eco1745, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1746(w_eco1746, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1747(w_eco1747, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1748(w_eco1748, prev_cnt[2], prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1749(w_eco1749, Tgdel[5], prev_cnt[1], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1750(w_eco1750, prev_cnt[4], prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1751(w_eco1751, prev_cnt[2], prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1752(w_eco1752, prev_cnt[2], prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1753(w_eco1753, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1754(w_eco1754, Tsync[5], !ena, !rst, !prev_state[3]);
	and _ECO_1755(w_eco1755, prev_cnt[1], prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1756(w_eco1756, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1757(w_eco1757, prev_cnt[1], prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1758(w_eco1758, prev_cnt[2], prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1759(w_eco1759, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1760(w_eco1760, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1761(w_eco1761, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1762(w_eco1762, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1763(w_eco1763, prev_cnt[4], prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1764(w_eco1764, Tgdel[5], prev_cnt[2], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1765(w_eco1765, prev_cnt[0], prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1766(w_eco1766, prev_cnt[4], prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1767(w_eco1767, prev_cnt[4], prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1768(w_eco1768, prev_cnt[1], prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1769(w_eco1769, prev_cnt[4], prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1770(w_eco1770, prev_cnt[2], prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1771(w_eco1771, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1772(w_eco1772, prev_cnt[2], prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1773(w_eco1773, prev_cnt[2], prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1774(w_eco1774, Tgdel[5], prev_cnt[1], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1775(w_eco1775, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1776(w_eco1776, prev_cnt[2], prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1777(w_eco1777, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1778(w_eco1778, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_1779(w_eco1779, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1780(w_eco1780, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1781(w_eco1781, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1782(w_eco1782, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1783(w_eco1783, prev_cnt[0], prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1784(w_eco1784, Tgdel[5], prev_cnt[4], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1785(w_eco1785, prev_cnt[1], prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1786(w_eco1786, prev_cnt[3], prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1787(w_eco1787, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[9], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1788(w_eco1788, prev_cnt[0], prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1789(w_eco1789, prev_cnt[0], prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1790(w_eco1790, prev_cnt[0], prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1791(w_eco1791, prev_cnt[4], prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1792(w_eco1792, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1793(w_eco1793, prev_cnt[4], prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1794(w_eco1794, prev_cnt[4], prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1795(w_eco1795, Tgdel[5], prev_cnt[2], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1796(w_eco1796, prev_cnt[1], prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1797(w_eco1797, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1798(w_eco1798, prev_cnt[4], prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1799(w_eco1799, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1800(w_eco1800, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1801(w_eco1801, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1802(w_eco1802, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1803(w_eco1803, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1804(w_eco1804, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1805(w_eco1805, prev_cnt[3], prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1806(w_eco1806, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[9], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1807(w_eco1807, Tgdel[5], prev_cnt[0], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1808(w_eco1808, Tgate[5], prev_cnt[1], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1809(w_eco1809, prev_cnt[2], prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1810(w_eco1810, prev_cnt[3], prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1811(w_eco1811, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1812(w_eco1812, prev_cnt[3], prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1813(w_eco1813, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !ena, !rst, !prev_state[0]);
	and _ECO_1814(w_eco1814, prev_cnt[3], prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1815(w_eco1815, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[9], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1816(w_eco1816, prev_cnt[0], prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1817(w_eco1817, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1818(w_eco1818, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1819(w_eco1819, prev_cnt[0], prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1820(w_eco1820, prev_cnt[0], prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1821(w_eco1821, Tgdel[5], prev_cnt[4], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1822(w_eco1822, prev_cnt[1], prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1823(w_eco1823, prev_cnt[2], prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1824(w_eco1824, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1825(w_eco1825, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1826(w_eco1826, prev_cnt[0], prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1827(w_eco1827, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_1828(w_eco1828, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1829(w_eco1829, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1830(w_eco1830, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1831(w_eco1831, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1832(w_eco1832, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_1833(w_eco1833, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1834(w_eco1834, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1835(w_eco1835, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1836(w_eco1836, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1837(w_eco1837, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1838(w_eco1838, Tgdel[5], prev_cnt[3], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1839(w_eco1839, Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1840(w_eco1840, prev_cnt[1], prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1841(w_eco1841, Tgate[5], prev_cnt[2], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1842(w_eco1842, prev_cnt[4], prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1843(w_eco1843, prev_cnt[3], prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1844(w_eco1844, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1845(w_eco1845, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1846(w_eco1846, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1847(w_eco1847, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1848(w_eco1848, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1849(w_eco1849, prev_cnt[3], prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1850(w_eco1850, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !ena, !rst, !prev_state[3]);
	and _ECO_1851(w_eco1851, prev_cnt[3], prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1852(w_eco1852, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[9], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1853(w_eco1853, Tgdel[5], prev_cnt[0], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1854(w_eco1854, Tgate[5], prev_cnt[1], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1855(w_eco1855, prev_cnt[2], prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1856(w_eco1856, prev_cnt[4], prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1857(w_eco1857, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1858(w_eco1858, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1859(w_eco1859, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1860(w_eco1860, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1861(w_eco1861, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1862(w_eco1862, prev_cnt[3], prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1863(w_eco1863, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_1864(w_eco1864, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_1865(w_eco1865, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_1866(w_eco1866, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1867(w_eco1867, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1868(w_eco1868, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1869(w_eco1869, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_1870(w_eco1870, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1871(w_eco1871, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1872(w_eco1872, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1873(w_eco1873, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1874(w_eco1874, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1875(w_eco1875, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1876(w_eco1876, prev_cnt[1], prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1877(w_eco1877, prev_cnt[2], prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1878(w_eco1878, Tgate[5], prev_cnt[4], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1879(w_eco1879, prev_cnt[0], prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1880(w_eco1880, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1881(w_eco1881, Tgdel[5], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_1882(w_eco1882, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1883(w_eco1883, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1884(w_eco1884, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1885(w_eco1885, Tgdel[5], prev_cnt[3], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1886(w_eco1886, Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1887(w_eco1887, prev_cnt[1], prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1888(w_eco1888, Tgate[5], prev_cnt[2], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1889(w_eco1889, prev_cnt[4], prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1890(w_eco1890, prev_cnt[0], prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1891(w_eco1891, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1892(w_eco1892, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1893(w_eco1893, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1894(w_eco1894, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1895(w_eco1895, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1896(w_eco1896, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1897(w_eco1897, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_1898(w_eco1898, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_1899(w_eco1899, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_1900(w_eco1900, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_1901(w_eco1901, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_1902(w_eco1902, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1903(w_eco1903, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1904(w_eco1904, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_1905(w_eco1905, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_1906(w_eco1906, Tgdel[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !ena, !rst, !prev_state[0]);
	and _ECO_1907(w_eco1907, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1908(w_eco1908, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1909(w_eco1909, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1910(w_eco1910, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1911(w_eco1911, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1912(w_eco1912, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1913(w_eco1913, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1914(w_eco1914, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1915(w_eco1915, Tgdel[5], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_1916(w_eco1916, prev_cnt[1], prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1917(w_eco1917, prev_cnt[2], prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1918(w_eco1918, prev_cnt[4], prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1919(w_eco1919, Tgate[5], prev_cnt[0], prev_cnt[5], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1920(w_eco1920, prev_cnt[3], prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1921(w_eco1921, Tgdel[5], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_1922(w_eco1922, prev_cnt[14], prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1923(w_eco1923, Tgdel[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_1924(w_eco1924, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1925(w_eco1925, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1926(w_eco1926, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1927(w_eco1927, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1928(w_eco1928, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1929(w_eco1929, prev_cnt[1], prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1930(w_eco1930, prev_cnt[2], prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1931(w_eco1931, Tgate[5], prev_cnt[4], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1932(w_eco1932, prev_cnt[0], prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1933(w_eco1933, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1934(w_eco1934, prev_cnt[3], prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1935(w_eco1935, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_1936(w_eco1936, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1937(w_eco1937, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1938(w_eco1938, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1939(w_eco1939, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1940(w_eco1940, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1941(w_eco1941, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1942(w_eco1942, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1943(w_eco1943, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1944(w_eco1944, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1945(w_eco1945, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_1946(w_eco1946, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_1947(w_eco1947, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_1948(w_eco1948, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_1949(w_eco1949, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_1950(w_eco1950, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1951(w_eco1951, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_1952(w_eco1952, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_1953(w_eco1953, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_1954(w_eco1954, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1955(w_eco1955, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1956(w_eco1956, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1957(w_eco1957, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1958(w_eco1958, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1959(w_eco1959, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1960(w_eco1960, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1961(w_eco1961, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1962(w_eco1962, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1963(w_eco1963, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_1964(w_eco1964, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_1965(w_eco1965, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1966(w_eco1966, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_1967(w_eco1967, prev_cnt[1], prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1968(w_eco1968, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1969(w_eco1969, prev_cnt[2], prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1970(w_eco1970, prev_cnt[4], prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1971(w_eco1971, prev_cnt[0], prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1972(w_eco1972, prev_cnt[3], prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1973(w_eco1973, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_1974(w_eco1974, Tgdel[5], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_1975(w_eco1975, Tgdel[5], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_1976(w_eco1976, prev_cnt[14], prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_1977(w_eco1977, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !ena, !rst, !prev_state[0]);
	and _ECO_1978(w_eco1978, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[3], prev_state[1]);
	and _ECO_1979(w_eco1979, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1980(w_eco1980, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1981(w_eco1981, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1982(w_eco1982, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1983(w_eco1983, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1984(w_eco1984, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_1985(w_eco1985, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1986(w_eco1986, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_1987(w_eco1987, Tgdel[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !ena, !rst, !prev_state[3]);
	and _ECO_1988(w_eco1988, prev_cnt[1], prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1989(w_eco1989, prev_cnt[2], prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1990(w_eco1990, prev_cnt[4], prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1991(w_eco1991, Tgate[5], prev_cnt[0], prev_cnt[5], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1992(w_eco1992, prev_cnt[3], prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_1993(w_eco1993, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1994(w_eco1994, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1995(w_eco1995, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1996(w_eco1996, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1997(w_eco1997, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1998(w_eco1998, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_1999(w_eco1999, prev_cnt[1], prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2000(w_eco2000, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2001(w_eco2001, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2002(w_eco2002, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2003(w_eco2003, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2004(w_eco2004, prev_cnt[14], prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2005(w_eco2005, Tgdel[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_2006(w_eco2006, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2007(w_eco2007, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2008(w_eco2008, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2009(w_eco2009, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_2010(w_eco2010, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_2011(w_eco2011, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_2012(w_eco2012, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_2013(w_eco2013, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_2014(w_eco2014, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_2015(w_eco2015, Tgdel[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !ena, !rst, !prev_state[0]);
	and _ECO_2016(w_eco2016, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2017(w_eco2017, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2018(w_eco2018, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2019(w_eco2019, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2020(w_eco2020, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2021(w_eco2021, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2022(w_eco2022, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2023(w_eco2023, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2024(w_eco2024, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2025(w_eco2025, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2026(w_eco2026, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2027(w_eco2027, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2028(w_eco2028, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2029(w_eco2029, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2030(w_eco2030, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2031(w_eco2031, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2032(w_eco2032, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2033(w_eco2033, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2034(w_eco2034, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2035(w_eco2035, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2036(w_eco2036, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2037(w_eco2037, prev_cnt[2], prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2038(w_eco2038, prev_cnt[4], prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2039(w_eco2039, prev_cnt[0], prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2040(w_eco2040, prev_cnt[3], prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2041(w_eco2041, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[11], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2042(w_eco2042, Tgdel[5], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2043(w_eco2043, Tgdel[5], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2044(w_eco2044, Tgdel[5], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2045(w_eco2045, Tgdel[5], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2046(w_eco2046, prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2047(w_eco2047, prev_cnt[14], prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2048(w_eco2048, Tgdel[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_2049(w_eco2049, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2050(w_eco2050, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2051(w_eco2051, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2052(w_eco2052, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2053(w_eco2053, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2054(w_eco2054, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2055(w_eco2055, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2056(w_eco2056, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2057(w_eco2057, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2058(w_eco2058, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2059(w_eco2059, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2060(w_eco2060, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !ena, !rst, !prev_state[3]);
	and _ECO_2061(w_eco2061, prev_cnt[1], prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2062(w_eco2062, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2063(w_eco2063, prev_cnt[2], prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2064(w_eco2064, prev_cnt[4], prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2065(w_eco2065, prev_cnt[0], prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2066(w_eco2066, prev_cnt[3], prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2067(w_eco2067, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2068(w_eco2068, Tgdel[5], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2069(w_eco2069, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2070(w_eco2070, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2071(w_eco2071, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2072(w_eco2072, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2073(w_eco2073, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2074(w_eco2074, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2075(w_eco2075, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2076(w_eco2076, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2077(w_eco2077, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2078(w_eco2078, prev_cnt[1], prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2079(w_eco2079, prev_cnt[2], prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2080(w_eco2080, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2081(w_eco2081, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2082(w_eco2082, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2083(w_eco2083, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2084(w_eco2084, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2085(w_eco2085, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2086(w_eco2086, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2087(w_eco2087, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2088(w_eco2088, prev_cnt[14], prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2089(w_eco2089, Tgate[5], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_2090(w_eco2090, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2091(w_eco2091, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_2092(w_eco2092, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_2093(w_eco2093, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_2094(w_eco2094, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_2095(w_eco2095, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_2096(w_eco2096, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2097(w_eco2097, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2098(w_eco2098, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2099(w_eco2099, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2100(w_eco2100, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2101(w_eco2101, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2102(w_eco2102, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2103(w_eco2103, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2104(w_eco2104, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2105(w_eco2105, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2106(w_eco2106, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2107(w_eco2107, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2108(w_eco2108, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2109(w_eco2109, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2110(w_eco2110, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2111(w_eco2111, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2112(w_eco2112, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2113(w_eco2113, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2114(w_eco2114, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2115(w_eco2115, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2116(w_eco2116, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2117(w_eco2117, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2118(w_eco2118, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2119(w_eco2119, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2120(w_eco2120, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2121(w_eco2121, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2122(w_eco2122, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2123(w_eco2123, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2124(w_eco2124, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2125(w_eco2125, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2126(w_eco2126, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2127(w_eco2127, prev_cnt[4], prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2128(w_eco2128, prev_cnt[0], prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2129(w_eco2129, prev_cnt[3], prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2130(w_eco2130, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2131(w_eco2131, Tgdel[5], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2132(w_eco2132, Tgdel[5], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2133(w_eco2133, Tgdel[5], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2134(w_eco2134, prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2135(w_eco2135, prev_cnt[14], prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2136(w_eco2136, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !ena, !rst, !prev_state[0]);
	and _ECO_2137(w_eco2137, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[3], prev_state[1]);
	and _ECO_2138(w_eco2138, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2139(w_eco2139, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2140(w_eco2140, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2141(w_eco2141, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2142(w_eco2142, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2143(w_eco2143, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2144(w_eco2144, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2145(w_eco2145, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2146(w_eco2146, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2147(w_eco2147, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2148(w_eco2148, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2149(w_eco2149, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2150(w_eco2150, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2151(w_eco2151, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2152(w_eco2152, Tgdel[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !ena, !rst, !prev_state[3]);
	and _ECO_2153(w_eco2153, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2154(w_eco2154, prev_cnt[2], prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2155(w_eco2155, prev_cnt[4], prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2156(w_eco2156, prev_cnt[0], prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2157(w_eco2157, prev_cnt[3], prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2158(w_eco2158, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[11], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2159(w_eco2159, Tgdel[5], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2160(w_eco2160, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2161(w_eco2161, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2162(w_eco2162, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2163(w_eco2163, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2164(w_eco2164, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2165(w_eco2165, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2166(w_eco2166, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2167(w_eco2167, prev_cnt[1], prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2168(w_eco2168, prev_cnt[2], prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2169(w_eco2169, prev_cnt[4], prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2170(w_eco2170, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2171(w_eco2171, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2172(w_eco2172, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2173(w_eco2173, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2174(w_eco2174, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2175(w_eco2175, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2176(w_eco2176, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2177(w_eco2177, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2178(w_eco2178, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2179(w_eco2179, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2180(w_eco2180, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2181(w_eco2181, prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2182(w_eco2182, prev_cnt[14], prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2183(w_eco2183, Tgdel[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_2184(w_eco2184, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2185(w_eco2185, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2186(w_eco2186, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_2187(w_eco2187, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_2188(w_eco2188, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_2189(w_eco2189, !Tgate[5], !Tgdel[5], !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_2190(w_eco2190, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_state[3], prev_state[0]);
	and _ECO_2191(w_eco2191, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2192(w_eco2192, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2193(w_eco2193, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2194(w_eco2194, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2195(w_eco2195, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2196(w_eco2196, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2197(w_eco2197, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2198(w_eco2198, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2199(w_eco2199, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2200(w_eco2200, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2201(w_eco2201, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2202(w_eco2202, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2203(w_eco2203, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2204(w_eco2204, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2205(w_eco2205, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2206(w_eco2206, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2207(w_eco2207, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2208(w_eco2208, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2209(w_eco2209, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2210(w_eco2210, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2211(w_eco2211, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2212(w_eco2212, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2213(w_eco2213, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2214(w_eco2214, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2215(w_eco2215, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2216(w_eco2216, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2217(w_eco2217, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2218(w_eco2218, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2219(w_eco2219, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2220(w_eco2220, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2221(w_eco2221, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2222(w_eco2222, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2223(w_eco2223, prev_cnt[0], prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2224(w_eco2224, prev_cnt[3], prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2225(w_eco2225, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[10], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2226(w_eco2226, Tgdel[5], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2227(w_eco2227, Tgdel[5], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2228(w_eco2228, Tgdel[5], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2229(w_eco2229, Tgdel[5], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2230(w_eco2230, prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2231(w_eco2231, prev_cnt[14], prev_cnt[3], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2232(w_eco2232, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2233(w_eco2233, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2234(w_eco2234, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2235(w_eco2235, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2236(w_eco2236, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2237(w_eco2237, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2238(w_eco2238, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2239(w_eco2239, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2240(w_eco2240, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2241(w_eco2241, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2242(w_eco2242, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2243(w_eco2243, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2244(w_eco2244, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2245(w_eco2245, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2246(w_eco2246, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2247(w_eco2247, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2248(w_eco2248, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2249(w_eco2249, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2250(w_eco2250, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2251(w_eco2251, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !ena, !rst, !prev_state[3]);
	and _ECO_2252(w_eco2252, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2253(w_eco2253, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2254(w_eco2254, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2255(w_eco2255, prev_cnt[4], prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2256(w_eco2256, prev_cnt[0], prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2257(w_eco2257, prev_cnt[3], prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2258(w_eco2258, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2259(w_eco2259, Tgdel[5], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2260(w_eco2260, Tgdel[5], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2261(w_eco2261, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2262(w_eco2262, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2263(w_eco2263, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2264(w_eco2264, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2265(w_eco2265, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2266(w_eco2266, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2267(w_eco2267, prev_cnt[0], prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2268(w_eco2268, prev_cnt[1], prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2269(w_eco2269, prev_cnt[2], prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2270(w_eco2270, prev_cnt[4], prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2271(w_eco2271, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2272(w_eco2272, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2273(w_eco2273, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2274(w_eco2274, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2275(w_eco2275, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2276(w_eco2276, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2277(w_eco2277, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2278(w_eco2278, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2279(w_eco2279, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2280(w_eco2280, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2281(w_eco2281, prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2282(w_eco2282, prev_cnt[14], prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2283(w_eco2283, Tgate[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_2284(w_eco2284, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2285(w_eco2285, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2286(w_eco2286, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2287(w_eco2287, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_2288(w_eco2288, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_2289(w_eco2289, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2290(w_eco2290, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2291(w_eco2291, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2292(w_eco2292, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2293(w_eco2293, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2294(w_eco2294, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2295(w_eco2295, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2296(w_eco2296, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2297(w_eco2297, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2298(w_eco2298, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2299(w_eco2299, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2300(w_eco2300, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2301(w_eco2301, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2302(w_eco2302, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2303(w_eco2303, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2304(w_eco2304, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2305(w_eco2305, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2306(w_eco2306, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2307(w_eco2307, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2308(w_eco2308, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2309(w_eco2309, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2310(w_eco2310, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2311(w_eco2311, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2312(w_eco2312, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2313(w_eco2313, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2314(w_eco2314, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2315(w_eco2315, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2316(w_eco2316, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2317(w_eco2317, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2318(w_eco2318, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2319(w_eco2319, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2320(w_eco2320, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2321(w_eco2321, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2322(w_eco2322, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2323(w_eco2323, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2324(w_eco2324, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2325(w_eco2325, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2326(w_eco2326, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2327(w_eco2327, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2328(w_eco2328, prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2329(w_eco2329, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2330(w_eco2330, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2331(w_eco2331, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2332(w_eco2332, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[8], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2333(w_eco2333, Tgdel[5], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2334(w_eco2334, Tgdel[5], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2335(w_eco2335, Tgdel[5], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2336(w_eco2336, Tgdel[5], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2337(w_eco2337, prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2338(w_eco2338, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2339(w_eco2339, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2340(w_eco2340, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2341(w_eco2341, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2342(w_eco2342, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2343(w_eco2343, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2344(w_eco2344, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2345(w_eco2345, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2346(w_eco2346, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2347(w_eco2347, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2348(w_eco2348, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2349(w_eco2349, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2350(w_eco2350, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2351(w_eco2351, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2352(w_eco2352, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2353(w_eco2353, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2354(w_eco2354, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2355(w_eco2355, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2356(w_eco2356, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2357(w_eco2357, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2358(w_eco2358, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2359(w_eco2359, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2360(w_eco2360, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2361(w_eco2361, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2362(w_eco2362, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2363(w_eco2363, prev_cnt[0], prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2364(w_eco2364, prev_cnt[3], prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2365(w_eco2365, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[10], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2366(w_eco2366, Tgdel[5], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2367(w_eco2367, Tgdel[5], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2368(w_eco2368, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2369(w_eco2369, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2370(w_eco2370, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2371(w_eco2371, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2372(w_eco2372, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2373(w_eco2373, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2374(w_eco2374, prev_cnt[3], prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2375(w_eco2375, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[15], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2376(w_eco2376, prev_cnt[1], prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2377(w_eco2377, prev_cnt[2], prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2378(w_eco2378, prev_cnt[4], prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2379(w_eco2379, prev_cnt[0], prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2380(w_eco2380, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2381(w_eco2381, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2382(w_eco2382, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2383(w_eco2383, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2384(w_eco2384, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2385(w_eco2385, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2386(w_eco2386, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2387(w_eco2387, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2388(w_eco2388, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2389(w_eco2389, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2390(w_eco2390, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2391(w_eco2391, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2392(w_eco2392, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2393(w_eco2393, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2394(w_eco2394, prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2395(w_eco2395, prev_cnt[14], prev_cnt[3], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2396(w_eco2396, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2397(w_eco2397, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2398(w_eco2398, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2399(w_eco2399, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2400(w_eco2400, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2401(w_eco2401, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2402(w_eco2402, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2403(w_eco2403, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2404(w_eco2404, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2405(w_eco2405, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2406(w_eco2406, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2407(w_eco2407, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2408(w_eco2408, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2409(w_eco2409, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2410(w_eco2410, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2411(w_eco2411, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2412(w_eco2412, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2413(w_eco2413, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2414(w_eco2414, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2415(w_eco2415, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2416(w_eco2416, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2417(w_eco2417, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2418(w_eco2418, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2419(w_eco2419, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2420(w_eco2420, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2421(w_eco2421, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2422(w_eco2422, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2423(w_eco2423, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2424(w_eco2424, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2425(w_eco2425, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2426(w_eco2426, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2427(w_eco2427, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2428(w_eco2428, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2429(w_eco2429, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2430(w_eco2430, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2431(w_eco2431, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2432(w_eco2432, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2433(w_eco2433, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2434(w_eco2434, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2435(w_eco2435, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2436(w_eco2436, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2437(w_eco2437, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2438(w_eco2438, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2439(w_eco2439, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2440(w_eco2440, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2441(w_eco2441, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2442(w_eco2442, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2443(w_eco2443, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2444(w_eco2444, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2445(w_eco2445, prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2446(w_eco2446, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2447(w_eco2447, Tgdel[5], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2448(w_eco2448, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2449(w_eco2449, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2450(w_eco2450, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[12], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2451(w_eco2451, Tgdel[5], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2452(w_eco2452, Tgdel[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2453(w_eco2453, prev_cnt[3], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2454(w_eco2454, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2455(w_eco2455, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2456(w_eco2456, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2457(w_eco2457, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2458(w_eco2458, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2459(w_eco2459, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2460(w_eco2460, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2461(w_eco2461, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2462(w_eco2462, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2463(w_eco2463, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2464(w_eco2464, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2465(w_eco2465, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2466(w_eco2466, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2467(w_eco2467, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2468(w_eco2468, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2469(w_eco2469, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2470(w_eco2470, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2471(w_eco2471, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2472(w_eco2472, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2473(w_eco2473, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2474(w_eco2474, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2475(w_eco2475, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2476(w_eco2476, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2477(w_eco2477, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2478(w_eco2478, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2479(w_eco2479, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2480(w_eco2480, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2481(w_eco2481, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2482(w_eco2482, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2483(w_eco2483, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2484(w_eco2484, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2485(w_eco2485, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2486(w_eco2486, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2487(w_eco2487, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[8], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2488(w_eco2488, Tgdel[5], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2489(w_eco2489, Tgdel[5], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2490(w_eco2490, Tgdel[5], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2491(w_eco2491, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2492(w_eco2492, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2493(w_eco2493, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2494(w_eco2494, !Tgate[5], !Tgdel[5], !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2495(w_eco2495, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2496(w_eco2496, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2497(w_eco2497, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2498(w_eco2498, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2499(w_eco2499, prev_cnt[2], prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2500(w_eco2500, prev_cnt[4], prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2501(w_eco2501, prev_cnt[0], prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2502(w_eco2502, prev_cnt[3], prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2503(w_eco2503, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2504(w_eco2504, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2505(w_eco2505, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2506(w_eco2506, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2507(w_eco2507, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2508(w_eco2508, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2509(w_eco2509, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2510(w_eco2510, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2511(w_eco2511, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2512(w_eco2512, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2513(w_eco2513, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2514(w_eco2514, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2515(w_eco2515, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2516(w_eco2516, !Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2517(w_eco2517, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2518(w_eco2518, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2519(w_eco2519, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2520(w_eco2520, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2521(w_eco2521, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2522(w_eco2522, prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2523(w_eco2523, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2524(w_eco2524, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2525(w_eco2525, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2526(w_eco2526, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_2527(w_eco2527, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2528(w_eco2528, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2529(w_eco2529, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2530(w_eco2530, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2531(w_eco2531, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2532(w_eco2532, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2533(w_eco2533, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2534(w_eco2534, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2535(w_eco2535, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2536(w_eco2536, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2537(w_eco2537, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2538(w_eco2538, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2539(w_eco2539, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2540(w_eco2540, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2541(w_eco2541, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2542(w_eco2542, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2543(w_eco2543, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2544(w_eco2544, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2545(w_eco2545, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2546(w_eco2546, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2547(w_eco2547, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2548(w_eco2548, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2549(w_eco2549, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2550(w_eco2550, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2551(w_eco2551, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2552(w_eco2552, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2553(w_eco2553, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2554(w_eco2554, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2555(w_eco2555, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2556(w_eco2556, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2557(w_eco2557, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2558(w_eco2558, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2559(w_eco2559, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2560(w_eco2560, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2561(w_eco2561, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2562(w_eco2562, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2563(w_eco2563, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2564(w_eco2564, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2565(w_eco2565, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2566(w_eco2566, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2567(w_eco2567, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2568(w_eco2568, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2569(w_eco2569, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2570(w_eco2570, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2571(w_eco2571, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2572(w_eco2572, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2573(w_eco2573, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2574(w_eco2574, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2575(w_eco2575, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2576(w_eco2576, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2577(w_eco2577, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2578(w_eco2578, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2579(w_eco2579, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2580(w_eco2580, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2581(w_eco2581, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2582(w_eco2582, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2583(w_eco2583, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2584(w_eco2584, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2585(w_eco2585, prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2586(w_eco2586, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2587(w_eco2587, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2588(w_eco2588, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[13], !rst, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_2589(w_eco2589, Tgdel[5], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2590(w_eco2590, Tgdel[5], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_2591(w_eco2591, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_2592(w_eco2592, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2593(w_eco2593, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_2594(w_eco2594, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2595(w_eco2595, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2596(w_eco2596, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2597(w_eco2597, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2598(w_eco2598, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2599(w_eco2599, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2600(w_eco2600, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2601(w_eco2601, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2602(w_eco2602, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2603(w_eco2603, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2604(w_eco2604, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2605(w_eco2605, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2606(w_eco2606, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2607(w_eco2607, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2608(w_eco2608, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2609(w_eco2609, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2610(w_eco2610, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2611(w_eco2611, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2612(w_eco2612, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2613(w_eco2613, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2614(w_eco2614, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2615(w_eco2615, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2616(w_eco2616, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2617(w_eco2617, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2618(w_eco2618, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2619(w_eco2619, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2620(w_eco2620, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2621(w_eco2621, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2622(w_eco2622, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2623(w_eco2623, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2624(w_eco2624, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2625(w_eco2625, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2626(w_eco2626, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2627(w_eco2627, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2628(w_eco2628, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2629(w_eco2629, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[12], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2630(w_eco2630, Tgdel[5], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2631(w_eco2631, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2632(w_eco2632, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_2633(w_eco2633, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2634(w_eco2634, !prev_cnt[14], prev_cnt[1], prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2635(w_eco2635, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2636(w_eco2636, prev_cnt[4], prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2637(w_eco2637, prev_cnt[0], prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2638(w_eco2638, prev_cnt[3], prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2639(w_eco2639, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[11], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2640(w_eco2640, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2641(w_eco2641, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2642(w_eco2642, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2643(w_eco2643, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2644(w_eco2644, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2645(w_eco2645, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2646(w_eco2646, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2647(w_eco2647, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2648(w_eco2648, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2649(w_eco2649, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2650(w_eco2650, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2651(w_eco2651, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2652(w_eco2652, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2653(w_eco2653, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2654(w_eco2654, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2655(w_eco2655, !Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2656(w_eco2656, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2657(w_eco2657, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2658(w_eco2658, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2659(w_eco2659, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2660(w_eco2660, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2661(w_eco2661, prev_cnt[3], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2662(w_eco2662, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2663(w_eco2663, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2664(w_eco2664, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2665(w_eco2665, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2666(w_eco2666, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2667(w_eco2667, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2668(w_eco2668, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2669(w_eco2669, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2670(w_eco2670, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2671(w_eco2671, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2672(w_eco2672, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2673(w_eco2673, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2674(w_eco2674, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2675(w_eco2675, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2676(w_eco2676, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2677(w_eco2677, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2678(w_eco2678, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2679(w_eco2679, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2680(w_eco2680, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2681(w_eco2681, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2682(w_eco2682, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2683(w_eco2683, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2684(w_eco2684, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2685(w_eco2685, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2686(w_eco2686, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2687(w_eco2687, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2688(w_eco2688, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2689(w_eco2689, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2690(w_eco2690, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2691(w_eco2691, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2692(w_eco2692, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2693(w_eco2693, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2694(w_eco2694, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2695(w_eco2695, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2696(w_eco2696, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2697(w_eco2697, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2698(w_eco2698, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2699(w_eco2699, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2700(w_eco2700, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2701(w_eco2701, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2702(w_eco2702, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2703(w_eco2703, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2704(w_eco2704, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2705(w_eco2705, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2706(w_eco2706, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2707(w_eco2707, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2708(w_eco2708, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2709(w_eco2709, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2710(w_eco2710, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2711(w_eco2711, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2712(w_eco2712, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2713(w_eco2713, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2714(w_eco2714, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2715(w_eco2715, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2716(w_eco2716, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2717(w_eco2717, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2718(w_eco2718, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2719(w_eco2719, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2720(w_eco2720, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2721(w_eco2721, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2722(w_eco2722, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2723(w_eco2723, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2724(w_eco2724, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2725(w_eco2725, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2726(w_eco2726, prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2727(w_eco2727, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2728(w_eco2728, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2729(w_eco2729, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2730(w_eco2730, prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2731(w_eco2731, Tgdel[5], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[1], !prev_state[0]);
	and _ECO_2732(w_eco2732, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2733(w_eco2733, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2734(w_eco2734, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2735(w_eco2735, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2736(w_eco2736, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2737(w_eco2737, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2738(w_eco2738, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2739(w_eco2739, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2740(w_eco2740, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2741(w_eco2741, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2742(w_eco2742, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2743(w_eco2743, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2744(w_eco2744, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2745(w_eco2745, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2746(w_eco2746, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2747(w_eco2747, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2748(w_eco2748, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2749(w_eco2749, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2750(w_eco2750, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2751(w_eco2751, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2752(w_eco2752, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2753(w_eco2753, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2754(w_eco2754, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2755(w_eco2755, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2756(w_eco2756, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2757(w_eco2757, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2758(w_eco2758, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2759(w_eco2759, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2760(w_eco2760, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2761(w_eco2761, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2762(w_eco2762, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2763(w_eco2763, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2764(w_eco2764, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2765(w_eco2765, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2766(w_eco2766, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2767(w_eco2767, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2768(w_eco2768, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2769(w_eco2769, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2770(w_eco2770, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2771(w_eco2771, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2772(w_eco2772, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2773(w_eco2773, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2774(w_eco2774, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2775(w_eco2775, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[13], !rst, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_2776(w_eco2776, Tgdel[5], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2777(w_eco2777, Tgdel[5], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_2778(w_eco2778, !prev_cnt[14], prev_cnt[2], prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2779(w_eco2779, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2780(w_eco2780, prev_cnt[0], prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2781(w_eco2781, prev_cnt[3], prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2782(w_eco2782, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[6], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2783(w_eco2783, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2784(w_eco2784, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2785(w_eco2785, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2786(w_eco2786, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2787(w_eco2787, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2788(w_eco2788, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2789(w_eco2789, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2790(w_eco2790, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2791(w_eco2791, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2792(w_eco2792, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2793(w_eco2793, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2794(w_eco2794, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2795(w_eco2795, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2796(w_eco2796, !Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2797(w_eco2797, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2798(w_eco2798, !Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2799(w_eco2799, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2800(w_eco2800, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2801(w_eco2801, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2802(w_eco2802, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2803(w_eco2803, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_2804(w_eco2804, Tsync[5], !rst, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_2805(w_eco2805, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2806(w_eco2806, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2807(w_eco2807, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2808(w_eco2808, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2809(w_eco2809, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2810(w_eco2810, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2811(w_eco2811, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2812(w_eco2812, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2813(w_eco2813, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2814(w_eco2814, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2815(w_eco2815, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2816(w_eco2816, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2817(w_eco2817, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2818(w_eco2818, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2819(w_eco2819, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2820(w_eco2820, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2821(w_eco2821, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2822(w_eco2822, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2823(w_eco2823, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2824(w_eco2824, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2825(w_eco2825, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2826(w_eco2826, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2827(w_eco2827, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2828(w_eco2828, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2829(w_eco2829, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2830(w_eco2830, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2831(w_eco2831, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2832(w_eco2832, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2833(w_eco2833, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2834(w_eco2834, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2835(w_eco2835, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2836(w_eco2836, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2837(w_eco2837, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2838(w_eco2838, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2839(w_eco2839, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2840(w_eco2840, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2841(w_eco2841, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2842(w_eco2842, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2843(w_eco2843, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2844(w_eco2844, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2845(w_eco2845, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2846(w_eco2846, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2847(w_eco2847, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2848(w_eco2848, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2849(w_eco2849, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2850(w_eco2850, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2851(w_eco2851, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2852(w_eco2852, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2853(w_eco2853, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2854(w_eco2854, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2855(w_eco2855, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2856(w_eco2856, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2857(w_eco2857, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2858(w_eco2858, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2859(w_eco2859, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2860(w_eco2860, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2861(w_eco2861, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2862(w_eco2862, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2863(w_eco2863, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2864(w_eco2864, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2865(w_eco2865, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2866(w_eco2866, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2867(w_eco2867, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2868(w_eco2868, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2869(w_eco2869, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2870(w_eco2870, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2871(w_eco2871, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2872(w_eco2872, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2873(w_eco2873, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2874(w_eco2874, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2875(w_eco2875, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2876(w_eco2876, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2877(w_eco2877, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2878(w_eco2878, prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2879(w_eco2879, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2880(w_eco2880, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2881(w_eco2881, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2882(w_eco2882, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2883(w_eco2883, prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2884(w_eco2884, prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2885(w_eco2885, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2886(w_eco2886, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2887(w_eco2887, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2888(w_eco2888, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2889(w_eco2889, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2890(w_eco2890, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2891(w_eco2891, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2892(w_eco2892, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2893(w_eco2893, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2894(w_eco2894, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2895(w_eco2895, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2896(w_eco2896, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2897(w_eco2897, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2898(w_eco2898, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2899(w_eco2899, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2900(w_eco2900, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2901(w_eco2901, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2902(w_eco2902, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2903(w_eco2903, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2904(w_eco2904, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2905(w_eco2905, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2906(w_eco2906, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2907(w_eco2907, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2908(w_eco2908, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2909(w_eco2909, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2910(w_eco2910, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2911(w_eco2911, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2912(w_eco2912, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2913(w_eco2913, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2914(w_eco2914, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2915(w_eco2915, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2916(w_eco2916, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2917(w_eco2917, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2918(w_eco2918, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2919(w_eco2919, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2920(w_eco2920, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2921(w_eco2921, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2922(w_eco2922, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2923(w_eco2923, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2924(w_eco2924, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2925(w_eco2925, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2926(w_eco2926, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2927(w_eco2927, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2928(w_eco2928, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2929(w_eco2929, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2930(w_eco2930, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2931(w_eco2931, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2932(w_eco2932, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2933(w_eco2933, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2934(w_eco2934, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2935(w_eco2935, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2936(w_eco2936, !prev_cnt[14], prev_cnt[4], prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2937(w_eco2937, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2938(w_eco2938, prev_cnt[3], prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2939(w_eco2939, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[10], !rst, prev_state[1], !prev_state[0]);
	and _ECO_2940(w_eco2940, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2941(w_eco2941, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2942(w_eco2942, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2943(w_eco2943, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2944(w_eco2944, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2945(w_eco2945, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2946(w_eco2946, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2947(w_eco2947, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2948(w_eco2948, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2949(w_eco2949, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2950(w_eco2950, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2951(w_eco2951, !Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2952(w_eco2952, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2953(w_eco2953, !Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2954(w_eco2954, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2955(w_eco2955, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2956(w_eco2956, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_2957(w_eco2957, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2958(w_eco2958, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2959(w_eco2959, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2960(w_eco2960, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2961(w_eco2961, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2962(w_eco2962, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2963(w_eco2963, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2964(w_eco2964, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2965(w_eco2965, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2966(w_eco2966, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2967(w_eco2967, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2968(w_eco2968, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2969(w_eco2969, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2970(w_eco2970, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2971(w_eco2971, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2972(w_eco2972, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2973(w_eco2973, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2974(w_eco2974, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2975(w_eco2975, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2976(w_eco2976, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2977(w_eco2977, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2978(w_eco2978, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2979(w_eco2979, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2980(w_eco2980, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2981(w_eco2981, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2982(w_eco2982, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2983(w_eco2983, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2984(w_eco2984, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2985(w_eco2985, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2986(w_eco2986, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_2987(w_eco2987, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2988(w_eco2988, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2989(w_eco2989, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2990(w_eco2990, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2991(w_eco2991, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2992(w_eco2992, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_2993(w_eco2993, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2994(w_eco2994, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2995(w_eco2995, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2996(w_eco2996, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2997(w_eco2997, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_2998(w_eco2998, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_2999(w_eco2999, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3000(w_eco3000, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3001(w_eco3001, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3002(w_eco3002, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3003(w_eco3003, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3004(w_eco3004, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3005(w_eco3005, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3006(w_eco3006, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3007(w_eco3007, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3008(w_eco3008, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3009(w_eco3009, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3010(w_eco3010, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3011(w_eco3011, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3012(w_eco3012, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3013(w_eco3013, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3014(w_eco3014, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3015(w_eco3015, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3016(w_eco3016, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3017(w_eco3017, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3018(w_eco3018, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3019(w_eco3019, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3020(w_eco3020, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3021(w_eco3021, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3022(w_eco3022, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3023(w_eco3023, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3024(w_eco3024, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3025(w_eco3025, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3026(w_eco3026, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3027(w_eco3027, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3028(w_eco3028, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3029(w_eco3029, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3030(w_eco3030, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3031(w_eco3031, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3032(w_eco3032, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3033(w_eco3033, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3034(w_eco3034, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3035(w_eco3035, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3036(w_eco3036, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3037(w_eco3037, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3038(w_eco3038, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3039(w_eco3039, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3040(w_eco3040, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3041(w_eco3041, prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3042(w_eco3042, prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3043(w_eco3043, prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3044(w_eco3044, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3045(w_eco3045, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3046(w_eco3046, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3047(w_eco3047, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3048(w_eco3048, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3049(w_eco3049, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3050(w_eco3050, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3051(w_eco3051, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3052(w_eco3052, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3053(w_eco3053, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3054(w_eco3054, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3055(w_eco3055, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3056(w_eco3056, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3057(w_eco3057, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3058(w_eco3058, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3059(w_eco3059, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3060(w_eco3060, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3061(w_eco3061, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3062(w_eco3062, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3063(w_eco3063, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3064(w_eco3064, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3065(w_eco3065, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3066(w_eco3066, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3067(w_eco3067, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3068(w_eco3068, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3069(w_eco3069, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3070(w_eco3070, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3071(w_eco3071, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3072(w_eco3072, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3073(w_eco3073, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3074(w_eco3074, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3075(w_eco3075, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3076(w_eco3076, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3077(w_eco3077, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3078(w_eco3078, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3079(w_eco3079, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3080(w_eco3080, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3081(w_eco3081, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3082(w_eco3082, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3083(w_eco3083, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3084(w_eco3084, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3085(w_eco3085, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3086(w_eco3086, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3087(w_eco3087, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3088(w_eco3088, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3089(w_eco3089, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3090(w_eco3090, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3091(w_eco3091, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3092(w_eco3092, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3093(w_eco3093, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3094(w_eco3094, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3095(w_eco3095, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3096(w_eco3096, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3097(w_eco3097, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3098(w_eco3098, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3099(w_eco3099, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[9], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3100(w_eco3100, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3101(w_eco3101, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3102(w_eco3102, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3103(w_eco3103, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3104(w_eco3104, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3105(w_eco3105, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3106(w_eco3106, !prev_cnt[14], prev_cnt[0], prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3107(w_eco3107, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3108(w_eco3108, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[8], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3109(w_eco3109, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3110(w_eco3110, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3111(w_eco3111, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3112(w_eco3112, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3113(w_eco3113, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3114(w_eco3114, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3115(w_eco3115, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3116(w_eco3116, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3117(w_eco3117, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3118(w_eco3118, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3119(w_eco3119, !Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3120(w_eco3120, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3121(w_eco3121, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3122(w_eco3122, !Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3123(w_eco3123, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3124(w_eco3124, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3125(w_eco3125, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3126(w_eco3126, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3127(w_eco3127, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3128(w_eco3128, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3129(w_eco3129, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3130(w_eco3130, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3131(w_eco3131, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3132(w_eco3132, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3133(w_eco3133, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3134(w_eco3134, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3135(w_eco3135, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3136(w_eco3136, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3137(w_eco3137, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3138(w_eco3138, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3139(w_eco3139, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3140(w_eco3140, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3141(w_eco3141, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3142(w_eco3142, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3143(w_eco3143, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3144(w_eco3144, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3145(w_eco3145, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3146(w_eco3146, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3147(w_eco3147, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3148(w_eco3148, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3149(w_eco3149, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3150(w_eco3150, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3151(w_eco3151, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3152(w_eco3152, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3153(w_eco3153, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3154(w_eco3154, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3155(w_eco3155, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3156(w_eco3156, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3157(w_eco3157, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3158(w_eco3158, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3159(w_eco3159, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3160(w_eco3160, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3161(w_eco3161, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3162(w_eco3162, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3163(w_eco3163, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3164(w_eco3164, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3165(w_eco3165, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3166(w_eco3166, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3167(w_eco3167, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3168(w_eco3168, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3169(w_eco3169, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3170(w_eco3170, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3171(w_eco3171, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3172(w_eco3172, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3173(w_eco3173, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3174(w_eco3174, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3175(w_eco3175, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3176(w_eco3176, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3177(w_eco3177, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3178(w_eco3178, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3179(w_eco3179, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3180(w_eco3180, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3181(w_eco3181, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3182(w_eco3182, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3183(w_eco3183, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3184(w_eco3184, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3185(w_eco3185, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3186(w_eco3186, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3187(w_eco3187, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3188(w_eco3188, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3189(w_eco3189, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3190(w_eco3190, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3191(w_eco3191, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3192(w_eco3192, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3193(w_eco3193, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3194(w_eco3194, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3195(w_eco3195, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3196(w_eco3196, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3197(w_eco3197, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3198(w_eco3198, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3199(w_eco3199, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3200(w_eco3200, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3201(w_eco3201, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3202(w_eco3202, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3203(w_eco3203, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3204(w_eco3204, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3205(w_eco3205, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3206(w_eco3206, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3207(w_eco3207, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3208(w_eco3208, prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3209(w_eco3209, prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3210(w_eco3210, prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3211(w_eco3211, prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3212(w_eco3212, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3213(w_eco3213, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3214(w_eco3214, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3215(w_eco3215, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3216(w_eco3216, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3217(w_eco3217, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3218(w_eco3218, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3219(w_eco3219, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3220(w_eco3220, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3221(w_eco3221, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3222(w_eco3222, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3223(w_eco3223, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3224(w_eco3224, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3225(w_eco3225, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3226(w_eco3226, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3227(w_eco3227, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3228(w_eco3228, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3229(w_eco3229, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3230(w_eco3230, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3231(w_eco3231, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3232(w_eco3232, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3233(w_eco3233, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3234(w_eco3234, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3235(w_eco3235, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3236(w_eco3236, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3237(w_eco3237, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3238(w_eco3238, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3239(w_eco3239, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3240(w_eco3240, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3241(w_eco3241, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3242(w_eco3242, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3243(w_eco3243, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3244(w_eco3244, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3245(w_eco3245, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3246(w_eco3246, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3247(w_eco3247, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3248(w_eco3248, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3249(w_eco3249, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3250(w_eco3250, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3251(w_eco3251, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3252(w_eco3252, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3253(w_eco3253, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3254(w_eco3254, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3255(w_eco3255, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3256(w_eco3256, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3257(w_eco3257, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3258(w_eco3258, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3259(w_eco3259, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3260(w_eco3260, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3261(w_eco3261, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3262(w_eco3262, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3263(w_eco3263, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3264(w_eco3264, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3265(w_eco3265, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3266(w_eco3266, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3267(w_eco3267, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3268(w_eco3268, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3269(w_eco3269, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3270(w_eco3270, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3271(w_eco3271, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3272(w_eco3272, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3273(w_eco3273, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3274(w_eco3274, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3275(w_eco3275, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3276(w_eco3276, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3277(w_eco3277, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3278(w_eco3278, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3279(w_eco3279, !prev_cnt[14], prev_cnt[3], prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3280(w_eco3280, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[12], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3281(w_eco3281, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3282(w_eco3282, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3283(w_eco3283, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_3284(w_eco3284, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3285(w_eco3285, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3286(w_eco3286, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3287(w_eco3287, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3288(w_eco3288, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3289(w_eco3289, !Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3290(w_eco3290, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3291(w_eco3291, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3292(w_eco3292, !Tgate[5], !Tgdel[5], !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3293(w_eco3293, !Tgate[5], !Tgdel[5], !Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3294(w_eco3294, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3295(w_eco3295, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3296(w_eco3296, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3297(w_eco3297, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3298(w_eco3298, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3299(w_eco3299, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3300(w_eco3300, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3301(w_eco3301, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3302(w_eco3302, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3303(w_eco3303, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3304(w_eco3304, prev_cnt[1], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3305(w_eco3305, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3306(w_eco3306, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3307(w_eco3307, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3308(w_eco3308, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3309(w_eco3309, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3310(w_eco3310, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3311(w_eco3311, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3312(w_eco3312, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3313(w_eco3313, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3314(w_eco3314, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3315(w_eco3315, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3316(w_eco3316, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3317(w_eco3317, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3318(w_eco3318, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3319(w_eco3319, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3320(w_eco3320, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3321(w_eco3321, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3322(w_eco3322, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3323(w_eco3323, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3324(w_eco3324, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3325(w_eco3325, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3326(w_eco3326, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3327(w_eco3327, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3328(w_eco3328, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3329(w_eco3329, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3330(w_eco3330, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3331(w_eco3331, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3332(w_eco3332, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3333(w_eco3333, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3334(w_eco3334, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3335(w_eco3335, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3336(w_eco3336, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3337(w_eco3337, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3338(w_eco3338, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3339(w_eco3339, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3340(w_eco3340, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3341(w_eco3341, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3342(w_eco3342, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3343(w_eco3343, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3344(w_eco3344, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3345(w_eco3345, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3346(w_eco3346, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3347(w_eco3347, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3348(w_eco3348, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3349(w_eco3349, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3350(w_eco3350, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3351(w_eco3351, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3352(w_eco3352, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3353(w_eco3353, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3354(w_eco3354, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3355(w_eco3355, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3356(w_eco3356, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3357(w_eco3357, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3358(w_eco3358, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3359(w_eco3359, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3360(w_eco3360, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3361(w_eco3361, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3362(w_eco3362, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3363(w_eco3363, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3364(w_eco3364, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3365(w_eco3365, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3366(w_eco3366, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3367(w_eco3367, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3368(w_eco3368, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3369(w_eco3369, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3370(w_eco3370, prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3371(w_eco3371, prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3372(w_eco3372, prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3373(w_eco3373, prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3374(w_eco3374, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3375(w_eco3375, prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3376(w_eco3376, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3377(w_eco3377, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3378(w_eco3378, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3379(w_eco3379, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3380(w_eco3380, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3381(w_eco3381, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3382(w_eco3382, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3383(w_eco3383, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3384(w_eco3384, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3385(w_eco3385, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3386(w_eco3386, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3387(w_eco3387, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3388(w_eco3388, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3389(w_eco3389, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3390(w_eco3390, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3391(w_eco3391, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3392(w_eco3392, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3393(w_eco3393, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3394(w_eco3394, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3395(w_eco3395, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3396(w_eco3396, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3397(w_eco3397, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3398(w_eco3398, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3399(w_eco3399, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3400(w_eco3400, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3401(w_eco3401, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3402(w_eco3402, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3403(w_eco3403, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3404(w_eco3404, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3405(w_eco3405, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3406(w_eco3406, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3407(w_eco3407, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3408(w_eco3408, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3409(w_eco3409, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3410(w_eco3410, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3411(w_eco3411, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3412(w_eco3412, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3413(w_eco3413, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3414(w_eco3414, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3415(w_eco3415, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3416(w_eco3416, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3417(w_eco3417, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3418(w_eco3418, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3419(w_eco3419, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3420(w_eco3420, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3421(w_eco3421, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3422(w_eco3422, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3423(w_eco3423, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3424(w_eco3424, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3425(w_eco3425, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3426(w_eco3426, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3427(w_eco3427, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3428(w_eco3428, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3429(w_eco3429, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3430(w_eco3430, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3431(w_eco3431, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3432(w_eco3432, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3433(w_eco3433, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3434(w_eco3434, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3435(w_eco3435, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3436(w_eco3436, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3437(w_eco3437, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3438(w_eco3438, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3439(w_eco3439, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3440(w_eco3440, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3441(w_eco3441, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3442(w_eco3442, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3443(w_eco3443, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3444(w_eco3444, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3445(w_eco3445, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3446(w_eco3446, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3447(w_eco3447, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], prev_cnt[13], !rst, prev_state[1], !prev_state[0]);
	and _ECO_3448(w_eco3448, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3449(w_eco3449, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_3450(w_eco3450, !Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3451(w_eco3451, !Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3452(w_eco3452, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3453(w_eco3453, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3454(w_eco3454, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3455(w_eco3455, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3456(w_eco3456, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3457(w_eco3457, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3458(w_eco3458, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3459(w_eco3459, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3460(w_eco3460, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3461(w_eco3461, prev_cnt[2], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3462(w_eco3462, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3463(w_eco3463, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3464(w_eco3464, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3465(w_eco3465, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3466(w_eco3466, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3467(w_eco3467, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3468(w_eco3468, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3469(w_eco3469, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3470(w_eco3470, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3471(w_eco3471, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3472(w_eco3472, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3473(w_eco3473, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3474(w_eco3474, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3475(w_eco3475, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3476(w_eco3476, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3477(w_eco3477, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3478(w_eco3478, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3479(w_eco3479, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3480(w_eco3480, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3481(w_eco3481, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3482(w_eco3482, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3483(w_eco3483, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3484(w_eco3484, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3485(w_eco3485, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3486(w_eco3486, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3487(w_eco3487, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3488(w_eco3488, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3489(w_eco3489, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3490(w_eco3490, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3491(w_eco3491, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3492(w_eco3492, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3493(w_eco3493, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3494(w_eco3494, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3495(w_eco3495, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3496(w_eco3496, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3497(w_eco3497, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3498(w_eco3498, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3499(w_eco3499, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3500(w_eco3500, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3501(w_eco3501, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3502(w_eco3502, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3503(w_eco3503, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3504(w_eco3504, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3505(w_eco3505, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3506(w_eco3506, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3507(w_eco3507, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3508(w_eco3508, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3509(w_eco3509, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3510(w_eco3510, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3511(w_eco3511, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3512(w_eco3512, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3513(w_eco3513, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3514(w_eco3514, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3515(w_eco3515, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3516(w_eco3516, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3517(w_eco3517, prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3518(w_eco3518, prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3519(w_eco3519, prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3520(w_eco3520, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3521(w_eco3521, prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3522(w_eco3522, !Tgate[5], !Tgdel[5], prev_cnt[1], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3523(w_eco3523, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3524(w_eco3524, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3525(w_eco3525, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3526(w_eco3526, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3527(w_eco3527, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3528(w_eco3528, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3529(w_eco3529, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3530(w_eco3530, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3531(w_eco3531, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3532(w_eco3532, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3533(w_eco3533, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3534(w_eco3534, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3535(w_eco3535, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3536(w_eco3536, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3537(w_eco3537, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3538(w_eco3538, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3539(w_eco3539, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3540(w_eco3540, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3541(w_eco3541, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3542(w_eco3542, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3543(w_eco3543, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3544(w_eco3544, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3545(w_eco3545, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3546(w_eco3546, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3547(w_eco3547, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3548(w_eco3548, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3549(w_eco3549, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3550(w_eco3550, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3551(w_eco3551, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3552(w_eco3552, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3553(w_eco3553, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3554(w_eco3554, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3555(w_eco3555, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3556(w_eco3556, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3557(w_eco3557, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3558(w_eco3558, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3559(w_eco3559, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3560(w_eco3560, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3561(w_eco3561, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3562(w_eco3562, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3563(w_eco3563, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3564(w_eco3564, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3565(w_eco3565, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3566(w_eco3566, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3567(w_eco3567, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3568(w_eco3568, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3569(w_eco3569, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3570(w_eco3570, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3571(w_eco3571, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3572(w_eco3572, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3573(w_eco3573, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3574(w_eco3574, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3575(w_eco3575, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3576(w_eco3576, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3577(w_eco3577, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3578(w_eco3578, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3579(w_eco3579, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3580(w_eco3580, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3581(w_eco3581, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3582(w_eco3582, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3583(w_eco3583, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3584(w_eco3584, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3585(w_eco3585, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3586(w_eco3586, Tsync[5], prev_cnt[1], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3587(w_eco3587, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3588(w_eco3588, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3589(w_eco3589, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3590(w_eco3590, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3591(w_eco3591, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[15], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3592(w_eco3592, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3593(w_eco3593, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3594(w_eco3594, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3595(w_eco3595, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3596(w_eco3596, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3597(w_eco3597, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3598(w_eco3598, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3599(w_eco3599, prev_cnt[4], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3600(w_eco3600, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3601(w_eco3601, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3602(w_eco3602, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3603(w_eco3603, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3604(w_eco3604, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3605(w_eco3605, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3606(w_eco3606, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3607(w_eco3607, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3608(w_eco3608, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3609(w_eco3609, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3610(w_eco3610, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3611(w_eco3611, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3612(w_eco3612, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3613(w_eco3613, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3614(w_eco3614, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3615(w_eco3615, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3616(w_eco3616, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3617(w_eco3617, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3618(w_eco3618, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3619(w_eco3619, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3620(w_eco3620, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3621(w_eco3621, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3622(w_eco3622, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3623(w_eco3623, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3624(w_eco3624, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3625(w_eco3625, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3626(w_eco3626, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3627(w_eco3627, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3628(w_eco3628, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3629(w_eco3629, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3630(w_eco3630, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3631(w_eco3631, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3632(w_eco3632, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3633(w_eco3633, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3634(w_eco3634, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3635(w_eco3635, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3636(w_eco3636, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3637(w_eco3637, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3638(w_eco3638, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3639(w_eco3639, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3640(w_eco3640, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3641(w_eco3641, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3642(w_eco3642, !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3643(w_eco3643, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3644(w_eco3644, prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3645(w_eco3645, prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3646(w_eco3646, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3647(w_eco3647, prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3648(w_eco3648, !Tgate[5], !Tgdel[5], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3649(w_eco3649, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3650(w_eco3650, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3651(w_eco3651, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3652(w_eco3652, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3653(w_eco3653, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3654(w_eco3654, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3655(w_eco3655, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3656(w_eco3656, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3657(w_eco3657, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3658(w_eco3658, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3659(w_eco3659, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3660(w_eco3660, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3661(w_eco3661, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3662(w_eco3662, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3663(w_eco3663, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3664(w_eco3664, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3665(w_eco3665, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3666(w_eco3666, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3667(w_eco3667, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3668(w_eco3668, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3669(w_eco3669, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3670(w_eco3670, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3671(w_eco3671, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3672(w_eco3672, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3673(w_eco3673, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3674(w_eco3674, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3675(w_eco3675, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3676(w_eco3676, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3677(w_eco3677, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3678(w_eco3678, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3679(w_eco3679, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3680(w_eco3680, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3681(w_eco3681, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3682(w_eco3682, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3683(w_eco3683, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3684(w_eco3684, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3685(w_eco3685, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3686(w_eco3686, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3687(w_eco3687, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3688(w_eco3688, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3689(w_eco3689, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3690(w_eco3690, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3691(w_eco3691, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3692(w_eco3692, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3693(w_eco3693, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3694(w_eco3694, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3695(w_eco3695, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3696(w_eco3696, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3697(w_eco3697, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3698(w_eco3698, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3699(w_eco3699, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3700(w_eco3700, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3701(w_eco3701, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3702(w_eco3702, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3703(w_eco3703, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3704(w_eco3704, Tsync[5], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3705(w_eco3705, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3706(w_eco3706, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3707(w_eco3707, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3708(w_eco3708, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[11], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3709(w_eco3709, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[1], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3710(w_eco3710, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3711(w_eco3711, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3712(w_eco3712, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3713(w_eco3713, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3714(w_eco3714, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3715(w_eco3715, prev_cnt[0], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3716(w_eco3716, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3717(w_eco3717, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3718(w_eco3718, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3719(w_eco3719, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3720(w_eco3720, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3721(w_eco3721, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3722(w_eco3722, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3723(w_eco3723, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3724(w_eco3724, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3725(w_eco3725, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3726(w_eco3726, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3727(w_eco3727, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3728(w_eco3728, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3729(w_eco3729, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3730(w_eco3730, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3731(w_eco3731, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3732(w_eco3732, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3733(w_eco3733, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3734(w_eco3734, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3735(w_eco3735, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3736(w_eco3736, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3737(w_eco3737, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3738(w_eco3738, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3739(w_eco3739, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3740(w_eco3740, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3741(w_eco3741, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3742(w_eco3742, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3743(w_eco3743, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3744(w_eco3744, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3745(w_eco3745, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3746(w_eco3746, !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3747(w_eco3747, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3748(w_eco3748, prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3749(w_eco3749, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3750(w_eco3750, prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3751(w_eco3751, !Tgate[5], !Tgdel[5], prev_cnt[4], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3752(w_eco3752, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3753(w_eco3753, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3754(w_eco3754, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3755(w_eco3755, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3756(w_eco3756, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3757(w_eco3757, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3758(w_eco3758, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3759(w_eco3759, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3760(w_eco3760, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3761(w_eco3761, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3762(w_eco3762, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3763(w_eco3763, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3764(w_eco3764, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3765(w_eco3765, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3766(w_eco3766, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3767(w_eco3767, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3768(w_eco3768, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3769(w_eco3769, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3770(w_eco3770, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3771(w_eco3771, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3772(w_eco3772, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3773(w_eco3773, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3774(w_eco3774, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3775(w_eco3775, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3776(w_eco3776, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3777(w_eco3777, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3778(w_eco3778, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3779(w_eco3779, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3780(w_eco3780, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3781(w_eco3781, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3782(w_eco3782, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3783(w_eco3783, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3784(w_eco3784, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3785(w_eco3785, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3786(w_eco3786, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3787(w_eco3787, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3788(w_eco3788, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3789(w_eco3789, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3790(w_eco3790, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3791(w_eco3791, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3792(w_eco3792, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3793(w_eco3793, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3794(w_eco3794, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3795(w_eco3795, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3796(w_eco3796, Tsync[5], prev_cnt[4], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3797(w_eco3797, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3798(w_eco3798, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3799(w_eco3799, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[6], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3800(w_eco3800, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[2], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3801(w_eco3801, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3802(w_eco3802, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3803(w_eco3803, prev_cnt[3], prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3804(w_eco3804, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3805(w_eco3805, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3806(w_eco3806, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3807(w_eco3807, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3808(w_eco3808, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3809(w_eco3809, !Tgate[5], !Tgdel[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3810(w_eco3810, !Tgate[5], !Tgdel[5], prev_cnt[3], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3811(w_eco3811, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3812(w_eco3812, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3813(w_eco3813, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3814(w_eco3814, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3815(w_eco3815, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3816(w_eco3816, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3817(w_eco3817, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3818(w_eco3818, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3819(w_eco3819, !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3820(w_eco3820, !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3821(w_eco3821, !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3822(w_eco3822, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3823(w_eco3823, prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3824(w_eco3824, !Tgate[5], !Tgdel[5], prev_cnt[0], !prev_cnt[5], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3825(w_eco3825, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3826(w_eco3826, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3827(w_eco3827, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3828(w_eco3828, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3829(w_eco3829, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3830(w_eco3830, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3831(w_eco3831, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3832(w_eco3832, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3833(w_eco3833, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3834(w_eco3834, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3835(w_eco3835, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3836(w_eco3836, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3837(w_eco3837, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3838(w_eco3838, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3839(w_eco3839, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3840(w_eco3840, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3841(w_eco3841, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3842(w_eco3842, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3843(w_eco3843, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3844(w_eco3844, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3845(w_eco3845, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3846(w_eco3846, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3847(w_eco3847, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3848(w_eco3848, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3849(w_eco3849, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3850(w_eco3850, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3851(w_eco3851, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3852(w_eco3852, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3853(w_eco3853, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3854(w_eco3854, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3855(w_eco3855, Tsync[5], !prev_cnt[14], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3856(w_eco3856, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3857(w_eco3857, Tsync[5], prev_cnt[0], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3858(w_eco3858, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3859(w_eco3859, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[10], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3860(w_eco3860, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[4], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3861(w_eco3861, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3862(w_eco3862, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !rst, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3863(w_eco3863, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3864(w_eco3864, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3865(w_eco3865, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3866(w_eco3866, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3867(w_eco3867, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3868(w_eco3868, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3869(w_eco3869, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3870(w_eco3870, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3871(w_eco3871, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3872(w_eco3872, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3873(w_eco3873, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3874(w_eco3874, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3875(w_eco3875, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3876(w_eco3876, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3877(w_eco3877, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3878(w_eco3878, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_3879(w_eco3879, Tsync[5], !prev_cnt[14], prev_cnt[4], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3880(w_eco3880, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3881(w_eco3881, Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3882(w_eco3882, Tsync[5], prev_cnt[3], !prev_cnt[5], prev_cnt[8], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3883(w_eco3883, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[0], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3884(w_eco3884, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3885(w_eco3885, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3886(w_eco3886, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3887(w_eco3887, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3888(w_eco3888, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3889(w_eco3889, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3890(w_eco3890, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3891(w_eco3891, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3892(w_eco3892, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3893(w_eco3893, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[12], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3894(w_eco3894, !Tgate[5], !Tgdel[5], Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3895(w_eco3895, !Tgate[5], !Tgdel[5], Tsync[5], prev_cnt[3], !prev_cnt[5], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3896(w_eco3896, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3897(w_eco3897, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3898(w_eco3898, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_3899(w_eco3899, Tsync[5], !prev_cnt[14], prev_cnt[3], !prev_cnt[5], prev_cnt[13], ena, !rst, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_3900(w_eco3900, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914, w_eco1915, w_eco1916, w_eco1917, w_eco1918, w_eco1919, w_eco1920, w_eco1921, w_eco1922, w_eco1923, w_eco1924, w_eco1925, w_eco1926, w_eco1927, w_eco1928, w_eco1929, w_eco1930, w_eco1931, w_eco1932, w_eco1933, w_eco1934, w_eco1935, w_eco1936, w_eco1937, w_eco1938, w_eco1939, w_eco1940, w_eco1941, w_eco1942, w_eco1943, w_eco1944, w_eco1945, w_eco1946, w_eco1947, w_eco1948, w_eco1949, w_eco1950, w_eco1951, w_eco1952, w_eco1953, w_eco1954, w_eco1955, w_eco1956, w_eco1957, w_eco1958, w_eco1959, w_eco1960, w_eco1961, w_eco1962, w_eco1963, w_eco1964, w_eco1965, w_eco1966, w_eco1967, w_eco1968, w_eco1969, w_eco1970, w_eco1971, w_eco1972, w_eco1973, w_eco1974, w_eco1975, w_eco1976, w_eco1977, w_eco1978, w_eco1979, w_eco1980, w_eco1981, w_eco1982, w_eco1983, w_eco1984, w_eco1985, w_eco1986, w_eco1987, w_eco1988, w_eco1989, w_eco1990, w_eco1991, w_eco1992, w_eco1993, w_eco1994, w_eco1995, w_eco1996, w_eco1997, w_eco1998, w_eco1999, w_eco2000, w_eco2001, w_eco2002, w_eco2003, w_eco2004, w_eco2005, w_eco2006, w_eco2007, w_eco2008, w_eco2009, w_eco2010, w_eco2011, w_eco2012, w_eco2013, w_eco2014, w_eco2015, w_eco2016, w_eco2017, w_eco2018, w_eco2019, w_eco2020, w_eco2021, w_eco2022, w_eco2023, w_eco2024, w_eco2025, w_eco2026, w_eco2027, w_eco2028, w_eco2029, w_eco2030, w_eco2031, w_eco2032, w_eco2033, w_eco2034, w_eco2035, w_eco2036, w_eco2037, w_eco2038, w_eco2039, w_eco2040, w_eco2041, w_eco2042, w_eco2043, w_eco2044, w_eco2045, w_eco2046, w_eco2047, w_eco2048, w_eco2049, w_eco2050, w_eco2051, w_eco2052, w_eco2053, w_eco2054, w_eco2055, w_eco2056, w_eco2057, w_eco2058, w_eco2059, w_eco2060, w_eco2061, w_eco2062, w_eco2063, w_eco2064, w_eco2065, w_eco2066, w_eco2067, w_eco2068, w_eco2069, w_eco2070, w_eco2071, w_eco2072, w_eco2073, w_eco2074, w_eco2075, w_eco2076, w_eco2077, w_eco2078, w_eco2079, w_eco2080, w_eco2081, w_eco2082, w_eco2083, w_eco2084, w_eco2085, w_eco2086, w_eco2087, w_eco2088, w_eco2089, w_eco2090, w_eco2091, w_eco2092, w_eco2093, w_eco2094, w_eco2095, w_eco2096, w_eco2097, w_eco2098, w_eco2099, w_eco2100, w_eco2101, w_eco2102, w_eco2103, w_eco2104, w_eco2105, w_eco2106, w_eco2107, w_eco2108, w_eco2109, w_eco2110, w_eco2111, w_eco2112, w_eco2113, w_eco2114, w_eco2115, w_eco2116, w_eco2117, w_eco2118, w_eco2119, w_eco2120, w_eco2121, w_eco2122, w_eco2123, w_eco2124, w_eco2125, w_eco2126, w_eco2127, w_eco2128, w_eco2129, w_eco2130, w_eco2131, w_eco2132, w_eco2133, w_eco2134, w_eco2135, w_eco2136, w_eco2137, w_eco2138, w_eco2139, w_eco2140, w_eco2141, w_eco2142, w_eco2143, w_eco2144, w_eco2145, w_eco2146, w_eco2147, w_eco2148, w_eco2149, w_eco2150, w_eco2151, w_eco2152, w_eco2153, w_eco2154, w_eco2155, w_eco2156, w_eco2157, w_eco2158, w_eco2159, w_eco2160, w_eco2161, w_eco2162, w_eco2163, w_eco2164, w_eco2165, w_eco2166, w_eco2167, w_eco2168, w_eco2169, w_eco2170, w_eco2171, w_eco2172, w_eco2173, w_eco2174, w_eco2175, w_eco2176, w_eco2177, w_eco2178, w_eco2179, w_eco2180, w_eco2181, w_eco2182, w_eco2183, w_eco2184, w_eco2185, w_eco2186, w_eco2187, w_eco2188, w_eco2189, w_eco2190, w_eco2191, w_eco2192, w_eco2193, w_eco2194, w_eco2195, w_eco2196, w_eco2197, w_eco2198, w_eco2199, w_eco2200, w_eco2201, w_eco2202, w_eco2203, w_eco2204, w_eco2205, w_eco2206, w_eco2207, w_eco2208, w_eco2209, w_eco2210, w_eco2211, w_eco2212, w_eco2213, w_eco2214, w_eco2215, w_eco2216, w_eco2217, w_eco2218, w_eco2219, w_eco2220, w_eco2221, w_eco2222, w_eco2223, w_eco2224, w_eco2225, w_eco2226, w_eco2227, w_eco2228, w_eco2229, w_eco2230, w_eco2231, w_eco2232, w_eco2233, w_eco2234, w_eco2235, w_eco2236, w_eco2237, w_eco2238, w_eco2239, w_eco2240, w_eco2241, w_eco2242, w_eco2243, w_eco2244, w_eco2245, w_eco2246, w_eco2247, w_eco2248, w_eco2249, w_eco2250, w_eco2251, w_eco2252, w_eco2253, w_eco2254, w_eco2255, w_eco2256, w_eco2257, w_eco2258, w_eco2259, w_eco2260, w_eco2261, w_eco2262, w_eco2263, w_eco2264, w_eco2265, w_eco2266, w_eco2267, w_eco2268, w_eco2269, w_eco2270, w_eco2271, w_eco2272, w_eco2273, w_eco2274, w_eco2275, w_eco2276, w_eco2277, w_eco2278, w_eco2279, w_eco2280, w_eco2281, w_eco2282, w_eco2283, w_eco2284, w_eco2285, w_eco2286, w_eco2287, w_eco2288, w_eco2289, w_eco2290, w_eco2291, w_eco2292, w_eco2293, w_eco2294, w_eco2295, w_eco2296, w_eco2297, w_eco2298, w_eco2299, w_eco2300, w_eco2301, w_eco2302, w_eco2303, w_eco2304, w_eco2305, w_eco2306, w_eco2307, w_eco2308, w_eco2309, w_eco2310, w_eco2311, w_eco2312, w_eco2313, w_eco2314, w_eco2315, w_eco2316, w_eco2317, w_eco2318, w_eco2319, w_eco2320, w_eco2321, w_eco2322, w_eco2323, w_eco2324, w_eco2325, w_eco2326, w_eco2327, w_eco2328, w_eco2329, w_eco2330, w_eco2331, w_eco2332, w_eco2333, w_eco2334, w_eco2335, w_eco2336, w_eco2337, w_eco2338, w_eco2339, w_eco2340, w_eco2341, w_eco2342, w_eco2343, w_eco2344, w_eco2345, w_eco2346, w_eco2347, w_eco2348, w_eco2349, w_eco2350, w_eco2351, w_eco2352, w_eco2353, w_eco2354, w_eco2355, w_eco2356, w_eco2357, w_eco2358, w_eco2359, w_eco2360, w_eco2361, w_eco2362, w_eco2363, w_eco2364, w_eco2365, w_eco2366, w_eco2367, w_eco2368, w_eco2369, w_eco2370, w_eco2371, w_eco2372, w_eco2373, w_eco2374, w_eco2375, w_eco2376, w_eco2377, w_eco2378, w_eco2379, w_eco2380, w_eco2381, w_eco2382, w_eco2383, w_eco2384, w_eco2385, w_eco2386, w_eco2387, w_eco2388, w_eco2389, w_eco2390, w_eco2391, w_eco2392, w_eco2393, w_eco2394, w_eco2395, w_eco2396, w_eco2397, w_eco2398, w_eco2399, w_eco2400, w_eco2401, w_eco2402, w_eco2403, w_eco2404, w_eco2405, w_eco2406, w_eco2407, w_eco2408, w_eco2409, w_eco2410, w_eco2411, w_eco2412, w_eco2413, w_eco2414, w_eco2415, w_eco2416, w_eco2417, w_eco2418, w_eco2419, w_eco2420, w_eco2421, w_eco2422, w_eco2423, w_eco2424, w_eco2425, w_eco2426, w_eco2427, w_eco2428, w_eco2429, w_eco2430, w_eco2431, w_eco2432, w_eco2433, w_eco2434, w_eco2435, w_eco2436, w_eco2437, w_eco2438, w_eco2439, w_eco2440, w_eco2441, w_eco2442, w_eco2443, w_eco2444, w_eco2445, w_eco2446, w_eco2447, w_eco2448, w_eco2449, w_eco2450, w_eco2451, w_eco2452, w_eco2453, w_eco2454, w_eco2455, w_eco2456, w_eco2457, w_eco2458, w_eco2459, w_eco2460, w_eco2461, w_eco2462, w_eco2463, w_eco2464, w_eco2465, w_eco2466, w_eco2467, w_eco2468, w_eco2469, w_eco2470, w_eco2471, w_eco2472, w_eco2473, w_eco2474, w_eco2475, w_eco2476, w_eco2477, w_eco2478, w_eco2479, w_eco2480, w_eco2481, w_eco2482, w_eco2483, w_eco2484, w_eco2485, w_eco2486, w_eco2487, w_eco2488, w_eco2489, w_eco2490, w_eco2491, w_eco2492, w_eco2493, w_eco2494, w_eco2495, w_eco2496, w_eco2497, w_eco2498, w_eco2499, w_eco2500, w_eco2501, w_eco2502, w_eco2503, w_eco2504, w_eco2505, w_eco2506, w_eco2507, w_eco2508, w_eco2509, w_eco2510, w_eco2511, w_eco2512, w_eco2513, w_eco2514, w_eco2515, w_eco2516, w_eco2517, w_eco2518, w_eco2519, w_eco2520, w_eco2521, w_eco2522, w_eco2523, w_eco2524, w_eco2525, w_eco2526, w_eco2527, w_eco2528, w_eco2529, w_eco2530, w_eco2531, w_eco2532, w_eco2533, w_eco2534, w_eco2535, w_eco2536, w_eco2537, w_eco2538, w_eco2539, w_eco2540, w_eco2541, w_eco2542, w_eco2543, w_eco2544, w_eco2545, w_eco2546, w_eco2547, w_eco2548, w_eco2549, w_eco2550, w_eco2551, w_eco2552, w_eco2553, w_eco2554, w_eco2555, w_eco2556, w_eco2557, w_eco2558, w_eco2559, w_eco2560, w_eco2561, w_eco2562, w_eco2563, w_eco2564, w_eco2565, w_eco2566, w_eco2567, w_eco2568, w_eco2569, w_eco2570, w_eco2571, w_eco2572, w_eco2573, w_eco2574, w_eco2575, w_eco2576, w_eco2577, w_eco2578, w_eco2579, w_eco2580, w_eco2581, w_eco2582, w_eco2583, w_eco2584, w_eco2585, w_eco2586, w_eco2587, w_eco2588, w_eco2589, w_eco2590, w_eco2591, w_eco2592, w_eco2593, w_eco2594, w_eco2595, w_eco2596, w_eco2597, w_eco2598, w_eco2599, w_eco2600, w_eco2601, w_eco2602, w_eco2603, w_eco2604, w_eco2605, w_eco2606, w_eco2607, w_eco2608, w_eco2609, w_eco2610, w_eco2611, w_eco2612, w_eco2613, w_eco2614, w_eco2615, w_eco2616, w_eco2617, w_eco2618, w_eco2619, w_eco2620, w_eco2621, w_eco2622, w_eco2623, w_eco2624, w_eco2625, w_eco2626, w_eco2627, w_eco2628, w_eco2629, w_eco2630, w_eco2631, w_eco2632, w_eco2633, w_eco2634, w_eco2635, w_eco2636, w_eco2637, w_eco2638, w_eco2639, w_eco2640, w_eco2641, w_eco2642, w_eco2643, w_eco2644, w_eco2645, w_eco2646, w_eco2647, w_eco2648, w_eco2649, w_eco2650, w_eco2651, w_eco2652, w_eco2653, w_eco2654, w_eco2655, w_eco2656, w_eco2657, w_eco2658, w_eco2659, w_eco2660, w_eco2661, w_eco2662, w_eco2663, w_eco2664, w_eco2665, w_eco2666, w_eco2667, w_eco2668, w_eco2669, w_eco2670, w_eco2671, w_eco2672, w_eco2673, w_eco2674, w_eco2675, w_eco2676, w_eco2677, w_eco2678, w_eco2679, w_eco2680, w_eco2681, w_eco2682, w_eco2683, w_eco2684, w_eco2685, w_eco2686, w_eco2687, w_eco2688, w_eco2689, w_eco2690, w_eco2691, w_eco2692, w_eco2693, w_eco2694, w_eco2695, w_eco2696, w_eco2697, w_eco2698, w_eco2699, w_eco2700, w_eco2701, w_eco2702, w_eco2703, w_eco2704, w_eco2705, w_eco2706, w_eco2707, w_eco2708, w_eco2709, w_eco2710, w_eco2711, w_eco2712, w_eco2713, w_eco2714, w_eco2715, w_eco2716, w_eco2717, w_eco2718, w_eco2719, w_eco2720, w_eco2721, w_eco2722, w_eco2723, w_eco2724, w_eco2725, w_eco2726, w_eco2727, w_eco2728, w_eco2729, w_eco2730, w_eco2731, w_eco2732, w_eco2733, w_eco2734, w_eco2735, w_eco2736, w_eco2737, w_eco2738, w_eco2739, w_eco2740, w_eco2741, w_eco2742, w_eco2743, w_eco2744, w_eco2745, w_eco2746, w_eco2747, w_eco2748, w_eco2749, w_eco2750, w_eco2751, w_eco2752, w_eco2753, w_eco2754, w_eco2755, w_eco2756, w_eco2757, w_eco2758, w_eco2759, w_eco2760, w_eco2761, w_eco2762, w_eco2763, w_eco2764, w_eco2765, w_eco2766, w_eco2767, w_eco2768, w_eco2769, w_eco2770, w_eco2771, w_eco2772, w_eco2773, w_eco2774, w_eco2775, w_eco2776, w_eco2777, w_eco2778, w_eco2779, w_eco2780, w_eco2781, w_eco2782, w_eco2783, w_eco2784, w_eco2785, w_eco2786, w_eco2787, w_eco2788, w_eco2789, w_eco2790, w_eco2791, w_eco2792, w_eco2793, w_eco2794, w_eco2795, w_eco2796, w_eco2797, w_eco2798, w_eco2799, w_eco2800, w_eco2801, w_eco2802, w_eco2803, w_eco2804, w_eco2805, w_eco2806, w_eco2807, w_eco2808, w_eco2809, w_eco2810, w_eco2811, w_eco2812, w_eco2813, w_eco2814, w_eco2815, w_eco2816, w_eco2817, w_eco2818, w_eco2819, w_eco2820, w_eco2821, w_eco2822, w_eco2823, w_eco2824, w_eco2825, w_eco2826, w_eco2827, w_eco2828, w_eco2829, w_eco2830, w_eco2831, w_eco2832, w_eco2833, w_eco2834, w_eco2835, w_eco2836, w_eco2837, w_eco2838, w_eco2839, w_eco2840, w_eco2841, w_eco2842, w_eco2843, w_eco2844, w_eco2845, w_eco2846, w_eco2847, w_eco2848, w_eco2849, w_eco2850, w_eco2851, w_eco2852, w_eco2853, w_eco2854, w_eco2855, w_eco2856, w_eco2857, w_eco2858, w_eco2859, w_eco2860, w_eco2861, w_eco2862, w_eco2863, w_eco2864, w_eco2865, w_eco2866, w_eco2867, w_eco2868, w_eco2869, w_eco2870, w_eco2871, w_eco2872, w_eco2873, w_eco2874, w_eco2875, w_eco2876, w_eco2877, w_eco2878, w_eco2879, w_eco2880, w_eco2881, w_eco2882, w_eco2883, w_eco2884, w_eco2885, w_eco2886, w_eco2887, w_eco2888, w_eco2889, w_eco2890, w_eco2891, w_eco2892, w_eco2893, w_eco2894, w_eco2895, w_eco2896, w_eco2897, w_eco2898, w_eco2899, w_eco2900, w_eco2901, w_eco2902, w_eco2903, w_eco2904, w_eco2905, w_eco2906, w_eco2907, w_eco2908, w_eco2909, w_eco2910, w_eco2911, w_eco2912, w_eco2913, w_eco2914, w_eco2915, w_eco2916, w_eco2917, w_eco2918, w_eco2919, w_eco2920, w_eco2921, w_eco2922, w_eco2923, w_eco2924, w_eco2925, w_eco2926, w_eco2927, w_eco2928, w_eco2929, w_eco2930, w_eco2931, w_eco2932, w_eco2933, w_eco2934, w_eco2935, w_eco2936, w_eco2937, w_eco2938, w_eco2939, w_eco2940, w_eco2941, w_eco2942, w_eco2943, w_eco2944, w_eco2945, w_eco2946, w_eco2947, w_eco2948, w_eco2949, w_eco2950, w_eco2951, w_eco2952, w_eco2953, w_eco2954, w_eco2955, w_eco2956, w_eco2957, w_eco2958, w_eco2959, w_eco2960, w_eco2961, w_eco2962, w_eco2963, w_eco2964, w_eco2965, w_eco2966, w_eco2967, w_eco2968, w_eco2969, w_eco2970, w_eco2971, w_eco2972, w_eco2973, w_eco2974, w_eco2975, w_eco2976, w_eco2977, w_eco2978, w_eco2979, w_eco2980, w_eco2981, w_eco2982, w_eco2983, w_eco2984, w_eco2985, w_eco2986, w_eco2987, w_eco2988, w_eco2989, w_eco2990, w_eco2991, w_eco2992, w_eco2993, w_eco2994, w_eco2995, w_eco2996, w_eco2997, w_eco2998, w_eco2999, w_eco3000, w_eco3001, w_eco3002, w_eco3003, w_eco3004, w_eco3005, w_eco3006, w_eco3007, w_eco3008, w_eco3009, w_eco3010, w_eco3011, w_eco3012, w_eco3013, w_eco3014, w_eco3015, w_eco3016, w_eco3017, w_eco3018, w_eco3019, w_eco3020, w_eco3021, w_eco3022, w_eco3023, w_eco3024, w_eco3025, w_eco3026, w_eco3027, w_eco3028, w_eco3029, w_eco3030, w_eco3031, w_eco3032, w_eco3033, w_eco3034, w_eco3035, w_eco3036, w_eco3037, w_eco3038, w_eco3039, w_eco3040, w_eco3041, w_eco3042, w_eco3043, w_eco3044, w_eco3045, w_eco3046, w_eco3047, w_eco3048, w_eco3049, w_eco3050, w_eco3051, w_eco3052, w_eco3053, w_eco3054, w_eco3055, w_eco3056, w_eco3057, w_eco3058, w_eco3059, w_eco3060, w_eco3061, w_eco3062, w_eco3063, w_eco3064, w_eco3065, w_eco3066, w_eco3067, w_eco3068, w_eco3069, w_eco3070, w_eco3071, w_eco3072, w_eco3073, w_eco3074, w_eco3075, w_eco3076, w_eco3077, w_eco3078, w_eco3079, w_eco3080, w_eco3081, w_eco3082, w_eco3083, w_eco3084, w_eco3085, w_eco3086, w_eco3087, w_eco3088, w_eco3089, w_eco3090, w_eco3091, w_eco3092, w_eco3093, w_eco3094, w_eco3095, w_eco3096, w_eco3097, w_eco3098, w_eco3099, w_eco3100, w_eco3101, w_eco3102, w_eco3103, w_eco3104, w_eco3105, w_eco3106, w_eco3107, w_eco3108, w_eco3109, w_eco3110, w_eco3111, w_eco3112, w_eco3113, w_eco3114, w_eco3115, w_eco3116, w_eco3117, w_eco3118, w_eco3119, w_eco3120, w_eco3121, w_eco3122, w_eco3123, w_eco3124, w_eco3125, w_eco3126, w_eco3127, w_eco3128, w_eco3129, w_eco3130, w_eco3131, w_eco3132, w_eco3133, w_eco3134, w_eco3135, w_eco3136, w_eco3137, w_eco3138, w_eco3139, w_eco3140, w_eco3141, w_eco3142, w_eco3143, w_eco3144, w_eco3145, w_eco3146, w_eco3147, w_eco3148, w_eco3149, w_eco3150, w_eco3151, w_eco3152, w_eco3153, w_eco3154, w_eco3155, w_eco3156, w_eco3157, w_eco3158, w_eco3159, w_eco3160, w_eco3161, w_eco3162, w_eco3163, w_eco3164, w_eco3165, w_eco3166, w_eco3167, w_eco3168, w_eco3169, w_eco3170, w_eco3171, w_eco3172, w_eco3173, w_eco3174, w_eco3175, w_eco3176, w_eco3177, w_eco3178, w_eco3179, w_eco3180, w_eco3181, w_eco3182, w_eco3183, w_eco3184, w_eco3185, w_eco3186, w_eco3187, w_eco3188, w_eco3189, w_eco3190, w_eco3191, w_eco3192, w_eco3193, w_eco3194, w_eco3195, w_eco3196, w_eco3197, w_eco3198, w_eco3199, w_eco3200, w_eco3201, w_eco3202, w_eco3203, w_eco3204, w_eco3205, w_eco3206, w_eco3207, w_eco3208, w_eco3209, w_eco3210, w_eco3211, w_eco3212, w_eco3213, w_eco3214, w_eco3215, w_eco3216, w_eco3217, w_eco3218, w_eco3219, w_eco3220, w_eco3221, w_eco3222, w_eco3223, w_eco3224, w_eco3225, w_eco3226, w_eco3227, w_eco3228, w_eco3229, w_eco3230, w_eco3231, w_eco3232, w_eco3233, w_eco3234, w_eco3235, w_eco3236, w_eco3237, w_eco3238, w_eco3239, w_eco3240, w_eco3241, w_eco3242, w_eco3243, w_eco3244, w_eco3245, w_eco3246, w_eco3247, w_eco3248, w_eco3249, w_eco3250, w_eco3251, w_eco3252, w_eco3253, w_eco3254, w_eco3255, w_eco3256, w_eco3257, w_eco3258, w_eco3259, w_eco3260, w_eco3261, w_eco3262, w_eco3263, w_eco3264, w_eco3265, w_eco3266, w_eco3267, w_eco3268, w_eco3269, w_eco3270, w_eco3271, w_eco3272, w_eco3273, w_eco3274, w_eco3275, w_eco3276, w_eco3277, w_eco3278, w_eco3279, w_eco3280, w_eco3281, w_eco3282, w_eco3283, w_eco3284, w_eco3285, w_eco3286, w_eco3287, w_eco3288, w_eco3289, w_eco3290, w_eco3291, w_eco3292, w_eco3293, w_eco3294, w_eco3295, w_eco3296, w_eco3297, w_eco3298, w_eco3299, w_eco3300, w_eco3301, w_eco3302, w_eco3303, w_eco3304, w_eco3305, w_eco3306, w_eco3307, w_eco3308, w_eco3309, w_eco3310, w_eco3311, w_eco3312, w_eco3313, w_eco3314, w_eco3315, w_eco3316, w_eco3317, w_eco3318, w_eco3319, w_eco3320, w_eco3321, w_eco3322, w_eco3323, w_eco3324, w_eco3325, w_eco3326, w_eco3327, w_eco3328, w_eco3329, w_eco3330, w_eco3331, w_eco3332, w_eco3333, w_eco3334, w_eco3335, w_eco3336, w_eco3337, w_eco3338, w_eco3339, w_eco3340, w_eco3341, w_eco3342, w_eco3343, w_eco3344, w_eco3345, w_eco3346, w_eco3347, w_eco3348, w_eco3349, w_eco3350, w_eco3351, w_eco3352, w_eco3353, w_eco3354, w_eco3355, w_eco3356, w_eco3357, w_eco3358, w_eco3359, w_eco3360, w_eco3361, w_eco3362, w_eco3363, w_eco3364, w_eco3365, w_eco3366, w_eco3367, w_eco3368, w_eco3369, w_eco3370, w_eco3371, w_eco3372, w_eco3373, w_eco3374, w_eco3375, w_eco3376, w_eco3377, w_eco3378, w_eco3379, w_eco3380, w_eco3381, w_eco3382, w_eco3383, w_eco3384, w_eco3385, w_eco3386, w_eco3387, w_eco3388, w_eco3389, w_eco3390, w_eco3391, w_eco3392, w_eco3393, w_eco3394, w_eco3395, w_eco3396, w_eco3397, w_eco3398, w_eco3399, w_eco3400, w_eco3401, w_eco3402, w_eco3403, w_eco3404, w_eco3405, w_eco3406, w_eco3407, w_eco3408, w_eco3409, w_eco3410, w_eco3411, w_eco3412, w_eco3413, w_eco3414, w_eco3415, w_eco3416, w_eco3417, w_eco3418, w_eco3419, w_eco3420, w_eco3421, w_eco3422, w_eco3423, w_eco3424, w_eco3425, w_eco3426, w_eco3427, w_eco3428, w_eco3429, w_eco3430, w_eco3431, w_eco3432, w_eco3433, w_eco3434, w_eco3435, w_eco3436, w_eco3437, w_eco3438, w_eco3439, w_eco3440, w_eco3441, w_eco3442, w_eco3443, w_eco3444, w_eco3445, w_eco3446, w_eco3447, w_eco3448, w_eco3449, w_eco3450, w_eco3451, w_eco3452, w_eco3453, w_eco3454, w_eco3455, w_eco3456, w_eco3457, w_eco3458, w_eco3459, w_eco3460, w_eco3461, w_eco3462, w_eco3463, w_eco3464, w_eco3465, w_eco3466, w_eco3467, w_eco3468, w_eco3469, w_eco3470, w_eco3471, w_eco3472, w_eco3473, w_eco3474, w_eco3475, w_eco3476, w_eco3477, w_eco3478, w_eco3479, w_eco3480, w_eco3481, w_eco3482, w_eco3483, w_eco3484, w_eco3485, w_eco3486, w_eco3487, w_eco3488, w_eco3489, w_eco3490, w_eco3491, w_eco3492, w_eco3493, w_eco3494, w_eco3495, w_eco3496, w_eco3497, w_eco3498, w_eco3499, w_eco3500, w_eco3501, w_eco3502, w_eco3503, w_eco3504, w_eco3505, w_eco3506, w_eco3507, w_eco3508, w_eco3509, w_eco3510, w_eco3511, w_eco3512, w_eco3513, w_eco3514, w_eco3515, w_eco3516, w_eco3517, w_eco3518, w_eco3519, w_eco3520, w_eco3521, w_eco3522, w_eco3523, w_eco3524, w_eco3525, w_eco3526, w_eco3527, w_eco3528, w_eco3529, w_eco3530, w_eco3531, w_eco3532, w_eco3533, w_eco3534, w_eco3535, w_eco3536, w_eco3537, w_eco3538, w_eco3539, w_eco3540, w_eco3541, w_eco3542, w_eco3543, w_eco3544, w_eco3545, w_eco3546, w_eco3547, w_eco3548, w_eco3549, w_eco3550, w_eco3551, w_eco3552, w_eco3553, w_eco3554, w_eco3555, w_eco3556, w_eco3557, w_eco3558, w_eco3559, w_eco3560, w_eco3561, w_eco3562, w_eco3563, w_eco3564, w_eco3565, w_eco3566, w_eco3567, w_eco3568, w_eco3569, w_eco3570, w_eco3571, w_eco3572, w_eco3573, w_eco3574, w_eco3575, w_eco3576, w_eco3577, w_eco3578, w_eco3579, w_eco3580, w_eco3581, w_eco3582, w_eco3583, w_eco3584, w_eco3585, w_eco3586, w_eco3587, w_eco3588, w_eco3589, w_eco3590, w_eco3591, w_eco3592, w_eco3593, w_eco3594, w_eco3595, w_eco3596, w_eco3597, w_eco3598, w_eco3599, w_eco3600, w_eco3601, w_eco3602, w_eco3603, w_eco3604, w_eco3605, w_eco3606, w_eco3607, w_eco3608, w_eco3609, w_eco3610, w_eco3611, w_eco3612, w_eco3613, w_eco3614, w_eco3615, w_eco3616, w_eco3617, w_eco3618, w_eco3619, w_eco3620, w_eco3621, w_eco3622, w_eco3623, w_eco3624, w_eco3625, w_eco3626, w_eco3627, w_eco3628, w_eco3629, w_eco3630, w_eco3631, w_eco3632, w_eco3633, w_eco3634, w_eco3635, w_eco3636, w_eco3637, w_eco3638, w_eco3639, w_eco3640, w_eco3641, w_eco3642, w_eco3643, w_eco3644, w_eco3645, w_eco3646, w_eco3647, w_eco3648, w_eco3649, w_eco3650, w_eco3651, w_eco3652, w_eco3653, w_eco3654, w_eco3655, w_eco3656, w_eco3657, w_eco3658, w_eco3659, w_eco3660, w_eco3661, w_eco3662, w_eco3663, w_eco3664, w_eco3665, w_eco3666, w_eco3667, w_eco3668, w_eco3669, w_eco3670, w_eco3671, w_eco3672, w_eco3673, w_eco3674, w_eco3675, w_eco3676, w_eco3677, w_eco3678, w_eco3679, w_eco3680, w_eco3681, w_eco3682, w_eco3683, w_eco3684, w_eco3685, w_eco3686, w_eco3687, w_eco3688, w_eco3689, w_eco3690, w_eco3691, w_eco3692, w_eco3693, w_eco3694, w_eco3695, w_eco3696, w_eco3697, w_eco3698, w_eco3699, w_eco3700, w_eco3701, w_eco3702, w_eco3703, w_eco3704, w_eco3705, w_eco3706, w_eco3707, w_eco3708, w_eco3709, w_eco3710, w_eco3711, w_eco3712, w_eco3713, w_eco3714, w_eco3715, w_eco3716, w_eco3717, w_eco3718, w_eco3719, w_eco3720, w_eco3721, w_eco3722, w_eco3723, w_eco3724, w_eco3725, w_eco3726, w_eco3727, w_eco3728, w_eco3729, w_eco3730, w_eco3731, w_eco3732, w_eco3733, w_eco3734, w_eco3735, w_eco3736, w_eco3737, w_eco3738, w_eco3739, w_eco3740, w_eco3741, w_eco3742, w_eco3743, w_eco3744, w_eco3745, w_eco3746, w_eco3747, w_eco3748, w_eco3749, w_eco3750, w_eco3751, w_eco3752, w_eco3753, w_eco3754, w_eco3755, w_eco3756, w_eco3757, w_eco3758, w_eco3759, w_eco3760, w_eco3761, w_eco3762, w_eco3763, w_eco3764, w_eco3765, w_eco3766, w_eco3767, w_eco3768, w_eco3769, w_eco3770, w_eco3771, w_eco3772, w_eco3773, w_eco3774, w_eco3775, w_eco3776, w_eco3777, w_eco3778, w_eco3779, w_eco3780, w_eco3781, w_eco3782, w_eco3783, w_eco3784, w_eco3785, w_eco3786, w_eco3787, w_eco3788, w_eco3789, w_eco3790, w_eco3791, w_eco3792, w_eco3793, w_eco3794, w_eco3795, w_eco3796, w_eco3797, w_eco3798, w_eco3799, w_eco3800, w_eco3801, w_eco3802, w_eco3803, w_eco3804, w_eco3805, w_eco3806, w_eco3807, w_eco3808, w_eco3809, w_eco3810, w_eco3811, w_eco3812, w_eco3813, w_eco3814, w_eco3815, w_eco3816, w_eco3817, w_eco3818, w_eco3819, w_eco3820, w_eco3821, w_eco3822, w_eco3823, w_eco3824, w_eco3825, w_eco3826, w_eco3827, w_eco3828, w_eco3829, w_eco3830, w_eco3831, w_eco3832, w_eco3833, w_eco3834, w_eco3835, w_eco3836, w_eco3837, w_eco3838, w_eco3839, w_eco3840, w_eco3841, w_eco3842, w_eco3843, w_eco3844, w_eco3845, w_eco3846, w_eco3847, w_eco3848, w_eco3849, w_eco3850, w_eco3851, w_eco3852, w_eco3853, w_eco3854, w_eco3855, w_eco3856, w_eco3857, w_eco3858, w_eco3859, w_eco3860, w_eco3861, w_eco3862, w_eco3863, w_eco3864, w_eco3865, w_eco3866, w_eco3867, w_eco3868, w_eco3869, w_eco3870, w_eco3871, w_eco3872, w_eco3873, w_eco3874, w_eco3875, w_eco3876, w_eco3877, w_eco3878, w_eco3879, w_eco3880, w_eco3881, w_eco3882, w_eco3883, w_eco3884, w_eco3885, w_eco3886, w_eco3887, w_eco3888, w_eco3889, w_eco3890, w_eco3891, w_eco3892, w_eco3893, w_eco3894, w_eco3895, w_eco3896, w_eco3897, w_eco3898, w_eco3899);
	xor _ECO_out3(cnt[5], sub_wire3, w_eco3900);
	assign w_eco3901 = rst;
	and _ECO_3902(w_eco3902, Tsync[4], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3903(w_eco3903, Tsync[4], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_3904(w_eco3904, Tsync[4], !prev_cnt[3], ena, !prev_state[3], prev_state[1]);
	and _ECO_3905(w_eco3905, Tsync[4], !prev_cnt[3], ena, !prev_state[0]);
	and _ECO_3906(w_eco3906, Tsync[4], !Tsync[3], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_3907(w_eco3907, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_state[1]);
	and _ECO_3908(w_eco3908, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[11], !ena);
	and _ECO_3909(w_eco3909, Tgdel[4], prev_cnt[1], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3910(w_eco3910, Tgdel[4], prev_cnt[1], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3911(w_eco3911, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_state[3], !prev_state[2]);
	and _ECO_3912(w_eco3912, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_3913(w_eco3913, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_state[4], !prev_state[2]);
	and _ECO_3914(w_eco3914, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[15], !ena);
	and _ECO_3915(w_eco3915, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[11], !ena);
	and _ECO_3916(w_eco3916, Tgdel[4], !Tsync[3], prev_cnt[1], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_3917(w_eco3917, Tgdel[4], prev_cnt[2], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3918(w_eco3918, Tgate[4], prev_cnt[1], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3919(w_eco3919, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3920(w_eco3920, !Tsync[3], prev_cnt[1], prev_cnt[4], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_3921(w_eco3921, Tgdel[4], prev_cnt[2], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3922(w_eco3922, Tgate[4], prev_cnt[1], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3923(w_eco3923, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3924(w_eco3924, !Tsync[4], prev_cnt[3], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3925(w_eco3925, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_3926(w_eco3926, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], prev_state[1]);
	and _ECO_3927(w_eco3927, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_3928(w_eco3928, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_3929(w_eco3929, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[0]);
	and _ECO_3930(w_eco3930, Tgate[4], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_3931(w_eco3931, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_3932(w_eco3932, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[15], !ena);
	and _ECO_3933(w_eco3933, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[1], !prev_cnt[4], !ena);
	and _ECO_3934(w_eco3934, Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_3935(w_eco3935, Tgdel[4], !Tsync[3], prev_cnt[2], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_3936(w_eco3936, Tgdel[4], prev_cnt[3], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3937(w_eco3937, prev_cnt[1], prev_cnt[4], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3938(w_eco3938, Tgate[4], prev_cnt[2], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3939(w_eco3939, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], !ena);
	and _ECO_3940(w_eco3940, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3941(w_eco3941, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_3942(w_eco3942, !Tsync[3], prev_cnt[2], prev_cnt[4], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_3943(w_eco3943, Tgdel[4], prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3944(w_eco3944, prev_cnt[1], prev_cnt[4], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3945(w_eco3945, Tgate[4], prev_cnt[2], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3946(w_eco3946, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3947(w_eco3947, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_3948(w_eco3948, !Tsync[4], prev_cnt[3], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3949(w_eco3949, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_3950(w_eco3950, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], prev_state[1]);
	and _ECO_3951(w_eco3951, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_3952(w_eco3952, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_3953(w_eco3953, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_3954(w_eco3954, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[0]);
	and _ECO_3955(w_eco3955, Tgate[4], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_3956(w_eco3956, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_3957(w_eco3957, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[9], !ena);
	and _ECO_3958(w_eco3958, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[11], !ena);
	and _ECO_3959(w_eco3959, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !ena);
	and _ECO_3960(w_eco3960, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[2], !prev_cnt[4], !ena);
	and _ECO_3961(w_eco3961, Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_3962(w_eco3962, Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_3963(w_eco3963, Tgdel[4], !Tsync[3], prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_3964(w_eco3964, Tgdel[4], prev_cnt[0], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3965(w_eco3965, Tgdel[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3966(w_eco3966, prev_cnt[1], prev_cnt[4], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3967(w_eco3967, prev_cnt[2], prev_cnt[4], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3968(w_eco3968, Tgate[4], prev_cnt[3], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3969(w_eco3969, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], !ena);
	and _ECO_3970(w_eco3970, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3971(w_eco3971, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3972(w_eco3972, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_3973(w_eco3973, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_3974(w_eco3974, !Tsync[3], prev_cnt[3], prev_cnt[4], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_3975(w_eco3975, Tgate[4], !Tsync[3], prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_3976(w_eco3976, !Tsync[3], prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_3977(w_eco3977, Tgdel[4], prev_cnt[0], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3978(w_eco3978, Tgdel[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3979(w_eco3979, prev_cnt[1], prev_cnt[4], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3980(w_eco3980, prev_cnt[2], prev_cnt[4], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3981(w_eco3981, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3982(w_eco3982, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_3983(w_eco3983, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_3984(w_eco3984, !Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_3985(w_eco3985, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_3986(w_eco3986, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_3987(w_eco3987, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_3988(w_eco3988, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_state[1]);
	and _ECO_3989(w_eco3989, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_3990(w_eco3990, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_3991(w_eco3991, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_3992(w_eco3992, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_3993(w_eco3993, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[0]);
	and _ECO_3994(w_eco3994, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[0]);
	and _ECO_3995(w_eco3995, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[6], !ena);
	and _ECO_3996(w_eco3996, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[9], !ena);
	and _ECO_3997(w_eco3997, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[15], !ena);
	and _ECO_3998(w_eco3998, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !ena);
	and _ECO_3999(w_eco3999, Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4000(w_eco4000, Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4001(w_eco4001, !Tgate[4], !Tgdel[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4002(w_eco4002, prev_cnt[2], prev_cnt[4], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4003(w_eco4003, prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4004(w_eco4004, Tgate[4], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4005(w_eco4005, Tgate[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4006(w_eco4006, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], !ena);
	and _ECO_4007(w_eco4007, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4008(w_eco4008, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], prev_state[0]);
	and _ECO_4009(w_eco4009, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4010(w_eco4010, prev_cnt[2], prev_cnt[4], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4011(w_eco4011, Tgate[4], prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4012(w_eco4012, prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4013(w_eco4013, Tgate[4], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4014(w_eco4014, Tgate[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4015(w_eco4015, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], !prev_state[4], !prev_state[2]);
	and _ECO_4016(w_eco4016, !Tsync[4], prev_cnt[3], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4017(w_eco4017, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4018(w_eco4018, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], prev_state[1]);
	and _ECO_4019(w_eco4019, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_4020(w_eco4020, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4021(w_eco4021, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4022(w_eco4022, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4023(w_eco4023, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4024(w_eco4024, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_4025(w_eco4025, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_4026(w_eco4026, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_4027(w_eco4027, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_state[3], prev_state[0]);
	and _ECO_4028(w_eco4028, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_4029(w_eco4029, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_4030(w_eco4030, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[8], !ena);
	and _ECO_4031(w_eco4031, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[6], !ena);
	and _ECO_4032(w_eco4032, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[0], !prev_cnt[4], !ena);
	and _ECO_4033(w_eco4033, !Tgate[4], !Tgdel[4], !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], !ena);
	and _ECO_4034(w_eco4034, prev_cnt[1], prev_cnt[4], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4035(w_eco4035, prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4036(w_eco4036, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4037(w_eco4037, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], !ena);
	and _ECO_4038(w_eco4038, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4039(w_eco4039, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], prev_state[0]);
	and _ECO_4040(w_eco4040, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4041(w_eco4041, prev_cnt[1], prev_cnt[4], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4042(w_eco4042, prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4043(w_eco4043, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4044(w_eco4044, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_4045(w_eco4045, !Tsync[4], prev_cnt[3], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4046(w_eco4046, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], prev_state[1]);
	and _ECO_4047(w_eco4047, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4048(w_eco4048, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4049(w_eco4049, !Tgate[4], !Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], !prev_state[3], prev_state[0]);
	and _ECO_4050(w_eco4050, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4051(w_eco4051, Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4052(w_eco4052, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4053(w_eco4053, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4054(w_eco4054, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_4055(w_eco4055, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_4056(w_eco4056, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_4057(w_eco4057, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_state[3], prev_state[0]);
	and _ECO_4058(w_eco4058, !Tsync[4], prev_cnt[1], !prev_cnt[4], prev_cnt[10], !ena);
	and _ECO_4059(w_eco4059, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[8], !ena);
	and _ECO_4060(w_eco4060, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[9], !ena);
	and _ECO_4061(w_eco4061, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !ena);
	and _ECO_4062(w_eco4062, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4063(w_eco4063, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4064(w_eco4064, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4065(w_eco4065, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4066(w_eco4066, prev_cnt[1], prev_cnt[4], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4067(w_eco4067, prev_cnt[2], prev_cnt[4], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4068(w_eco4068, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4069(w_eco4069, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4070(w_eco4070, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], !ena);
	and _ECO_4071(w_eco4071, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4072(w_eco4072, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4073(w_eco4073, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_state[0]);
	and _ECO_4074(w_eco4074, Tgdel[4], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4075(w_eco4075, prev_cnt[1], prev_cnt[4], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4076(w_eco4076, prev_cnt[2], prev_cnt[4], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4077(w_eco4077, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4078(w_eco4078, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4079(w_eco4079, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_4080(w_eco4080, !Tsync[4], prev_cnt[3], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4081(w_eco4081, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], prev_state[1]);
	and _ECO_4082(w_eco4082, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_4083(w_eco4083, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4084(w_eco4084, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4085(w_eco4085, Tgdel[4], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4086(w_eco4086, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4087(w_eco4087, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4088(w_eco4088, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_4089(w_eco4089, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_4090(w_eco4090, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_state[3], prev_state[0]);
	and _ECO_4091(w_eco4091, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_state[3], prev_state[0]);
	and _ECO_4092(w_eco4092, !Tsync[4], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], !ena);
	and _ECO_4093(w_eco4093, !Tsync[4], prev_cnt[2], !prev_cnt[4], prev_cnt[10], !ena);
	and _ECO_4094(w_eco4094, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[6], !ena);
	and _ECO_4095(w_eco4095, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !ena);
	and _ECO_4096(w_eco4096, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4097(w_eco4097, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4098(w_eco4098, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4099(w_eco4099, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4100(w_eco4100, Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4101(w_eco4101, Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4102(w_eco4102, Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4103(w_eco4103, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4104(w_eco4104, prev_cnt[1], prev_cnt[4], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4105(w_eco4105, prev_cnt[2], prev_cnt[4], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4106(w_eco4106, prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4107(w_eco4107, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4108(w_eco4108, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], !ena);
	and _ECO_4109(w_eco4109, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4110(w_eco4110, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4111(w_eco4111, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], prev_state[0]);
	and _ECO_4112(w_eco4112, Tgdel[4], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4113(w_eco4113, prev_cnt[14], prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4114(w_eco4114, prev_cnt[1], prev_cnt[4], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4115(w_eco4115, prev_cnt[2], prev_cnt[4], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4116(w_eco4116, prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4117(w_eco4117, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4118(w_eco4118, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_4119(w_eco4119, !Tsync[4], prev_cnt[3], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4120(w_eco4120, Tgdel[4], prev_cnt[14], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4121(w_eco4121, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4122(w_eco4122, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4123(w_eco4123, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], prev_state[1]);
	and _ECO_4124(w_eco4124, Tgdel[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_4125(w_eco4125, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_4126(w_eco4126, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4127(w_eco4127, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4128(w_eco4128, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4129(w_eco4129, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4130(w_eco4130, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4131(w_eco4131, Tgdel[4], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4132(w_eco4132, prev_cnt[14], prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4133(w_eco4133, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4134(w_eco4134, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4135(w_eco4135, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_4136(w_eco4136, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_4137(w_eco4137, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_4138(w_eco4138, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_4139(w_eco4139, !Tsync[4], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], !ena);
	and _ECO_4140(w_eco4140, !Tsync[4], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], !ena);
	and _ECO_4141(w_eco4141, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[8], !ena);
	and _ECO_4142(w_eco4142, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !ena);
	and _ECO_4143(w_eco4143, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4144(w_eco4144, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4145(w_eco4145, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4146(w_eco4146, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4147(w_eco4147, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4148(w_eco4148, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4149(w_eco4149, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4150(w_eco4150, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4151(w_eco4151, Tgate[4], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4152(w_eco4152, prev_cnt[1], prev_cnt[4], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4153(w_eco4153, prev_cnt[2], prev_cnt[4], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4154(w_eco4154, prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4155(w_eco4155, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4156(w_eco4156, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4157(w_eco4157, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], !ena);
	and _ECO_4158(w_eco4158, Tgdel[4], prev_cnt[14], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4159(w_eco4159, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4160(w_eco4160, Tgdel[4], !Tsync[3], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_4161(w_eco4161, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4162(w_eco4162, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], prev_state[0]);
	and _ECO_4163(w_eco4163, Tgdel[4], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4164(w_eco4164, Tgdel[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4165(w_eco4165, prev_cnt[14], prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4166(w_eco4166, Tgate[4], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4167(w_eco4167, prev_cnt[1], prev_cnt[4], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4168(w_eco4168, prev_cnt[2], prev_cnt[4], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4169(w_eco4169, prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4170(w_eco4170, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4171(w_eco4171, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4172(w_eco4172, Tgdel[4], prev_cnt[14], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4173(w_eco4173, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_4174(w_eco4174, !Tsync[4], !prev_cnt[14], prev_cnt[3], prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4175(w_eco4175, Tgdel[4], prev_cnt[14], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4176(w_eco4176, prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4177(w_eco4177, Tgdel[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_4178(w_eco4178, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4179(w_eco4179, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4180(w_eco4180, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], prev_state[1]);
	and _ECO_4181(w_eco4181, Tgate[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_4182(w_eco4182, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_4183(w_eco4183, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4184(w_eco4184, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4185(w_eco4185, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_4186(w_eco4186, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4187(w_eco4187, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4188(w_eco4188, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4189(w_eco4189, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4190(w_eco4190, Tgdel[4], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4191(w_eco4191, Tgdel[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4192(w_eco4192, prev_cnt[14], prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4193(w_eco4193, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4194(w_eco4194, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4195(w_eco4195, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4196(w_eco4196, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4197(w_eco4197, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4198(w_eco4198, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_4199(w_eco4199, Tgdel[4], !Tsync[3], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_4200(w_eco4200, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_4201(w_eco4201, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_4202(w_eco4202, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_4203(w_eco4203, !Tsync[4], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], !ena);
	and _ECO_4204(w_eco4204, !Tsync[4], prev_cnt[0], !prev_cnt[4], prev_cnt[10], !ena);
	and _ECO_4205(w_eco4205, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !ena);
	and _ECO_4206(w_eco4206, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4207(w_eco4207, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4208(w_eco4208, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4209(w_eco4209, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4210(w_eco4210, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4211(w_eco4211, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4212(w_eco4212, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4213(w_eco4213, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4214(w_eco4214, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4215(w_eco4215, !prev_cnt[14], prev_cnt[1], prev_cnt[4], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4216(w_eco4216, prev_cnt[2], prev_cnt[4], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4217(w_eco4217, prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4218(w_eco4218, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4219(w_eco4219, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4220(w_eco4220, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], !ena);
	and _ECO_4221(w_eco4221, Tgdel[4], prev_cnt[14], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4222(w_eco4222, Tgate[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4223(w_eco4223, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4224(w_eco4224, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], prev_state[0]);
	and _ECO_4225(w_eco4225, Tgate[4], !Tsync[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_4226(w_eco4226, Tgdel[4], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4227(w_eco4227, Tgdel[4], prev_cnt[14], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4228(w_eco4228, prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4229(w_eco4229, prev_cnt[14], prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4230(w_eco4230, !prev_cnt[14], prev_cnt[1], prev_cnt[4], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4231(w_eco4231, prev_cnt[2], prev_cnt[4], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4232(w_eco4232, prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4233(w_eco4233, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4234(w_eco4234, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4235(w_eco4235, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_4236(w_eco4236, !Tsync[4], !prev_cnt[14], prev_cnt[3], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4237(w_eco4237, Tgdel[4], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4238(w_eco4238, prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4239(w_eco4239, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4240(w_eco4240, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4241(w_eco4241, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4242(w_eco4242, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4243(w_eco4243, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], prev_state[1]);
	and _ECO_4244(w_eco4244, Tgdel[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_4245(w_eco4245, !Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_4246(w_eco4246, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4247(w_eco4247, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4248(w_eco4248, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4249(w_eco4249, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_4250(w_eco4250, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4251(w_eco4251, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4252(w_eco4252, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4253(w_eco4253, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4254(w_eco4254, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4255(w_eco4255, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4256(w_eco4256, Tgdel[4], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4257(w_eco4257, prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4258(w_eco4258, prev_cnt[14], prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4259(w_eco4259, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4260(w_eco4260, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4261(w_eco4261, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4262(w_eco4262, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4263(w_eco4263, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4264(w_eco4264, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4265(w_eco4265, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_4266(w_eco4266, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_4267(w_eco4267, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_4268(w_eco4268, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_4269(w_eco4269, Tgate[4], !Tsync[3], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_4270(w_eco4270, !Tgate[4], Tgdel[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[0]);
	and _ECO_4271(w_eco4271, !Tsync[4], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], !ena);
	and _ECO_4272(w_eco4272, !Tsync[4], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !ena);
	and _ECO_4273(w_eco4273, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4274(w_eco4274, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4275(w_eco4275, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4276(w_eco4276, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4277(w_eco4277, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4278(w_eco4278, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4279(w_eco4279, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4280(w_eco4280, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4281(w_eco4281, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4282(w_eco4282, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4283(w_eco4283, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4284(w_eco4284, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4285(w_eco4285, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4286(w_eco4286, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4287(w_eco4287, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4288(w_eco4288, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4289(w_eco4289, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4290(w_eco4290, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4291(w_eco4291, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4292(w_eco4292, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4293(w_eco4293, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4294(w_eco4294, Tgate[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4295(w_eco4295, !prev_cnt[14], prev_cnt[1], prev_cnt[4], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4296(w_eco4296, !prev_cnt[14], prev_cnt[2], prev_cnt[4], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4297(w_eco4297, prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4298(w_eco4298, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4299(w_eco4299, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4300(w_eco4300, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], !ena);
	and _ECO_4301(w_eco4301, Tgdel[4], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4302(w_eco4302, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4303(w_eco4303, Tgdel[4], !Tsync[3], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_4304(w_eco4304, Tgdel[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_4305(w_eco4305, Tgdel[4], prev_cnt[14], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4306(w_eco4306, prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4307(w_eco4307, prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4308(w_eco4308, Tgdel[4], !Tsync[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_4309(w_eco4309, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4310(w_eco4310, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4311(w_eco4311, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4312(w_eco4312, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4313(w_eco4313, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4314(w_eco4314, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4315(w_eco4315, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4316(w_eco4316, Tgate[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4317(w_eco4317, !prev_cnt[14], prev_cnt[1], prev_cnt[4], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4318(w_eco4318, !prev_cnt[14], prev_cnt[2], prev_cnt[4], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4319(w_eco4319, prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4320(w_eco4320, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4321(w_eco4321, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4322(w_eco4322, Tgdel[4], prev_cnt[1], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4323(w_eco4323, Tgdel[4], prev_cnt[14], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4324(w_eco4324, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_4325(w_eco4325, Tgdel[4], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4326(w_eco4326, prev_cnt[1], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4327(w_eco4327, Tgdel[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_4328(w_eco4328, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4329(w_eco4329, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4330(w_eco4330, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4331(w_eco4331, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4332(w_eco4332, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4333(w_eco4333, Tgate[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_4334(w_eco4334, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_4335(w_eco4335, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4336(w_eco4336, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_4337(w_eco4337, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_4338(w_eco4338, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4339(w_eco4339, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_4340(w_eco4340, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4341(w_eco4341, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4342(w_eco4342, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4343(w_eco4343, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4344(w_eco4344, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_4345(w_eco4345, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4346(w_eco4346, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4347(w_eco4347, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4348(w_eco4348, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4349(w_eco4349, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4350(w_eco4350, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4351(w_eco4351, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4352(w_eco4352, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4353(w_eco4353, Tgdel[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4354(w_eco4354, prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4355(w_eco4355, prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4356(w_eco4356, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4357(w_eco4357, Tgdel[4], Tsync[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2]);
	and _ECO_4358(w_eco4358, Tgdel[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4359(w_eco4359, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4360(w_eco4360, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4361(w_eco4361, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4362(w_eco4362, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4363(w_eco4363, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4364(w_eco4364, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4365(w_eco4365, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_4366(w_eco4366, Tgdel[4], !Tsync[3], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_4367(w_eco4367, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_4368(w_eco4368, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_4369(w_eco4369, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_4370(w_eco4370, !Tsync[4], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], !ena);
	and _ECO_4371(w_eco4371, !Tsync[4], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !ena);
	and _ECO_4372(w_eco4372, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4373(w_eco4373, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4374(w_eco4374, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4375(w_eco4375, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4376(w_eco4376, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4377(w_eco4377, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4378(w_eco4378, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4379(w_eco4379, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4380(w_eco4380, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4381(w_eco4381, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4382(w_eco4382, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4383(w_eco4383, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4384(w_eco4384, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4385(w_eco4385, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4386(w_eco4386, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4387(w_eco4387, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4388(w_eco4388, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4389(w_eco4389, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4390(w_eco4390, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4391(w_eco4391, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4392(w_eco4392, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4393(w_eco4393, !prev_cnt[14], prev_cnt[2], prev_cnt[4], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4394(w_eco4394, !prev_cnt[14], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4395(w_eco4395, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4396(w_eco4396, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4397(w_eco4397, Tgdel[4], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4398(w_eco4398, Tgdel[4], prev_cnt[14], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4399(w_eco4399, Tgdel[4], prev_cnt[14], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4400(w_eco4400, Tgate[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_4401(w_eco4401, !Tgate[4], Tgdel[4], !Tsync[4], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[0]);
	and _ECO_4402(w_eco4402, Tgdel[4], !Tsync[3], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_4403(w_eco4403, !Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], prev_state[0]);
	and _ECO_4404(w_eco4404, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], prev_state[0]);
	and _ECO_4405(w_eco4405, Tgate[4], !Tsync[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_4406(w_eco4406, Tgdel[4], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4407(w_eco4407, Tgdel[4], prev_cnt[14], !prev_cnt[3], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4408(w_eco4408, prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4409(w_eco4409, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4410(w_eco4410, Tgate[4], !Tsync[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_4411(w_eco4411, !prev_cnt[14], prev_cnt[2], prev_cnt[4], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4412(w_eco4412, !prev_cnt[14], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4413(w_eco4413, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4414(w_eco4414, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4415(w_eco4415, Tgdel[4], prev_cnt[14], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4416(w_eco4416, Tgdel[4], prev_cnt[14], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4417(w_eco4417, prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4418(w_eco4418, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4419(w_eco4419, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4420(w_eco4420, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4421(w_eco4421, Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4422(w_eco4422, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4423(w_eco4423, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4424(w_eco4424, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4425(w_eco4425, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4426(w_eco4426, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4427(w_eco4427, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4428(w_eco4428, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4429(w_eco4429, !Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_4430(w_eco4430, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4431(w_eco4431, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4432(w_eco4432, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4433(w_eco4433, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4434(w_eco4434, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_4435(w_eco4435, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_4436(w_eco4436, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4437(w_eco4437, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4438(w_eco4438, prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4439(w_eco4439, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4440(w_eco4440, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4441(w_eco4441, Tgate[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4442(w_eco4442, Tgdel[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4443(w_eco4443, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4444(w_eco4444, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4445(w_eco4445, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4446(w_eco4446, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4447(w_eco4447, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4448(w_eco4448, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4449(w_eco4449, Tgate[4], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_4450(w_eco4450, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4451(w_eco4451, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4452(w_eco4452, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4453(w_eco4453, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4454(w_eco4454, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4455(w_eco4455, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4456(w_eco4456, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4457(w_eco4457, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4458(w_eco4458, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4459(w_eco4459, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4460(w_eco4460, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4461(w_eco4461, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4462(w_eco4462, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4463(w_eco4463, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4464(w_eco4464, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_4465(w_eco4465, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_4466(w_eco4466, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_4467(w_eco4467, Tgate[4], !Tsync[3], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_4468(w_eco4468, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4469(w_eco4469, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4470(w_eco4470, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4471(w_eco4471, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4472(w_eco4472, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4473(w_eco4473, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4474(w_eco4474, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4475(w_eco4475, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4476(w_eco4476, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4477(w_eco4477, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4478(w_eco4478, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4479(w_eco4479, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4480(w_eco4480, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4481(w_eco4481, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4482(w_eco4482, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4483(w_eco4483, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4484(w_eco4484, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4485(w_eco4485, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4486(w_eco4486, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4487(w_eco4487, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4488(w_eco4488, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4489(w_eco4489, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4490(w_eco4490, !prev_cnt[14], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4491(w_eco4491, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4492(w_eco4492, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4493(w_eco4493, Tgdel[4], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4494(w_eco4494, Tgdel[4], prev_cnt[14], !prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_4495(w_eco4495, prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4496(w_eco4496, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4497(w_eco4497, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4498(w_eco4498, Tgdel[4], !Tsync[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_4499(w_eco4499, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4500(w_eco4500, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4501(w_eco4501, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4502(w_eco4502, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4503(w_eco4503, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4504(w_eco4504, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4505(w_eco4505, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4506(w_eco4506, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4507(w_eco4507, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4508(w_eco4508, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4509(w_eco4509, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4510(w_eco4510, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4511(w_eco4511, !prev_cnt[14], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4512(w_eco4512, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4513(w_eco4513, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4514(w_eco4514, Tgdel[4], prev_cnt[2], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4515(w_eco4515, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4516(w_eco4516, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4517(w_eco4517, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4518(w_eco4518, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4519(w_eco4519, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4520(w_eco4520, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4521(w_eco4521, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4522(w_eco4522, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4523(w_eco4523, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4524(w_eco4524, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4525(w_eco4525, Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_4526(w_eco4526, Tgate[4], !Tsync[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_4527(w_eco4527, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4528(w_eco4528, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4529(w_eco4529, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4530(w_eco4530, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4531(w_eco4531, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_4532(w_eco4532, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_4533(w_eco4533, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_4534(w_eco4534, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_4535(w_eco4535, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4536(w_eco4536, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4537(w_eco4537, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4538(w_eco4538, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4539(w_eco4539, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4540(w_eco4540, prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4541(w_eco4541, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4542(w_eco4542, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4543(w_eco4543, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4544(w_eco4544, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4545(w_eco4545, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4546(w_eco4546, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4547(w_eco4547, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4548(w_eco4548, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4549(w_eco4549, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4550(w_eco4550, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4551(w_eco4551, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4552(w_eco4552, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4553(w_eco4553, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4554(w_eco4554, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4555(w_eco4555, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4556(w_eco4556, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4557(w_eco4557, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_4558(w_eco4558, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_4559(w_eco4559, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4560(w_eco4560, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4561(w_eco4561, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4562(w_eco4562, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4563(w_eco4563, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4564(w_eco4564, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4565(w_eco4565, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4566(w_eco4566, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4567(w_eco4567, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4568(w_eco4568, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4569(w_eco4569, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4570(w_eco4570, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4571(w_eco4571, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4572(w_eco4572, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4573(w_eco4573, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4574(w_eco4574, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4575(w_eco4575, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4576(w_eco4576, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4577(w_eco4577, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4578(w_eco4578, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4579(w_eco4579, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4580(w_eco4580, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4581(w_eco4581, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4582(w_eco4582, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4583(w_eco4583, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4584(w_eco4584, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4585(w_eco4585, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4586(w_eco4586, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4587(w_eco4587, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4588(w_eco4588, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4589(w_eco4589, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4590(w_eco4590, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4591(w_eco4591, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4592(w_eco4592, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4593(w_eco4593, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4594(w_eco4594, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4595(w_eco4595, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4596(w_eco4596, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4597(w_eco4597, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4598(w_eco4598, Tgdel[4], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4599(w_eco4599, Tgdel[4], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_4600(w_eco4600, Tgdel[4], !Tsync[3], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_4601(w_eco4601, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], prev_state[0]);
	and _ECO_4602(w_eco4602, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_4603(w_eco4603, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4604(w_eco4604, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4605(w_eco4605, Tgdel[4], prev_cnt[0], !prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4606(w_eco4606, Tgdel[4], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_4607(w_eco4607, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_4608(w_eco4608, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_4609(w_eco4609, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4610(w_eco4610, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_4611(w_eco4611, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4612(w_eco4612, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4613(w_eco4613, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4614(w_eco4614, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4615(w_eco4615, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4616(w_eco4616, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4617(w_eco4617, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4618(w_eco4618, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4619(w_eco4619, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4620(w_eco4620, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4621(w_eco4621, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4622(w_eco4622, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4623(w_eco4623, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4624(w_eco4624, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4625(w_eco4625, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4626(w_eco4626, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4627(w_eco4627, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4628(w_eco4628, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4629(w_eco4629, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4630(w_eco4630, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4631(w_eco4631, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4632(w_eco4632, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_4633(w_eco4633, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4634(w_eco4634, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4635(w_eco4635, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4636(w_eco4636, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4637(w_eco4637, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4638(w_eco4638, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_4639(w_eco4639, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_4640(w_eco4640, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_4641(w_eco4641, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4642(w_eco4642, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4643(w_eco4643, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4644(w_eco4644, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_4645(w_eco4645, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4646(w_eco4646, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4647(w_eco4647, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4648(w_eco4648, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4649(w_eco4649, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4650(w_eco4650, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4651(w_eco4651, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4652(w_eco4652, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4653(w_eco4653, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4654(w_eco4654, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4655(w_eco4655, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4656(w_eco4656, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4657(w_eco4657, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4658(w_eco4658, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4659(w_eco4659, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4660(w_eco4660, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4661(w_eco4661, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4662(w_eco4662, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_4663(w_eco4663, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_4664(w_eco4664, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4665(w_eco4665, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4666(w_eco4666, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4667(w_eco4667, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4668(w_eco4668, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4669(w_eco4669, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4670(w_eco4670, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4671(w_eco4671, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4672(w_eco4672, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4673(w_eco4673, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4674(w_eco4674, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4675(w_eco4675, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4676(w_eco4676, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4677(w_eco4677, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4678(w_eco4678, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4679(w_eco4679, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4680(w_eco4680, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4681(w_eco4681, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4682(w_eco4682, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4683(w_eco4683, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4684(w_eco4684, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4685(w_eco4685, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4686(w_eco4686, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4687(w_eco4687, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4688(w_eco4688, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4689(w_eco4689, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4690(w_eco4690, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4691(w_eco4691, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4692(w_eco4692, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4693(w_eco4693, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4694(w_eco4694, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4695(w_eco4695, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4696(w_eco4696, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4697(w_eco4697, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_4698(w_eco4698, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_4699(w_eco4699, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_4700(w_eco4700, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4701(w_eco4701, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4702(w_eco4702, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4703(w_eco4703, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4704(w_eco4704, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4705(w_eco4705, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4706(w_eco4706, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4707(w_eco4707, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4708(w_eco4708, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4709(w_eco4709, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4710(w_eco4710, prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4711(w_eco4711, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4712(w_eco4712, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4713(w_eco4713, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4714(w_eco4714, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4715(w_eco4715, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4716(w_eco4716, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4717(w_eco4717, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4718(w_eco4718, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_4719(w_eco4719, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4720(w_eco4720, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4721(w_eco4721, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_4722(w_eco4722, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4723(w_eco4723, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4724(w_eco4724, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4725(w_eco4725, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4726(w_eco4726, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4727(w_eco4727, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4728(w_eco4728, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4729(w_eco4729, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4730(w_eco4730, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4731(w_eco4731, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4732(w_eco4732, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4733(w_eco4733, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4734(w_eco4734, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4735(w_eco4735, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4736(w_eco4736, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4737(w_eco4737, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4738(w_eco4738, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4739(w_eco4739, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4740(w_eco4740, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4741(w_eco4741, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4742(w_eco4742, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4743(w_eco4743, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4744(w_eco4744, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4745(w_eco4745, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4746(w_eco4746, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4747(w_eco4747, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4748(w_eco4748, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4749(w_eco4749, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4750(w_eco4750, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4751(w_eco4751, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4752(w_eco4752, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4753(w_eco4753, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4754(w_eco4754, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4755(w_eco4755, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4756(w_eco4756, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4757(w_eco4757, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4758(w_eco4758, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4759(w_eco4759, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4760(w_eco4760, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4761(w_eco4761, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4762(w_eco4762, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4763(w_eco4763, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4764(w_eco4764, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4765(w_eco4765, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4766(w_eco4766, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4767(w_eco4767, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4768(w_eco4768, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4769(w_eco4769, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4770(w_eco4770, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4771(w_eco4771, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4772(w_eco4772, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4773(w_eco4773, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4774(w_eco4774, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4775(w_eco4775, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4776(w_eco4776, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4777(w_eco4777, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4778(w_eco4778, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4779(w_eco4779, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4780(w_eco4780, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4781(w_eco4781, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4782(w_eco4782, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4783(w_eco4783, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4784(w_eco4784, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4785(w_eco4785, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4786(w_eco4786, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4787(w_eco4787, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4788(w_eco4788, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4789(w_eco4789, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4790(w_eco4790, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4791(w_eco4791, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4792(w_eco4792, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4793(w_eco4793, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4794(w_eco4794, Tsync[4], !Tsync[3], !prev_cnt[3], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4795(w_eco4795, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_4796(w_eco4796, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_4797(w_eco4797, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4798(w_eco4798, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4799(w_eco4799, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4800(w_eco4800, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4801(w_eco4801, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4802(w_eco4802, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4803(w_eco4803, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4804(w_eco4804, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4805(w_eco4805, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4806(w_eco4806, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4807(w_eco4807, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4808(w_eco4808, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4809(w_eco4809, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4810(w_eco4810, prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4811(w_eco4811, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4812(w_eco4812, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4813(w_eco4813, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4814(w_eco4814, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4815(w_eco4815, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4816(w_eco4816, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4817(w_eco4817, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4818(w_eco4818, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_4819(w_eco4819, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4820(w_eco4820, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4821(w_eco4821, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4822(w_eco4822, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4823(w_eco4823, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4824(w_eco4824, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4825(w_eco4825, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4826(w_eco4826, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4827(w_eco4827, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4828(w_eco4828, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4829(w_eco4829, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4830(w_eco4830, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4831(w_eco4831, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4832(w_eco4832, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4833(w_eco4833, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4834(w_eco4834, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4835(w_eco4835, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4836(w_eco4836, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4837(w_eco4837, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4838(w_eco4838, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4839(w_eco4839, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4840(w_eco4840, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4841(w_eco4841, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4842(w_eco4842, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4843(w_eco4843, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4844(w_eco4844, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4845(w_eco4845, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4846(w_eco4846, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4847(w_eco4847, Tsync[4], !Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4848(w_eco4848, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4849(w_eco4849, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4850(w_eco4850, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4851(w_eco4851, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4852(w_eco4852, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4853(w_eco4853, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4854(w_eco4854, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4855(w_eco4855, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4856(w_eco4856, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4857(w_eco4857, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4858(w_eco4858, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4859(w_eco4859, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4860(w_eco4860, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4861(w_eco4861, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4862(w_eco4862, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4863(w_eco4863, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4864(w_eco4864, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4865(w_eco4865, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4866(w_eco4866, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4867(w_eco4867, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4868(w_eco4868, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4869(w_eco4869, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4870(w_eco4870, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4871(w_eco4871, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4872(w_eco4872, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4873(w_eco4873, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4874(w_eco4874, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4875(w_eco4875, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4876(w_eco4876, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4877(w_eco4877, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4878(w_eco4878, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4879(w_eco4879, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4880(w_eco4880, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4881(w_eco4881, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4882(w_eco4882, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4883(w_eco4883, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4884(w_eco4884, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4885(w_eco4885, Tsync[4], !Tsync[3], !prev_cnt[3], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4886(w_eco4886, Tsync[4], !Tsync[3], !prev_cnt[3], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4887(w_eco4887, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4888(w_eco4888, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4889(w_eco4889, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4890(w_eco4890, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4891(w_eco4891, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4892(w_eco4892, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4893(w_eco4893, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4894(w_eco4894, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4895(w_eco4895, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4896(w_eco4896, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4897(w_eco4897, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4898(w_eco4898, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_4899(w_eco4899, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_4900(w_eco4900, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4901(w_eco4901, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4902(w_eco4902, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4903(w_eco4903, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_4904(w_eco4904, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4905(w_eco4905, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4906(w_eco4906, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4907(w_eco4907, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4908(w_eco4908, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4909(w_eco4909, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4910(w_eco4910, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4911(w_eco4911, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4912(w_eco4912, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4913(w_eco4913, !Tgate[4], !Tgdel[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4914(w_eco4914, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4915(w_eco4915, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4916(w_eco4916, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4917(w_eco4917, Tsync[4], !prev_cnt[3], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4918(w_eco4918, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4919(w_eco4919, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4920(w_eco4920, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4921(w_eco4921, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4922(w_eco4922, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4923(w_eco4923, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4924(w_eco4924, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_4925(w_eco4925, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4926(w_eco4926, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_4927(w_eco4927, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4928(w_eco4928, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4929(w_eco4929, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4930(w_eco4930, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4931(w_eco4931, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4932(w_eco4932, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4933(w_eco4933, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4934(w_eco4934, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4935(w_eco4935, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4936(w_eco4936, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4937(w_eco4937, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4938(w_eco4938, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4939(w_eco4939, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4940(w_eco4940, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4941(w_eco4941, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4942(w_eco4942, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4943(w_eco4943, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4944(w_eco4944, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4945(w_eco4945, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4946(w_eco4946, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4947(w_eco4947, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4948(w_eco4948, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4949(w_eco4949, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4950(w_eco4950, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4951(w_eco4951, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4952(w_eco4952, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4953(w_eco4953, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4954(w_eco4954, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4955(w_eco4955, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4956(w_eco4956, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4957(w_eco4957, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4958(w_eco4958, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4959(w_eco4959, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4960(w_eco4960, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4961(w_eco4961, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4962(w_eco4962, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4963(w_eco4963, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4964(w_eco4964, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4965(w_eco4965, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4966(w_eco4966, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4967(w_eco4967, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4968(w_eco4968, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4969(w_eco4969, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4970(w_eco4970, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4971(w_eco4971, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4972(w_eco4972, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4973(w_eco4973, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4974(w_eco4974, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4975(w_eco4975, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4976(w_eco4976, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4977(w_eco4977, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4978(w_eco4978, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4979(w_eco4979, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4980(w_eco4980, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4981(w_eco4981, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4982(w_eco4982, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4983(w_eco4983, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4984(w_eco4984, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4985(w_eco4985, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4986(w_eco4986, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4987(w_eco4987, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4988(w_eco4988, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4989(w_eco4989, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4990(w_eco4990, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4991(w_eco4991, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4992(w_eco4992, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4993(w_eco4993, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4994(w_eco4994, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_4995(w_eco4995, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_4996(w_eco4996, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4997(w_eco4997, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_4998(w_eco4998, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_4999(w_eco4999, Tsync[4], !Tsync[3], !prev_cnt[3], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5000(w_eco5000, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_5001(w_eco5001, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_5002(w_eco5002, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_5003(w_eco5003, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5004(w_eco5004, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5005(w_eco5005, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5006(w_eco5006, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5007(w_eco5007, !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5008(w_eco5008, !Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5009(w_eco5009, !Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5010(w_eco5010, !Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5011(w_eco5011, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5012(w_eco5012, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5013(w_eco5013, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5014(w_eco5014, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5015(w_eco5015, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5016(w_eco5016, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5017(w_eco5017, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5018(w_eco5018, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5019(w_eco5019, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5020(w_eco5020, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5021(w_eco5021, prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5022(w_eco5022, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5023(w_eco5023, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5024(w_eco5024, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5025(w_eco5025, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5026(w_eco5026, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5027(w_eco5027, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5028(w_eco5028, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5029(w_eco5029, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5030(w_eco5030, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5031(w_eco5031, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5032(w_eco5032, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5033(w_eco5033, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5034(w_eco5034, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5035(w_eco5035, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5036(w_eco5036, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5037(w_eco5037, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5038(w_eco5038, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5039(w_eco5039, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5040(w_eco5040, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5041(w_eco5041, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5042(w_eco5042, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5043(w_eco5043, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5044(w_eco5044, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5045(w_eco5045, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5046(w_eco5046, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5047(w_eco5047, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5048(w_eco5048, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5049(w_eco5049, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5050(w_eco5050, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5051(w_eco5051, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5052(w_eco5052, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5053(w_eco5053, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5054(w_eco5054, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5055(w_eco5055, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5056(w_eco5056, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5057(w_eco5057, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5058(w_eco5058, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5059(w_eco5059, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5060(w_eco5060, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5061(w_eco5061, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5062(w_eco5062, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5063(w_eco5063, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5064(w_eco5064, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5065(w_eco5065, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5066(w_eco5066, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5067(w_eco5067, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5068(w_eco5068, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5069(w_eco5069, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5070(w_eco5070, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5071(w_eco5071, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5072(w_eco5072, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5073(w_eco5073, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5074(w_eco5074, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5075(w_eco5075, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5076(w_eco5076, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5077(w_eco5077, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5078(w_eco5078, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5079(w_eco5079, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5080(w_eco5080, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5081(w_eco5081, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5082(w_eco5082, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5083(w_eco5083, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5084(w_eco5084, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5085(w_eco5085, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5086(w_eco5086, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5087(w_eco5087, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5088(w_eco5088, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5089(w_eco5089, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5090(w_eco5090, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5091(w_eco5091, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5092(w_eco5092, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5093(w_eco5093, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5094(w_eco5094, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5095(w_eco5095, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5096(w_eco5096, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5097(w_eco5097, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5098(w_eco5098, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5099(w_eco5099, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5100(w_eco5100, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5101(w_eco5101, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5102(w_eco5102, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5103(w_eco5103, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5104(w_eco5104, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5105(w_eco5105, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5106(w_eco5106, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5107(w_eco5107, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5108(w_eco5108, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5109(w_eco5109, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5110(w_eco5110, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5111(w_eco5111, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5112(w_eco5112, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5113(w_eco5113, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5114(w_eco5114, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5115(w_eco5115, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5116(w_eco5116, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5117(w_eco5117, Tsync[4], !Tsync[3], !prev_cnt[3], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5118(w_eco5118, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5119(w_eco5119, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5120(w_eco5120, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5121(w_eco5121, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5122(w_eco5122, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5123(w_eco5123, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5124(w_eco5124, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5125(w_eco5125, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5126(w_eco5126, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5127(w_eco5127, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5128(w_eco5128, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5129(w_eco5129, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5130(w_eco5130, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5131(w_eco5131, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5132(w_eco5132, !Tgate[4], !Tgdel[4], !Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5133(w_eco5133, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5134(w_eco5134, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5135(w_eco5135, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5136(w_eco5136, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5137(w_eco5137, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5138(w_eco5138, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5139(w_eco5139, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5140(w_eco5140, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5141(w_eco5141, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5142(w_eco5142, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5143(w_eco5143, prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5144(w_eco5144, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5145(w_eco5145, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5146(w_eco5146, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5147(w_eco5147, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5148(w_eco5148, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5149(w_eco5149, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5150(w_eco5150, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5151(w_eco5151, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5152(w_eco5152, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5153(w_eco5153, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5154(w_eco5154, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5155(w_eco5155, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5156(w_eco5156, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5157(w_eco5157, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5158(w_eco5158, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5159(w_eco5159, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5160(w_eco5160, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5161(w_eco5161, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5162(w_eco5162, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5163(w_eco5163, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5164(w_eco5164, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5165(w_eco5165, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5166(w_eco5166, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5167(w_eco5167, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5168(w_eco5168, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5169(w_eco5169, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5170(w_eco5170, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5171(w_eco5171, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5172(w_eco5172, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5173(w_eco5173, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5174(w_eco5174, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5175(w_eco5175, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5176(w_eco5176, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5177(w_eco5177, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5178(w_eco5178, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5179(w_eco5179, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5180(w_eco5180, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5181(w_eco5181, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5182(w_eco5182, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5183(w_eco5183, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5184(w_eco5184, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5185(w_eco5185, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5186(w_eco5186, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5187(w_eco5187, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5188(w_eco5188, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5189(w_eco5189, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5190(w_eco5190, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5191(w_eco5191, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5192(w_eco5192, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5193(w_eco5193, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5194(w_eco5194, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5195(w_eco5195, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5196(w_eco5196, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5197(w_eco5197, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5198(w_eco5198, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5199(w_eco5199, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5200(w_eco5200, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5201(w_eco5201, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5202(w_eco5202, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5203(w_eco5203, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5204(w_eco5204, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5205(w_eco5205, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5206(w_eco5206, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5207(w_eco5207, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5208(w_eco5208, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5209(w_eco5209, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5210(w_eco5210, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5211(w_eco5211, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5212(w_eco5212, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5213(w_eco5213, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5214(w_eco5214, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5215(w_eco5215, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5216(w_eco5216, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5217(w_eco5217, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5218(w_eco5218, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5219(w_eco5219, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5220(w_eco5220, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5221(w_eco5221, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5222(w_eco5222, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5223(w_eco5223, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5224(w_eco5224, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5225(w_eco5225, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5226(w_eco5226, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5227(w_eco5227, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5228(w_eco5228, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5229(w_eco5229, !Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5230(w_eco5230, !Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5231(w_eco5231, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5232(w_eco5232, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5233(w_eco5233, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5234(w_eco5234, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5235(w_eco5235, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5236(w_eco5236, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5237(w_eco5237, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5238(w_eco5238, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5239(w_eco5239, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5240(w_eco5240, prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5241(w_eco5241, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5242(w_eco5242, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5243(w_eco5243, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5244(w_eco5244, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5245(w_eco5245, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5246(w_eco5246, prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5247(w_eco5247, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5248(w_eco5248, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5249(w_eco5249, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5250(w_eco5250, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5251(w_eco5251, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5252(w_eco5252, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5253(w_eco5253, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5254(w_eco5254, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5255(w_eco5255, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5256(w_eco5256, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5257(w_eco5257, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5258(w_eco5258, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5259(w_eco5259, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5260(w_eco5260, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5261(w_eco5261, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5262(w_eco5262, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5263(w_eco5263, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5264(w_eco5264, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5265(w_eco5265, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5266(w_eco5266, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5267(w_eco5267, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5268(w_eco5268, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5269(w_eco5269, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5270(w_eco5270, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5271(w_eco5271, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5272(w_eco5272, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5273(w_eco5273, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5274(w_eco5274, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5275(w_eco5275, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5276(w_eco5276, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5277(w_eco5277, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5278(w_eco5278, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5279(w_eco5279, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5280(w_eco5280, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5281(w_eco5281, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5282(w_eco5282, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5283(w_eco5283, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5284(w_eco5284, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5285(w_eco5285, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5286(w_eco5286, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5287(w_eco5287, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5288(w_eco5288, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5289(w_eco5289, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5290(w_eco5290, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5291(w_eco5291, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5292(w_eco5292, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5293(w_eco5293, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5294(w_eco5294, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5295(w_eco5295, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5296(w_eco5296, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5297(w_eco5297, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5298(w_eco5298, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5299(w_eco5299, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5300(w_eco5300, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5301(w_eco5301, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5302(w_eco5302, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5303(w_eco5303, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5304(w_eco5304, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5305(w_eco5305, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5306(w_eco5306, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5307(w_eco5307, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5308(w_eco5308, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5309(w_eco5309, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5310(w_eco5310, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5311(w_eco5311, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5312(w_eco5312, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5313(w_eco5313, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5314(w_eco5314, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5315(w_eco5315, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5316(w_eco5316, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5317(w_eco5317, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5318(w_eco5318, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5319(w_eco5319, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5320(w_eco5320, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5321(w_eco5321, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5322(w_eco5322, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5323(w_eco5323, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5324(w_eco5324, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5325(w_eco5325, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5326(w_eco5326, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5327(w_eco5327, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5328(w_eco5328, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5329(w_eco5329, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5330(w_eco5330, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5331(w_eco5331, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5332(w_eco5332, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5333(w_eco5333, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5334(w_eco5334, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5335(w_eco5335, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5336(w_eco5336, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5337(w_eco5337, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5338(w_eco5338, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5339(w_eco5339, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5340(w_eco5340, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5341(w_eco5341, prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5342(w_eco5342, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5343(w_eco5343, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5344(w_eco5344, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5345(w_eco5345, prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5346(w_eco5346, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5347(w_eco5347, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5348(w_eco5348, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5349(w_eco5349, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5350(w_eco5350, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5351(w_eco5351, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5352(w_eco5352, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5353(w_eco5353, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5354(w_eco5354, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5355(w_eco5355, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5356(w_eco5356, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5357(w_eco5357, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5358(w_eco5358, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5359(w_eco5359, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5360(w_eco5360, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5361(w_eco5361, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5362(w_eco5362, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5363(w_eco5363, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5364(w_eco5364, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5365(w_eco5365, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5366(w_eco5366, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5367(w_eco5367, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5368(w_eco5368, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5369(w_eco5369, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5370(w_eco5370, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5371(w_eco5371, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5372(w_eco5372, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5373(w_eco5373, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5374(w_eco5374, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5375(w_eco5375, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5376(w_eco5376, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5377(w_eco5377, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5378(w_eco5378, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5379(w_eco5379, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5380(w_eco5380, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5381(w_eco5381, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5382(w_eco5382, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5383(w_eco5383, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5384(w_eco5384, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5385(w_eco5385, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5386(w_eco5386, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5387(w_eco5387, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5388(w_eco5388, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5389(w_eco5389, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5390(w_eco5390, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5391(w_eco5391, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5392(w_eco5392, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5393(w_eco5393, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5394(w_eco5394, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5395(w_eco5395, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5396(w_eco5396, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5397(w_eco5397, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5398(w_eco5398, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5399(w_eco5399, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5400(w_eco5400, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5401(w_eco5401, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5402(w_eco5402, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5403(w_eco5403, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5404(w_eco5404, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5405(w_eco5405, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5406(w_eco5406, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5407(w_eco5407, !Tgate[4], !Tsync[4], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5408(w_eco5408, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5409(w_eco5409, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5410(w_eco5410, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5411(w_eco5411, prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5412(w_eco5412, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5413(w_eco5413, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5414(w_eco5414, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5415(w_eco5415, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5416(w_eco5416, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5417(w_eco5417, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5418(w_eco5418, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5419(w_eco5419, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[4], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5420(w_eco5420, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5421(w_eco5421, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5422(w_eco5422, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5423(w_eco5423, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5424(w_eco5424, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5425(w_eco5425, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5426(w_eco5426, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5427(w_eco5427, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5428(w_eco5428, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5429(w_eco5429, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5430(w_eco5430, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5431(w_eco5431, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5432(w_eco5432, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5433(w_eco5433, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5434(w_eco5434, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5435(w_eco5435, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5436(w_eco5436, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5437(w_eco5437, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5438(w_eco5438, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5439(w_eco5439, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5440(w_eco5440, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5441(w_eco5441, Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5442(w_eco5442, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5443(w_eco5443, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5444(w_eco5444, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5445(w_eco5445, !Tgate[4], !Tgdel[4], Tsync[4], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5446(w_eco5446, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5447(w_eco5447, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5448(w_eco5448, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5449(w_eco5449, Tsync[4], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5450(w_eco5450, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5451(w_eco5451, !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5452(w_eco5452, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5453(w_eco5453, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5454(w_eco5454, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5455(w_eco5455, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5456(w_eco5456, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5457(w_eco5457, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5458(w_eco5458, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5459(w_eco5459, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5460(w_eco5460, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5461(w_eco5461, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5462(w_eco5462, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5463(w_eco5463, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5464(w_eco5464, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5465(w_eco5465, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5466(w_eco5466, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5467(w_eco5467, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5468(w_eco5468, !Tgate[4], !Tgdel[4], Tsync[4], Tsync[3], prev_cnt[3], !prev_cnt[4], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5469(w_eco5469, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5470(w_eco5470, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5471(w_eco5471, !Tgate[4], !Tsync[4], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5472(w_eco5472, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5473(w_eco5473, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5474(w_eco5474, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5475(w_eco5475, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5476(w_eco5476, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5477(w_eco5477, Tsync[4], !prev_cnt[14], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5478(w_eco5478, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5479(w_eco5479, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_5480(w_eco5480, w_eco3901, w_eco3902, w_eco3903, w_eco3904, w_eco3905, w_eco3906, w_eco3907, w_eco3908, w_eco3909, w_eco3910, w_eco3911, w_eco3912, w_eco3913, w_eco3914, w_eco3915, w_eco3916, w_eco3917, w_eco3918, w_eco3919, w_eco3920, w_eco3921, w_eco3922, w_eco3923, w_eco3924, w_eco3925, w_eco3926, w_eco3927, w_eco3928, w_eco3929, w_eco3930, w_eco3931, w_eco3932, w_eco3933, w_eco3934, w_eco3935, w_eco3936, w_eco3937, w_eco3938, w_eco3939, w_eco3940, w_eco3941, w_eco3942, w_eco3943, w_eco3944, w_eco3945, w_eco3946, w_eco3947, w_eco3948, w_eco3949, w_eco3950, w_eco3951, w_eco3952, w_eco3953, w_eco3954, w_eco3955, w_eco3956, w_eco3957, w_eco3958, w_eco3959, w_eco3960, w_eco3961, w_eco3962, w_eco3963, w_eco3964, w_eco3965, w_eco3966, w_eco3967, w_eco3968, w_eco3969, w_eco3970, w_eco3971, w_eco3972, w_eco3973, w_eco3974, w_eco3975, w_eco3976, w_eco3977, w_eco3978, w_eco3979, w_eco3980, w_eco3981, w_eco3982, w_eco3983, w_eco3984, w_eco3985, w_eco3986, w_eco3987, w_eco3988, w_eco3989, w_eco3990, w_eco3991, w_eco3992, w_eco3993, w_eco3994, w_eco3995, w_eco3996, w_eco3997, w_eco3998, w_eco3999, w_eco4000, w_eco4001, w_eco4002, w_eco4003, w_eco4004, w_eco4005, w_eco4006, w_eco4007, w_eco4008, w_eco4009, w_eco4010, w_eco4011, w_eco4012, w_eco4013, w_eco4014, w_eco4015, w_eco4016, w_eco4017, w_eco4018, w_eco4019, w_eco4020, w_eco4021, w_eco4022, w_eco4023, w_eco4024, w_eco4025, w_eco4026, w_eco4027, w_eco4028, w_eco4029, w_eco4030, w_eco4031, w_eco4032, w_eco4033, w_eco4034, w_eco4035, w_eco4036, w_eco4037, w_eco4038, w_eco4039, w_eco4040, w_eco4041, w_eco4042, w_eco4043, w_eco4044, w_eco4045, w_eco4046, w_eco4047, w_eco4048, w_eco4049, w_eco4050, w_eco4051, w_eco4052, w_eco4053, w_eco4054, w_eco4055, w_eco4056, w_eco4057, w_eco4058, w_eco4059, w_eco4060, w_eco4061, w_eco4062, w_eco4063, w_eco4064, w_eco4065, w_eco4066, w_eco4067, w_eco4068, w_eco4069, w_eco4070, w_eco4071, w_eco4072, w_eco4073, w_eco4074, w_eco4075, w_eco4076, w_eco4077, w_eco4078, w_eco4079, w_eco4080, w_eco4081, w_eco4082, w_eco4083, w_eco4084, w_eco4085, w_eco4086, w_eco4087, w_eco4088, w_eco4089, w_eco4090, w_eco4091, w_eco4092, w_eco4093, w_eco4094, w_eco4095, w_eco4096, w_eco4097, w_eco4098, w_eco4099, w_eco4100, w_eco4101, w_eco4102, w_eco4103, w_eco4104, w_eco4105, w_eco4106, w_eco4107, w_eco4108, w_eco4109, w_eco4110, w_eco4111, w_eco4112, w_eco4113, w_eco4114, w_eco4115, w_eco4116, w_eco4117, w_eco4118, w_eco4119, w_eco4120, w_eco4121, w_eco4122, w_eco4123, w_eco4124, w_eco4125, w_eco4126, w_eco4127, w_eco4128, w_eco4129, w_eco4130, w_eco4131, w_eco4132, w_eco4133, w_eco4134, w_eco4135, w_eco4136, w_eco4137, w_eco4138, w_eco4139, w_eco4140, w_eco4141, w_eco4142, w_eco4143, w_eco4144, w_eco4145, w_eco4146, w_eco4147, w_eco4148, w_eco4149, w_eco4150, w_eco4151, w_eco4152, w_eco4153, w_eco4154, w_eco4155, w_eco4156, w_eco4157, w_eco4158, w_eco4159, w_eco4160, w_eco4161, w_eco4162, w_eco4163, w_eco4164, w_eco4165, w_eco4166, w_eco4167, w_eco4168, w_eco4169, w_eco4170, w_eco4171, w_eco4172, w_eco4173, w_eco4174, w_eco4175, w_eco4176, w_eco4177, w_eco4178, w_eco4179, w_eco4180, w_eco4181, w_eco4182, w_eco4183, w_eco4184, w_eco4185, w_eco4186, w_eco4187, w_eco4188, w_eco4189, w_eco4190, w_eco4191, w_eco4192, w_eco4193, w_eco4194, w_eco4195, w_eco4196, w_eco4197, w_eco4198, w_eco4199, w_eco4200, w_eco4201, w_eco4202, w_eco4203, w_eco4204, w_eco4205, w_eco4206, w_eco4207, w_eco4208, w_eco4209, w_eco4210, w_eco4211, w_eco4212, w_eco4213, w_eco4214, w_eco4215, w_eco4216, w_eco4217, w_eco4218, w_eco4219, w_eco4220, w_eco4221, w_eco4222, w_eco4223, w_eco4224, w_eco4225, w_eco4226, w_eco4227, w_eco4228, w_eco4229, w_eco4230, w_eco4231, w_eco4232, w_eco4233, w_eco4234, w_eco4235, w_eco4236, w_eco4237, w_eco4238, w_eco4239, w_eco4240, w_eco4241, w_eco4242, w_eco4243, w_eco4244, w_eco4245, w_eco4246, w_eco4247, w_eco4248, w_eco4249, w_eco4250, w_eco4251, w_eco4252, w_eco4253, w_eco4254, w_eco4255, w_eco4256, w_eco4257, w_eco4258, w_eco4259, w_eco4260, w_eco4261, w_eco4262, w_eco4263, w_eco4264, w_eco4265, w_eco4266, w_eco4267, w_eco4268, w_eco4269, w_eco4270, w_eco4271, w_eco4272, w_eco4273, w_eco4274, w_eco4275, w_eco4276, w_eco4277, w_eco4278, w_eco4279, w_eco4280, w_eco4281, w_eco4282, w_eco4283, w_eco4284, w_eco4285, w_eco4286, w_eco4287, w_eco4288, w_eco4289, w_eco4290, w_eco4291, w_eco4292, w_eco4293, w_eco4294, w_eco4295, w_eco4296, w_eco4297, w_eco4298, w_eco4299, w_eco4300, w_eco4301, w_eco4302, w_eco4303, w_eco4304, w_eco4305, w_eco4306, w_eco4307, w_eco4308, w_eco4309, w_eco4310, w_eco4311, w_eco4312, w_eco4313, w_eco4314, w_eco4315, w_eco4316, w_eco4317, w_eco4318, w_eco4319, w_eco4320, w_eco4321, w_eco4322, w_eco4323, w_eco4324, w_eco4325, w_eco4326, w_eco4327, w_eco4328, w_eco4329, w_eco4330, w_eco4331, w_eco4332, w_eco4333, w_eco4334, w_eco4335, w_eco4336, w_eco4337, w_eco4338, w_eco4339, w_eco4340, w_eco4341, w_eco4342, w_eco4343, w_eco4344, w_eco4345, w_eco4346, w_eco4347, w_eco4348, w_eco4349, w_eco4350, w_eco4351, w_eco4352, w_eco4353, w_eco4354, w_eco4355, w_eco4356, w_eco4357, w_eco4358, w_eco4359, w_eco4360, w_eco4361, w_eco4362, w_eco4363, w_eco4364, w_eco4365, w_eco4366, w_eco4367, w_eco4368, w_eco4369, w_eco4370, w_eco4371, w_eco4372, w_eco4373, w_eco4374, w_eco4375, w_eco4376, w_eco4377, w_eco4378, w_eco4379, w_eco4380, w_eco4381, w_eco4382, w_eco4383, w_eco4384, w_eco4385, w_eco4386, w_eco4387, w_eco4388, w_eco4389, w_eco4390, w_eco4391, w_eco4392, w_eco4393, w_eco4394, w_eco4395, w_eco4396, w_eco4397, w_eco4398, w_eco4399, w_eco4400, w_eco4401, w_eco4402, w_eco4403, w_eco4404, w_eco4405, w_eco4406, w_eco4407, w_eco4408, w_eco4409, w_eco4410, w_eco4411, w_eco4412, w_eco4413, w_eco4414, w_eco4415, w_eco4416, w_eco4417, w_eco4418, w_eco4419, w_eco4420, w_eco4421, w_eco4422, w_eco4423, w_eco4424, w_eco4425, w_eco4426, w_eco4427, w_eco4428, w_eco4429, w_eco4430, w_eco4431, w_eco4432, w_eco4433, w_eco4434, w_eco4435, w_eco4436, w_eco4437, w_eco4438, w_eco4439, w_eco4440, w_eco4441, w_eco4442, w_eco4443, w_eco4444, w_eco4445, w_eco4446, w_eco4447, w_eco4448, w_eco4449, w_eco4450, w_eco4451, w_eco4452, w_eco4453, w_eco4454, w_eco4455, w_eco4456, w_eco4457, w_eco4458, w_eco4459, w_eco4460, w_eco4461, w_eco4462, w_eco4463, w_eco4464, w_eco4465, w_eco4466, w_eco4467, w_eco4468, w_eco4469, w_eco4470, w_eco4471, w_eco4472, w_eco4473, w_eco4474, w_eco4475, w_eco4476, w_eco4477, w_eco4478, w_eco4479, w_eco4480, w_eco4481, w_eco4482, w_eco4483, w_eco4484, w_eco4485, w_eco4486, w_eco4487, w_eco4488, w_eco4489, w_eco4490, w_eco4491, w_eco4492, w_eco4493, w_eco4494, w_eco4495, w_eco4496, w_eco4497, w_eco4498, w_eco4499, w_eco4500, w_eco4501, w_eco4502, w_eco4503, w_eco4504, w_eco4505, w_eco4506, w_eco4507, w_eco4508, w_eco4509, w_eco4510, w_eco4511, w_eco4512, w_eco4513, w_eco4514, w_eco4515, w_eco4516, w_eco4517, w_eco4518, w_eco4519, w_eco4520, w_eco4521, w_eco4522, w_eco4523, w_eco4524, w_eco4525, w_eco4526, w_eco4527, w_eco4528, w_eco4529, w_eco4530, w_eco4531, w_eco4532, w_eco4533, w_eco4534, w_eco4535, w_eco4536, w_eco4537, w_eco4538, w_eco4539, w_eco4540, w_eco4541, w_eco4542, w_eco4543, w_eco4544, w_eco4545, w_eco4546, w_eco4547, w_eco4548, w_eco4549, w_eco4550, w_eco4551, w_eco4552, w_eco4553, w_eco4554, w_eco4555, w_eco4556, w_eco4557, w_eco4558, w_eco4559, w_eco4560, w_eco4561, w_eco4562, w_eco4563, w_eco4564, w_eco4565, w_eco4566, w_eco4567, w_eco4568, w_eco4569, w_eco4570, w_eco4571, w_eco4572, w_eco4573, w_eco4574, w_eco4575, w_eco4576, w_eco4577, w_eco4578, w_eco4579, w_eco4580, w_eco4581, w_eco4582, w_eco4583, w_eco4584, w_eco4585, w_eco4586, w_eco4587, w_eco4588, w_eco4589, w_eco4590, w_eco4591, w_eco4592, w_eco4593, w_eco4594, w_eco4595, w_eco4596, w_eco4597, w_eco4598, w_eco4599, w_eco4600, w_eco4601, w_eco4602, w_eco4603, w_eco4604, w_eco4605, w_eco4606, w_eco4607, w_eco4608, w_eco4609, w_eco4610, w_eco4611, w_eco4612, w_eco4613, w_eco4614, w_eco4615, w_eco4616, w_eco4617, w_eco4618, w_eco4619, w_eco4620, w_eco4621, w_eco4622, w_eco4623, w_eco4624, w_eco4625, w_eco4626, w_eco4627, w_eco4628, w_eco4629, w_eco4630, w_eco4631, w_eco4632, w_eco4633, w_eco4634, w_eco4635, w_eco4636, w_eco4637, w_eco4638, w_eco4639, w_eco4640, w_eco4641, w_eco4642, w_eco4643, w_eco4644, w_eco4645, w_eco4646, w_eco4647, w_eco4648, w_eco4649, w_eco4650, w_eco4651, w_eco4652, w_eco4653, w_eco4654, w_eco4655, w_eco4656, w_eco4657, w_eco4658, w_eco4659, w_eco4660, w_eco4661, w_eco4662, w_eco4663, w_eco4664, w_eco4665, w_eco4666, w_eco4667, w_eco4668, w_eco4669, w_eco4670, w_eco4671, w_eco4672, w_eco4673, w_eco4674, w_eco4675, w_eco4676, w_eco4677, w_eco4678, w_eco4679, w_eco4680, w_eco4681, w_eco4682, w_eco4683, w_eco4684, w_eco4685, w_eco4686, w_eco4687, w_eco4688, w_eco4689, w_eco4690, w_eco4691, w_eco4692, w_eco4693, w_eco4694, w_eco4695, w_eco4696, w_eco4697, w_eco4698, w_eco4699, w_eco4700, w_eco4701, w_eco4702, w_eco4703, w_eco4704, w_eco4705, w_eco4706, w_eco4707, w_eco4708, w_eco4709, w_eco4710, w_eco4711, w_eco4712, w_eco4713, w_eco4714, w_eco4715, w_eco4716, w_eco4717, w_eco4718, w_eco4719, w_eco4720, w_eco4721, w_eco4722, w_eco4723, w_eco4724, w_eco4725, w_eco4726, w_eco4727, w_eco4728, w_eco4729, w_eco4730, w_eco4731, w_eco4732, w_eco4733, w_eco4734, w_eco4735, w_eco4736, w_eco4737, w_eco4738, w_eco4739, w_eco4740, w_eco4741, w_eco4742, w_eco4743, w_eco4744, w_eco4745, w_eco4746, w_eco4747, w_eco4748, w_eco4749, w_eco4750, w_eco4751, w_eco4752, w_eco4753, w_eco4754, w_eco4755, w_eco4756, w_eco4757, w_eco4758, w_eco4759, w_eco4760, w_eco4761, w_eco4762, w_eco4763, w_eco4764, w_eco4765, w_eco4766, w_eco4767, w_eco4768, w_eco4769, w_eco4770, w_eco4771, w_eco4772, w_eco4773, w_eco4774, w_eco4775, w_eco4776, w_eco4777, w_eco4778, w_eco4779, w_eco4780, w_eco4781, w_eco4782, w_eco4783, w_eco4784, w_eco4785, w_eco4786, w_eco4787, w_eco4788, w_eco4789, w_eco4790, w_eco4791, w_eco4792, w_eco4793, w_eco4794, w_eco4795, w_eco4796, w_eco4797, w_eco4798, w_eco4799, w_eco4800, w_eco4801, w_eco4802, w_eco4803, w_eco4804, w_eco4805, w_eco4806, w_eco4807, w_eco4808, w_eco4809, w_eco4810, w_eco4811, w_eco4812, w_eco4813, w_eco4814, w_eco4815, w_eco4816, w_eco4817, w_eco4818, w_eco4819, w_eco4820, w_eco4821, w_eco4822, w_eco4823, w_eco4824, w_eco4825, w_eco4826, w_eco4827, w_eco4828, w_eco4829, w_eco4830, w_eco4831, w_eco4832, w_eco4833, w_eco4834, w_eco4835, w_eco4836, w_eco4837, w_eco4838, w_eco4839, w_eco4840, w_eco4841, w_eco4842, w_eco4843, w_eco4844, w_eco4845, w_eco4846, w_eco4847, w_eco4848, w_eco4849, w_eco4850, w_eco4851, w_eco4852, w_eco4853, w_eco4854, w_eco4855, w_eco4856, w_eco4857, w_eco4858, w_eco4859, w_eco4860, w_eco4861, w_eco4862, w_eco4863, w_eco4864, w_eco4865, w_eco4866, w_eco4867, w_eco4868, w_eco4869, w_eco4870, w_eco4871, w_eco4872, w_eco4873, w_eco4874, w_eco4875, w_eco4876, w_eco4877, w_eco4878, w_eco4879, w_eco4880, w_eco4881, w_eco4882, w_eco4883, w_eco4884, w_eco4885, w_eco4886, w_eco4887, w_eco4888, w_eco4889, w_eco4890, w_eco4891, w_eco4892, w_eco4893, w_eco4894, w_eco4895, w_eco4896, w_eco4897, w_eco4898, w_eco4899, w_eco4900, w_eco4901, w_eco4902, w_eco4903, w_eco4904, w_eco4905, w_eco4906, w_eco4907, w_eco4908, w_eco4909, w_eco4910, w_eco4911, w_eco4912, w_eco4913, w_eco4914, w_eco4915, w_eco4916, w_eco4917, w_eco4918, w_eco4919, w_eco4920, w_eco4921, w_eco4922, w_eco4923, w_eco4924, w_eco4925, w_eco4926, w_eco4927, w_eco4928, w_eco4929, w_eco4930, w_eco4931, w_eco4932, w_eco4933, w_eco4934, w_eco4935, w_eco4936, w_eco4937, w_eco4938, w_eco4939, w_eco4940, w_eco4941, w_eco4942, w_eco4943, w_eco4944, w_eco4945, w_eco4946, w_eco4947, w_eco4948, w_eco4949, w_eco4950, w_eco4951, w_eco4952, w_eco4953, w_eco4954, w_eco4955, w_eco4956, w_eco4957, w_eco4958, w_eco4959, w_eco4960, w_eco4961, w_eco4962, w_eco4963, w_eco4964, w_eco4965, w_eco4966, w_eco4967, w_eco4968, w_eco4969, w_eco4970, w_eco4971, w_eco4972, w_eco4973, w_eco4974, w_eco4975, w_eco4976, w_eco4977, w_eco4978, w_eco4979, w_eco4980, w_eco4981, w_eco4982, w_eco4983, w_eco4984, w_eco4985, w_eco4986, w_eco4987, w_eco4988, w_eco4989, w_eco4990, w_eco4991, w_eco4992, w_eco4993, w_eco4994, w_eco4995, w_eco4996, w_eco4997, w_eco4998, w_eco4999, w_eco5000, w_eco5001, w_eco5002, w_eco5003, w_eco5004, w_eco5005, w_eco5006, w_eco5007, w_eco5008, w_eco5009, w_eco5010, w_eco5011, w_eco5012, w_eco5013, w_eco5014, w_eco5015, w_eco5016, w_eco5017, w_eco5018, w_eco5019, w_eco5020, w_eco5021, w_eco5022, w_eco5023, w_eco5024, w_eco5025, w_eco5026, w_eco5027, w_eco5028, w_eco5029, w_eco5030, w_eco5031, w_eco5032, w_eco5033, w_eco5034, w_eco5035, w_eco5036, w_eco5037, w_eco5038, w_eco5039, w_eco5040, w_eco5041, w_eco5042, w_eco5043, w_eco5044, w_eco5045, w_eco5046, w_eco5047, w_eco5048, w_eco5049, w_eco5050, w_eco5051, w_eco5052, w_eco5053, w_eco5054, w_eco5055, w_eco5056, w_eco5057, w_eco5058, w_eco5059, w_eco5060, w_eco5061, w_eco5062, w_eco5063, w_eco5064, w_eco5065, w_eco5066, w_eco5067, w_eco5068, w_eco5069, w_eco5070, w_eco5071, w_eco5072, w_eco5073, w_eco5074, w_eco5075, w_eco5076, w_eco5077, w_eco5078, w_eco5079, w_eco5080, w_eco5081, w_eco5082, w_eco5083, w_eco5084, w_eco5085, w_eco5086, w_eco5087, w_eco5088, w_eco5089, w_eco5090, w_eco5091, w_eco5092, w_eco5093, w_eco5094, w_eco5095, w_eco5096, w_eco5097, w_eco5098, w_eco5099, w_eco5100, w_eco5101, w_eco5102, w_eco5103, w_eco5104, w_eco5105, w_eco5106, w_eco5107, w_eco5108, w_eco5109, w_eco5110, w_eco5111, w_eco5112, w_eco5113, w_eco5114, w_eco5115, w_eco5116, w_eco5117, w_eco5118, w_eco5119, w_eco5120, w_eco5121, w_eco5122, w_eco5123, w_eco5124, w_eco5125, w_eco5126, w_eco5127, w_eco5128, w_eco5129, w_eco5130, w_eco5131, w_eco5132, w_eco5133, w_eco5134, w_eco5135, w_eco5136, w_eco5137, w_eco5138, w_eco5139, w_eco5140, w_eco5141, w_eco5142, w_eco5143, w_eco5144, w_eco5145, w_eco5146, w_eco5147, w_eco5148, w_eco5149, w_eco5150, w_eco5151, w_eco5152, w_eco5153, w_eco5154, w_eco5155, w_eco5156, w_eco5157, w_eco5158, w_eco5159, w_eco5160, w_eco5161, w_eco5162, w_eco5163, w_eco5164, w_eco5165, w_eco5166, w_eco5167, w_eco5168, w_eco5169, w_eco5170, w_eco5171, w_eco5172, w_eco5173, w_eco5174, w_eco5175, w_eco5176, w_eco5177, w_eco5178, w_eco5179, w_eco5180, w_eco5181, w_eco5182, w_eco5183, w_eco5184, w_eco5185, w_eco5186, w_eco5187, w_eco5188, w_eco5189, w_eco5190, w_eco5191, w_eco5192, w_eco5193, w_eco5194, w_eco5195, w_eco5196, w_eco5197, w_eco5198, w_eco5199, w_eco5200, w_eco5201, w_eco5202, w_eco5203, w_eco5204, w_eco5205, w_eco5206, w_eco5207, w_eco5208, w_eco5209, w_eco5210, w_eco5211, w_eco5212, w_eco5213, w_eco5214, w_eco5215, w_eco5216, w_eco5217, w_eco5218, w_eco5219, w_eco5220, w_eco5221, w_eco5222, w_eco5223, w_eco5224, w_eco5225, w_eco5226, w_eco5227, w_eco5228, w_eco5229, w_eco5230, w_eco5231, w_eco5232, w_eco5233, w_eco5234, w_eco5235, w_eco5236, w_eco5237, w_eco5238, w_eco5239, w_eco5240, w_eco5241, w_eco5242, w_eco5243, w_eco5244, w_eco5245, w_eco5246, w_eco5247, w_eco5248, w_eco5249, w_eco5250, w_eco5251, w_eco5252, w_eco5253, w_eco5254, w_eco5255, w_eco5256, w_eco5257, w_eco5258, w_eco5259, w_eco5260, w_eco5261, w_eco5262, w_eco5263, w_eco5264, w_eco5265, w_eco5266, w_eco5267, w_eco5268, w_eco5269, w_eco5270, w_eco5271, w_eco5272, w_eco5273, w_eco5274, w_eco5275, w_eco5276, w_eco5277, w_eco5278, w_eco5279, w_eco5280, w_eco5281, w_eco5282, w_eco5283, w_eco5284, w_eco5285, w_eco5286, w_eco5287, w_eco5288, w_eco5289, w_eco5290, w_eco5291, w_eco5292, w_eco5293, w_eco5294, w_eco5295, w_eco5296, w_eco5297, w_eco5298, w_eco5299, w_eco5300, w_eco5301, w_eco5302, w_eco5303, w_eco5304, w_eco5305, w_eco5306, w_eco5307, w_eco5308, w_eco5309, w_eco5310, w_eco5311, w_eco5312, w_eco5313, w_eco5314, w_eco5315, w_eco5316, w_eco5317, w_eco5318, w_eco5319, w_eco5320, w_eco5321, w_eco5322, w_eco5323, w_eco5324, w_eco5325, w_eco5326, w_eco5327, w_eco5328, w_eco5329, w_eco5330, w_eco5331, w_eco5332, w_eco5333, w_eco5334, w_eco5335, w_eco5336, w_eco5337, w_eco5338, w_eco5339, w_eco5340, w_eco5341, w_eco5342, w_eco5343, w_eco5344, w_eco5345, w_eco5346, w_eco5347, w_eco5348, w_eco5349, w_eco5350, w_eco5351, w_eco5352, w_eco5353, w_eco5354, w_eco5355, w_eco5356, w_eco5357, w_eco5358, w_eco5359, w_eco5360, w_eco5361, w_eco5362, w_eco5363, w_eco5364, w_eco5365, w_eco5366, w_eco5367, w_eco5368, w_eco5369, w_eco5370, w_eco5371, w_eco5372, w_eco5373, w_eco5374, w_eco5375, w_eco5376, w_eco5377, w_eco5378, w_eco5379, w_eco5380, w_eco5381, w_eco5382, w_eco5383, w_eco5384, w_eco5385, w_eco5386, w_eco5387, w_eco5388, w_eco5389, w_eco5390, w_eco5391, w_eco5392, w_eco5393, w_eco5394, w_eco5395, w_eco5396, w_eco5397, w_eco5398, w_eco5399, w_eco5400, w_eco5401, w_eco5402, w_eco5403, w_eco5404, w_eco5405, w_eco5406, w_eco5407, w_eco5408, w_eco5409, w_eco5410, w_eco5411, w_eco5412, w_eco5413, w_eco5414, w_eco5415, w_eco5416, w_eco5417, w_eco5418, w_eco5419, w_eco5420, w_eco5421, w_eco5422, w_eco5423, w_eco5424, w_eco5425, w_eco5426, w_eco5427, w_eco5428, w_eco5429, w_eco5430, w_eco5431, w_eco5432, w_eco5433, w_eco5434, w_eco5435, w_eco5436, w_eco5437, w_eco5438, w_eco5439, w_eco5440, w_eco5441, w_eco5442, w_eco5443, w_eco5444, w_eco5445, w_eco5446, w_eco5447, w_eco5448, w_eco5449, w_eco5450, w_eco5451, w_eco5452, w_eco5453, w_eco5454, w_eco5455, w_eco5456, w_eco5457, w_eco5458, w_eco5459, w_eco5460, w_eco5461, w_eco5462, w_eco5463, w_eco5464, w_eco5465, w_eco5466, w_eco5467, w_eco5468, w_eco5469, w_eco5470, w_eco5471, w_eco5472, w_eco5473, w_eco5474, w_eco5475, w_eco5476, w_eco5477, w_eco5478, w_eco5479);
	xor _ECO_out4(cnt[4], sub_wire4, w_eco5480);
	assign w_eco5481 = rst;
	and _ECO_5482(w_eco5482, Tgate[3], prev_cnt[1], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5483(w_eco5483, Tgate[3], prev_cnt[1], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5484(w_eco5484, Tgate[3], prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1]);
	and _ECO_5485(w_eco5485, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5486(w_eco5486, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], !ena);
	and _ECO_5487(w_eco5487, prev_cnt[1], prev_cnt[3], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5488(w_eco5488, Tgate[3], prev_cnt[2], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5489(w_eco5489, Tgate[3], prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_5490(w_eco5490, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5491(w_eco5491, !Tsync[4], prev_cnt[1], prev_cnt[3], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5492(w_eco5492, Tsync[3], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5493(w_eco5493, prev_cnt[1], prev_cnt[3], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5494(w_eco5494, Tgate[3], prev_cnt[2], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5495(w_eco5495, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5496(w_eco5496, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_5497(w_eco5497, Tgate[3], prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1]);
	and _ECO_5498(w_eco5498, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5499(w_eco5499, Tsync[3], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5500(w_eco5500, !Tsync[4], prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[0]);
	and _ECO_5501(w_eco5501, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_5502(w_eco5502, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], !ena);
	and _ECO_5503(w_eco5503, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], !ena);
	and _ECO_5504(w_eco5504, Tgate[3], prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_5505(w_eco5505, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5506(w_eco5506, !Tsync[4], prev_cnt[2], prev_cnt[3], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5507(w_eco5507, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5508(w_eco5508, !Tsync[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5509(w_eco5509, Tsync[3], !prev_cnt[4], ena, !prev_state[0]);
	and _ECO_5510(w_eco5510, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_5511(w_eco5511, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_5512(w_eco5512, !Tsync[4], prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[0]);
	and _ECO_5513(w_eco5513, !Tgate[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5514(w_eco5514, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], !ena);
	and _ECO_5515(w_eco5515, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], !ena);
	and _ECO_5516(w_eco5516, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], !ena);
	and _ECO_5517(w_eco5517, prev_cnt[1], prev_cnt[3], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5518(w_eco5518, prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5519(w_eco5519, Tgate[3], prev_cnt[0], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5520(w_eco5520, Tgate[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5521(w_eco5521, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[1]);
	and _ECO_5522(w_eco5522, !Tsync[4], Tsync[3], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_5523(w_eco5523, !Tsync[4], Tgate[3], prev_cnt[1], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5524(w_eco5524, !Tsync[4], prev_cnt[1], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5525(w_eco5525, prev_cnt[1], prev_cnt[3], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5526(w_eco5526, prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5527(w_eco5527, Tgate[3], prev_cnt[0], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5528(w_eco5528, Tgate[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5529(w_eco5529, !Tsync[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5530(w_eco5530, Tsync[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1]);
	and _ECO_5531(w_eco5531, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5532(w_eco5532, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[1]);
	and _ECO_5533(w_eco5533, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[1]);
	and _ECO_5534(w_eco5534, Tgate[3], prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1]);
	and _ECO_5535(w_eco5535, Tgate[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1]);
	and _ECO_5536(w_eco5536, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5537(w_eco5537, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5538(w_eco5538, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5539(w_eco5539, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5540(w_eco5540, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_state[1]);
	and _ECO_5541(w_eco5541, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_5542(w_eco5542, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], !ena);
	and _ECO_5543(w_eco5543, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], !ena);
	and _ECO_5544(w_eco5544, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], !ena);
	and _ECO_5545(w_eco5545, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5546(w_eco5546, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5547(w_eco5547, !Tsync[4], Tgate[3], prev_cnt[0], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5548(w_eco5548, !Tsync[4], Tgate[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5549(w_eco5549, !Tsync[4], prev_cnt[0], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5550(w_eco5550, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5551(w_eco5551, prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5552(w_eco5552, prev_cnt[0], prev_cnt[3], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5553(w_eco5553, Tgate[3], prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_5554(w_eco5554, Tgate[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0]);
	and _ECO_5555(w_eco5555, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5556(w_eco5556, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5557(w_eco5557, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5558(w_eco5558, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5559(w_eco5559, !Tsync[4], prev_cnt[0], prev_cnt[3], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5560(w_eco5560, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5561(w_eco5561, prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5562(w_eco5562, prev_cnt[0], prev_cnt[3], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5563(w_eco5563, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5564(w_eco5564, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5565(w_eco5565, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_5566(w_eco5566, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_5567(w_eco5567, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_5568(w_eco5568, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_state[3], !prev_state[2]);
	and _ECO_5569(w_eco5569, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_5570(w_eco5570, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_5571(w_eco5571, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5572(w_eco5572, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[1]);
	and _ECO_5573(w_eco5573, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[1]);
	and _ECO_5574(w_eco5574, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], prev_state[1]);
	and _ECO_5575(w_eco5575, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_5576(w_eco5576, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_state[4], !prev_state[2]);
	and _ECO_5577(w_eco5577, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5578(w_eco5578, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5579(w_eco5579, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5580(w_eco5580, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5581(w_eco5581, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5582(w_eco5582, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5583(w_eco5583, !Tsync[4], prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[0]);
	and _ECO_5584(w_eco5584, !Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[0]);
	and _ECO_5585(w_eco5585, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_5586(w_eco5586, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_5587(w_eco5587, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], !ena);
	and _ECO_5588(w_eco5588, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], !ena);
	and _ECO_5589(w_eco5589, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5590(w_eco5590, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5591(w_eco5591, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5592(w_eco5592, Tgdel[3], prev_cnt[1], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5593(w_eco5593, prev_cnt[0], prev_cnt[3], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5594(w_eco5594, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5595(w_eco5595, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5596(w_eco5596, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5597(w_eco5597, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5598(w_eco5598, !Tsync[4], Tgate[3], prev_cnt[2], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5599(w_eco5599, !Tsync[4], prev_cnt[2], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5600(w_eco5600, Tgdel[3], prev_cnt[1], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5601(w_eco5601, prev_cnt[0], prev_cnt[3], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5602(w_eco5602, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5603(w_eco5603, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_5604(w_eco5604, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_5605(w_eco5605, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_5606(w_eco5606, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_5607(w_eco5607, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_5608(w_eco5608, !Tsync[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5609(w_eco5609, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5610(w_eco5610, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5611(w_eco5611, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[1]);
	and _ECO_5612(w_eco5612, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[1]);
	and _ECO_5613(w_eco5613, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], prev_state[1]);
	and _ECO_5614(w_eco5614, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_5615(w_eco5615, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_5616(w_eco5616, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5617(w_eco5617, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5618(w_eco5618, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5619(w_eco5619, !Tgate[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5620(w_eco5620, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], !ena);
	and _ECO_5621(w_eco5621, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], !ena);
	and _ECO_5622(w_eco5622, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], !ena);
	and _ECO_5623(w_eco5623, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], !ena);
	and _ECO_5624(w_eco5624, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5625(w_eco5625, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5626(w_eco5626, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5627(w_eco5627, prev_cnt[1], prev_cnt[3], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5628(w_eco5628, Tgdel[3], prev_cnt[2], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5629(w_eco5629, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5630(w_eco5630, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5631(w_eco5631, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5632(w_eco5632, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5633(w_eco5633, prev_cnt[1], prev_cnt[3], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5634(w_eco5634, Tgdel[3], prev_cnt[2], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5635(w_eco5635, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5636(w_eco5636, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_5637(w_eco5637, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_5638(w_eco5638, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_5639(w_eco5639, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_5640(w_eco5640, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_5641(w_eco5641, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_5642(w_eco5642, !Tsync[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5643(w_eco5643, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5644(w_eco5644, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5645(w_eco5645, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5646(w_eco5646, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[1]);
	and _ECO_5647(w_eco5647, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[1]);
	and _ECO_5648(w_eco5648, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_5649(w_eco5649, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_5650(w_eco5650, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_5651(w_eco5651, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5652(w_eco5652, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5653(w_eco5653, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5654(w_eco5654, !Tgate[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5655(w_eco5655, !Tgate[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_5656(w_eco5656, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5657(w_eco5657, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], !ena);
	and _ECO_5658(w_eco5658, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], !ena);
	and _ECO_5659(w_eco5659, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], !ena);
	and _ECO_5660(w_eco5660, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], !ena);
	and _ECO_5661(w_eco5661, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5662(w_eco5662, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5663(w_eco5663, prev_cnt[1], prev_cnt[3], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5664(w_eco5664, prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5665(w_eco5665, Tgdel[3], prev_cnt[0], prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5666(w_eco5666, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5667(w_eco5667, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5668(w_eco5668, prev_cnt[14], prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5669(w_eco5669, prev_cnt[1], prev_cnt[3], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5670(w_eco5670, prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5671(w_eco5671, Tgdel[3], prev_cnt[0], prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5672(w_eco5672, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_5673(w_eco5673, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_5674(w_eco5674, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_5675(w_eco5675, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_5676(w_eco5676, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_5677(w_eco5677, !Tsync[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5678(w_eco5678, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5679(w_eco5679, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5680(w_eco5680, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5681(w_eco5681, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[1]);
	and _ECO_5682(w_eco5682, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[1]);
	and _ECO_5683(w_eco5683, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[1]);
	and _ECO_5684(w_eco5684, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], prev_state[1]);
	and _ECO_5685(w_eco5685, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_5686(w_eco5686, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_5687(w_eco5687, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_5688(w_eco5688, prev_cnt[14], prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5689(w_eco5689, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5690(w_eco5690, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5691(w_eco5691, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_5692(w_eco5692, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5693(w_eco5693, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], !ena);
	and _ECO_5694(w_eco5694, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], !ena);
	and _ECO_5695(w_eco5695, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], !ena);
	and _ECO_5696(w_eco5696, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], !ena);
	and _ECO_5697(w_eco5697, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], !ena);
	and _ECO_5698(w_eco5698, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5699(w_eco5699, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5700(w_eco5700, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5701(w_eco5701, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5702(w_eco5702, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5703(w_eco5703, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5704(w_eco5704, Tgate[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5705(w_eco5705, prev_cnt[1], prev_cnt[3], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5706(w_eco5706, prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5707(w_eco5707, prev_cnt[0], prev_cnt[3], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5708(w_eco5708, Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5709(w_eco5709, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5710(w_eco5710, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5711(w_eco5711, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5712(w_eco5712, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5713(w_eco5713, Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5714(w_eco5714, prev_cnt[14], prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5715(w_eco5715, Tgate[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5716(w_eco5716, prev_cnt[1], prev_cnt[3], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5717(w_eco5717, prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5718(w_eco5718, prev_cnt[0], prev_cnt[3], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5719(w_eco5719, Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5720(w_eco5720, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_5721(w_eco5721, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_5722(w_eco5722, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_5723(w_eco5723, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_5724(w_eco5724, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_5725(w_eco5725, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_5726(w_eco5726, !Tsync[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5727(w_eco5727, prev_cnt[14], prev_cnt[1], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5728(w_eco5728, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5729(w_eco5729, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5730(w_eco5730, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[1]);
	and _ECO_5731(w_eco5731, Tgate[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_5732(w_eco5732, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[1]);
	and _ECO_5733(w_eco5733, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[1]);
	and _ECO_5734(w_eco5734, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], prev_state[1]);
	and _ECO_5735(w_eco5735, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_5736(w_eco5736, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_5737(w_eco5737, Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5738(w_eco5738, prev_cnt[14], prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5739(w_eco5739, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5740(w_eco5740, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5741(w_eco5741, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5742(w_eco5742, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5743(w_eco5743, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5744(w_eco5744, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5745(w_eco5745, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_5746(w_eco5746, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_5747(w_eco5747, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5748(w_eco5748, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5749(w_eco5749, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], !ena);
	and _ECO_5750(w_eco5750, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], !ena);
	and _ECO_5751(w_eco5751, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], !ena);
	and _ECO_5752(w_eco5752, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], !ena);
	and _ECO_5753(w_eco5753, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], !ena);
	and _ECO_5754(w_eco5754, Tsync[4], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5755(w_eco5755, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5756(w_eco5756, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5757(w_eco5757, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5758(w_eco5758, !Tsync[4], Tgate[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5759(w_eco5759, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5760(w_eco5760, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5761(w_eco5761, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5762(w_eco5762, prev_cnt[1], prev_cnt[3], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5763(w_eco5763, prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5764(w_eco5764, prev_cnt[0], prev_cnt[3], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5765(w_eco5765, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5766(w_eco5766, Tgate[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_5767(w_eco5767, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5768(w_eco5768, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5769(w_eco5769, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5770(w_eco5770, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5771(w_eco5771, !Tsync[4], Tgate[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5772(w_eco5772, prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5773(w_eco5773, Tgdel[3], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5774(w_eco5774, prev_cnt[14], prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5775(w_eco5775, prev_cnt[1], prev_cnt[3], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5776(w_eco5776, prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5777(w_eco5777, prev_cnt[0], prev_cnt[3], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5778(w_eco5778, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5779(w_eco5779, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_5780(w_eco5780, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_5781(w_eco5781, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_5782(w_eco5782, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_5783(w_eco5783, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_5784(w_eco5784, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_5785(w_eco5785, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_5786(w_eco5786, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_5787(w_eco5787, !Tsync[3], !prev_cnt[14], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5788(w_eco5788, !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5789(w_eco5789, Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_5790(w_eco5790, prev_cnt[14], prev_cnt[2], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5791(w_eco5791, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5792(w_eco5792, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5793(w_eco5793, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5794(w_eco5794, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5795(w_eco5795, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5796(w_eco5796, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5797(w_eco5797, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[1]);
	and _ECO_5798(w_eco5798, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_state[1]);
	and _ECO_5799(w_eco5799, Tgdel[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5800(w_eco5800, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[1]);
	and _ECO_5801(w_eco5801, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[1]);
	and _ECO_5802(w_eco5802, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], prev_state[1]);
	and _ECO_5803(w_eco5803, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_5804(w_eco5804, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_5805(w_eco5805, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_5806(w_eco5806, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_5807(w_eco5807, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5808(w_eco5808, prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5809(w_eco5809, Tgdel[3], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5810(w_eco5810, prev_cnt[14], prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5811(w_eco5811, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5812(w_eco5812, Tgate[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5813(w_eco5813, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5814(w_eco5814, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5815(w_eco5815, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5816(w_eco5816, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5817(w_eco5817, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5818(w_eco5818, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5819(w_eco5819, !Tsync[4], Tgate[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_5820(w_eco5820, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_5821(w_eco5821, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_5822(w_eco5822, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5823(w_eco5823, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5824(w_eco5824, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], !ena);
	and _ECO_5825(w_eco5825, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], !ena);
	and _ECO_5826(w_eco5826, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], !ena);
	and _ECO_5827(w_eco5827, !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !ena);
	and _ECO_5828(w_eco5828, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], !ena);
	and _ECO_5829(w_eco5829, Tsync[4], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5830(w_eco5830, Tsync[4], !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5831(w_eco5831, Tsync[4], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5832(w_eco5832, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5833(w_eco5833, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5834(w_eco5834, !Tsync[4], Tgdel[3], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5835(w_eco5835, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5836(w_eco5836, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5837(w_eco5837, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5838(w_eco5838, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5839(w_eco5839, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5840(w_eco5840, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5841(w_eco5841, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5842(w_eco5842, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5843(w_eco5843, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5844(w_eco5844, Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_5845(w_eco5845, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5846(w_eco5846, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5847(w_eco5847, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5848(w_eco5848, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5849(w_eco5849, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5850(w_eco5850, !Tsync[4], Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_5851(w_eco5851, Tgdel[3], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5852(w_eco5852, prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5853(w_eco5853, Tgdel[3], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5854(w_eco5854, Tgdel[3], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5855(w_eco5855, !prev_cnt[14], prev_cnt[1], prev_cnt[3], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5856(w_eco5856, prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5857(w_eco5857, prev_cnt[0], prev_cnt[3], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5858(w_eco5858, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5859(w_eco5859, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5860(w_eco5860, Tgdel[3], prev_cnt[14], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_5861(w_eco5861, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_5862(w_eco5862, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_state[3], prev_state[0]);
	and _ECO_5863(w_eco5863, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_5864(w_eco5864, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_5865(w_eco5865, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_5866(w_eco5866, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_5867(w_eco5867, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_5868(w_eco5868, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_5869(w_eco5869, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_5870(w_eco5870, !Tsync[3], !prev_cnt[14], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5871(w_eco5871, prev_cnt[1], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5872(w_eco5872, !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5873(w_eco5873, Tgdel[3], prev_cnt[14], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_5874(w_eco5874, prev_cnt[14], prev_cnt[0], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5875(w_eco5875, Tgdel[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_5876(w_eco5876, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5877(w_eco5877, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5878(w_eco5878, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5879(w_eco5879, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5880(w_eco5880, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5881(w_eco5881, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5882(w_eco5882, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5883(w_eco5883, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[1]);
	and _ECO_5884(w_eco5884, Tgate[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_5885(w_eco5885, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[1]);
	and _ECO_5886(w_eco5886, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_state[1]);
	and _ECO_5887(w_eco5887, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[1]);
	and _ECO_5888(w_eco5888, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], prev_state[1]);
	and _ECO_5889(w_eco5889, !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_5890(w_eco5890, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_5891(w_eco5891, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_5892(w_eco5892, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_5893(w_eco5893, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5894(w_eco5894, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_5895(w_eco5895, Tgdel[3], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5896(w_eco5896, prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5897(w_eco5897, Tgdel[3], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5898(w_eco5898, Tgdel[3], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5899(w_eco5899, !prev_cnt[14], prev_cnt[1], prev_cnt[3], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5900(w_eco5900, prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5901(w_eco5901, prev_cnt[0], prev_cnt[3], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5902(w_eco5902, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5903(w_eco5903, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5904(w_eco5904, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5905(w_eco5905, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5906(w_eco5906, Tgdel[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_5907(w_eco5907, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5908(w_eco5908, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5909(w_eco5909, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5910(w_eco5910, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5911(w_eco5911, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5912(w_eco5912, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5913(w_eco5913, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5914(w_eco5914, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5915(w_eco5915, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5916(w_eco5916, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5917(w_eco5917, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5918(w_eco5918, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5919(w_eco5919, !Tsync[4], Tgdel[3], prev_cnt[14], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_5920(w_eco5920, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5921(w_eco5921, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5922(w_eco5922, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_5923(w_eco5923, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_5924(w_eco5924, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_5925(w_eco5925, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5926(w_eco5926, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], !ena);
	and _ECO_5927(w_eco5927, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], !ena);
	and _ECO_5928(w_eco5928, Tsync[4], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5929(w_eco5929, Tsync[4], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5930(w_eco5930, Tsync[4], !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5931(w_eco5931, Tsync[4], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5932(w_eco5932, Tsync[4], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5933(w_eco5933, !Tsync[4], Tgate[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_5934(w_eco5934, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5935(w_eco5935, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5936(w_eco5936, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5937(w_eco5937, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5938(w_eco5938, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5939(w_eco5939, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5940(w_eco5940, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_5941(w_eco5941, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5942(w_eco5942, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5943(w_eco5943, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5944(w_eco5944, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5945(w_eco5945, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5946(w_eco5946, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5947(w_eco5947, Tgate[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_5948(w_eco5948, Tgdel[3], prev_cnt[14], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_5949(w_eco5949, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5950(w_eco5950, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5951(w_eco5951, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5952(w_eco5952, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5953(w_eco5953, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_5954(w_eco5954, !Tsync[4], Tgate[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_5955(w_eco5955, Tgdel[3], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_5956(w_eco5956, prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5957(w_eco5957, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5958(w_eco5958, Tgdel[3], prev_cnt[14], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_5959(w_eco5959, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_5960(w_eco5960, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_5961(w_eco5961, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_state[3], prev_state[0]);
	and _ECO_5962(w_eco5962, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_5963(w_eco5963, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_5964(w_eco5964, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_5965(w_eco5965, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], !prev_state[4], !prev_state[2]);
	and _ECO_5966(w_eco5966, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_5967(w_eco5967, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_5968(w_eco5968, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_5969(w_eco5969, Tgdel[3], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_5970(w_eco5970, prev_cnt[2], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5971(w_eco5971, !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5972(w_eco5972, Tgdel[3], prev_cnt[14], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_5973(w_eco5973, !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5974(w_eco5974, Tgdel[3], prev_cnt[14], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_5975(w_eco5975, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5976(w_eco5976, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5977(w_eco5977, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5978(w_eco5978, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5979(w_eco5979, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_5980(w_eco5980, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_5981(w_eco5981, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5982(w_eco5982, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5983(w_eco5983, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_5984(w_eco5984, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5985(w_eco5985, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5986(w_eco5986, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_5987(w_eco5987, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_5988(w_eco5988, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_5989(w_eco5989, Tgate[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5990(w_eco5990, !prev_cnt[14], prev_cnt[1], prev_cnt[3], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5991(w_eco5991, !prev_cnt[14], prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5992(w_eco5992, prev_cnt[0], prev_cnt[3], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5993(w_eco5993, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_5994(w_eco5994, Tgdel[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_5995(w_eco5995, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[1]);
	and _ECO_5996(w_eco5996, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[1]);
	and _ECO_5997(w_eco5997, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], prev_state[1]);
	and _ECO_5998(w_eco5998, !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_state[1]);
	and _ECO_5999(w_eco5999, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_state[1]);
	and _ECO_6000(w_eco6000, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_6001(w_eco6001, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], !prev_state[3], prev_state[0]);
	and _ECO_6002(w_eco6002, !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_6003(w_eco6003, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_6004(w_eco6004, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_6005(w_eco6005, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6006(w_eco6006, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6007(w_eco6007, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6008(w_eco6008, Tgdel[3], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6009(w_eco6009, prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6010(w_eco6010, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_6011(w_eco6011, !Tgate[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_6012(w_eco6012, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6013(w_eco6013, Tgate[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_6014(w_eco6014, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6015(w_eco6015, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6016(w_eco6016, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6017(w_eco6017, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6018(w_eco6018, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6019(w_eco6019, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6020(w_eco6020, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6021(w_eco6021, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6022(w_eco6022, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6023(w_eco6023, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6024(w_eco6024, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6025(w_eco6025, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6026(w_eco6026, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6027(w_eco6027, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6028(w_eco6028, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6029(w_eco6029, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6030(w_eco6030, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6031(w_eco6031, !Tsync[4], Tgate[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_6032(w_eco6032, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6033(w_eco6033, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_6034(w_eco6034, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_6035(w_eco6035, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_6036(w_eco6036, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6037(w_eco6037, Tsync[4], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6038(w_eco6038, Tsync[4], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6039(w_eco6039, Tsync[4], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6040(w_eco6040, Tsync[4], !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6041(w_eco6041, Tsync[4], !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6042(w_eco6042, !Tsync[4], Tgdel[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_6043(w_eco6043, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6044(w_eco6044, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6045(w_eco6045, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6046(w_eco6046, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6047(w_eco6047, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6048(w_eco6048, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6049(w_eco6049, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6050(w_eco6050, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6051(w_eco6051, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6052(w_eco6052, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6053(w_eco6053, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6054(w_eco6054, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6055(w_eco6055, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6056(w_eco6056, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6057(w_eco6057, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6058(w_eco6058, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6059(w_eco6059, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6060(w_eco6060, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6061(w_eco6061, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6062(w_eco6062, Tgdel[3], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6063(w_eco6063, Tgdel[3], prev_cnt[14], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6064(w_eco6064, Tgdel[3], prev_cnt[14], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6065(w_eco6065, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6066(w_eco6066, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6067(w_eco6067, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6068(w_eco6068, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6069(w_eco6069, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6070(w_eco6070, !Tsync[4], Tgdel[3], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_6071(w_eco6071, !Tsync[4], Tgdel[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_6072(w_eco6072, Tgdel[3], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_6073(w_eco6073, Tgdel[3], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_6074(w_eco6074, !prev_cnt[14], prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6075(w_eco6075, !prev_cnt[14], prev_cnt[0], prev_cnt[3], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6076(w_eco6076, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6077(w_eco6077, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6078(w_eco6078, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6079(w_eco6079, Tgate[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6080(w_eco6080, !prev_cnt[14], prev_cnt[1], prev_cnt[3], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6081(w_eco6081, !prev_cnt[14], prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6082(w_eco6082, prev_cnt[0], prev_cnt[3], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6083(w_eco6083, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6084(w_eco6084, Tgdel[3], prev_cnt[1], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6085(w_eco6085, Tgdel[3], prev_cnt[14], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6086(w_eco6086, Tgdel[3], prev_cnt[14], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6087(w_eco6087, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_6088(w_eco6088, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_6089(w_eco6089, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_6090(w_eco6090, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_state[3], prev_state[0]);
	and _ECO_6091(w_eco6091, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_state[3], prev_state[0]);
	and _ECO_6092(w_eco6092, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_6093(w_eco6093, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_6094(w_eco6094, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_state[4], !prev_state[2]);
	and _ECO_6095(w_eco6095, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_6096(w_eco6096, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_6097(w_eco6097, Tgdel[3], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_6098(w_eco6098, prev_cnt[0], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6099(w_eco6099, Tgdel[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_6100(w_eco6100, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6101(w_eco6101, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6102(w_eco6102, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6103(w_eco6103, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6104(w_eco6104, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6105(w_eco6105, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6106(w_eco6106, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6107(w_eco6107, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6108(w_eco6108, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6109(w_eco6109, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6110(w_eco6110, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6111(w_eco6111, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6112(w_eco6112, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6113(w_eco6113, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6114(w_eco6114, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6115(w_eco6115, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6116(w_eco6116, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6117(w_eco6117, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6118(w_eco6118, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[1]);
	and _ECO_6119(w_eco6119, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], prev_state[1]);
	and _ECO_6120(w_eco6120, !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_6121(w_eco6121, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_6122(w_eco6122, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_state[3], prev_state[0]);
	and _ECO_6123(w_eco6123, !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_6124(w_eco6124, !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_6125(w_eco6125, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6126(w_eco6126, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6127(w_eco6127, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6128(w_eco6128, Tgdel[3], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6129(w_eco6129, Tgdel[3], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6130(w_eco6130, !prev_cnt[14], prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6131(w_eco6131, !prev_cnt[14], prev_cnt[0], prev_cnt[3], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6132(w_eco6132, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6133(w_eco6133, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6134(w_eco6134, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_6135(w_eco6135, !Tgate[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_6136(w_eco6136, Tgdel[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_6137(w_eco6137, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6138(w_eco6138, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6139(w_eco6139, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6140(w_eco6140, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6141(w_eco6141, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6142(w_eco6142, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6143(w_eco6143, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6144(w_eco6144, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6145(w_eco6145, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6146(w_eco6146, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6147(w_eco6147, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6148(w_eco6148, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6149(w_eco6149, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6150(w_eco6150, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6151(w_eco6151, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6152(w_eco6152, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6153(w_eco6153, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6154(w_eco6154, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6155(w_eco6155, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6156(w_eco6156, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6157(w_eco6157, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6158(w_eco6158, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6159(w_eco6159, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6160(w_eco6160, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6161(w_eco6161, !Tsync[4], Tgdel[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_6162(w_eco6162, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6163(w_eco6163, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_6164(w_eco6164, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_6165(w_eco6165, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_6166(w_eco6166, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_6167(w_eco6167, Tsync[4], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6168(w_eco6168, Tsync[4], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6169(w_eco6169, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6170(w_eco6170, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6171(w_eco6171, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6172(w_eco6172, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6173(w_eco6173, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6174(w_eco6174, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6175(w_eco6175, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6176(w_eco6176, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6177(w_eco6177, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6178(w_eco6178, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6179(w_eco6179, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6180(w_eco6180, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6181(w_eco6181, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6182(w_eco6182, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6183(w_eco6183, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6184(w_eco6184, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6185(w_eco6185, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6186(w_eco6186, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6187(w_eco6187, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6188(w_eco6188, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6189(w_eco6189, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6190(w_eco6190, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6191(w_eco6191, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6192(w_eco6192, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6193(w_eco6193, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6194(w_eco6194, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6195(w_eco6195, !prev_cnt[14], prev_cnt[0], prev_cnt[3], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6196(w_eco6196, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6197(w_eco6197, Tgdel[3], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6198(w_eco6198, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6199(w_eco6199, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_6200(w_eco6200, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6201(w_eco6201, !prev_cnt[14], prev_cnt[0], prev_cnt[3], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6202(w_eco6202, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6203(w_eco6203, Tgdel[3], prev_cnt[2], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6204(w_eco6204, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_6205(w_eco6205, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_6206(w_eco6206, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_6207(w_eco6207, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_6208(w_eco6208, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_6209(w_eco6209, !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], !prev_state[4], !prev_state[2]);
	and _ECO_6210(w_eco6210, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_state[4], !prev_state[2]);
	and _ECO_6211(w_eco6211, Tgdel[3], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_6212(w_eco6212, Tgdel[3], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_6213(w_eco6213, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6214(w_eco6214, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6215(w_eco6215, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6216(w_eco6216, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6217(w_eco6217, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6218(w_eco6218, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6219(w_eco6219, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6220(w_eco6220, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6221(w_eco6221, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6222(w_eco6222, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6223(w_eco6223, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6224(w_eco6224, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6225(w_eco6225, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6226(w_eco6226, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6227(w_eco6227, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6228(w_eco6228, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6229(w_eco6229, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6230(w_eco6230, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6231(w_eco6231, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6232(w_eco6232, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6233(w_eco6233, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6234(w_eco6234, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6235(w_eco6235, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6236(w_eco6236, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6237(w_eco6237, !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_6238(w_eco6238, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_6239(w_eco6239, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_6240(w_eco6240, !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], !prev_state[3], prev_state[0]);
	and _ECO_6241(w_eco6241, !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], !prev_state[3], prev_state[0]);
	and _ECO_6242(w_eco6242, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6243(w_eco6243, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6244(w_eco6244, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_6245(w_eco6245, !Tgate[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_6246(w_eco6246, !Tgate[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_6247(w_eco6247, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6248(w_eco6248, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6249(w_eco6249, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6250(w_eco6250, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6251(w_eco6251, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6252(w_eco6252, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6253(w_eco6253, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6254(w_eco6254, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6255(w_eco6255, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6256(w_eco6256, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6257(w_eco6257, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6258(w_eco6258, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6259(w_eco6259, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6260(w_eco6260, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6261(w_eco6261, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6262(w_eco6262, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6263(w_eco6263, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6264(w_eco6264, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6265(w_eco6265, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6266(w_eco6266, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6267(w_eco6267, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6268(w_eco6268, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6269(w_eco6269, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6270(w_eco6270, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6271(w_eco6271, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6272(w_eco6272, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6273(w_eco6273, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6274(w_eco6274, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6275(w_eco6275, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6276(w_eco6276, prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_6277(w_eco6277, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_6278(w_eco6278, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_6279(w_eco6279, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_6280(w_eco6280, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6281(w_eco6281, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6282(w_eco6282, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6283(w_eco6283, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6284(w_eco6284, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6285(w_eco6285, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6286(w_eco6286, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6287(w_eco6287, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6288(w_eco6288, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6289(w_eco6289, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6290(w_eco6290, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6291(w_eco6291, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6292(w_eco6292, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6293(w_eco6293, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6294(w_eco6294, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6295(w_eco6295, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6296(w_eco6296, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6297(w_eco6297, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6298(w_eco6298, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6299(w_eco6299, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6300(w_eco6300, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6301(w_eco6301, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6302(w_eco6302, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6303(w_eco6303, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6304(w_eco6304, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6305(w_eco6305, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6306(w_eco6306, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6307(w_eco6307, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6308(w_eco6308, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6309(w_eco6309, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6310(w_eco6310, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6311(w_eco6311, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6312(w_eco6312, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6313(w_eco6313, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_6314(w_eco6314, Tgdel[3], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6315(w_eco6315, Tgdel[3], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_6316(w_eco6316, !Tsync[4], Tgdel[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_6317(w_eco6317, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6318(w_eco6318, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_6319(w_eco6319, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_6320(w_eco6320, Tgdel[3], prev_cnt[3], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6321(w_eco6321, Tgdel[3], prev_cnt[0], !prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_6322(w_eco6322, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_6323(w_eco6323, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_6324(w_eco6324, !prev_cnt[14], prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_6325(w_eco6325, prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_6326(w_eco6326, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_6327(w_eco6327, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_6328(w_eco6328, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6329(w_eco6329, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6330(w_eco6330, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6331(w_eco6331, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6332(w_eco6332, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6333(w_eco6333, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6334(w_eco6334, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6335(w_eco6335, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6336(w_eco6336, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6337(w_eco6337, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6338(w_eco6338, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6339(w_eco6339, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6340(w_eco6340, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6341(w_eco6341, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6342(w_eco6342, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6343(w_eco6343, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6344(w_eco6344, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6345(w_eco6345, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6346(w_eco6346, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6347(w_eco6347, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6348(w_eco6348, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6349(w_eco6349, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6350(w_eco6350, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6351(w_eco6351, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6352(w_eco6352, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6353(w_eco6353, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6354(w_eco6354, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6355(w_eco6355, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6356(w_eco6356, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6357(w_eco6357, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6358(w_eco6358, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6359(w_eco6359, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6360(w_eco6360, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6361(w_eco6361, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6362(w_eco6362, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6363(w_eco6363, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6364(w_eco6364, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6365(w_eco6365, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6366(w_eco6366, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6367(w_eco6367, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6368(w_eco6368, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6369(w_eco6369, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_6370(w_eco6370, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6371(w_eco6371, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6372(w_eco6372, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6373(w_eco6373, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6374(w_eco6374, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6375(w_eco6375, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6376(w_eco6376, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6377(w_eco6377, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6378(w_eco6378, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6379(w_eco6379, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6380(w_eco6380, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6381(w_eco6381, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6382(w_eco6382, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6383(w_eco6383, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6384(w_eco6384, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6385(w_eco6385, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6386(w_eco6386, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6387(w_eco6387, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6388(w_eco6388, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6389(w_eco6389, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6390(w_eco6390, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6391(w_eco6391, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6392(w_eco6392, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6393(w_eco6393, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6394(w_eco6394, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6395(w_eco6395, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6396(w_eco6396, !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_6397(w_eco6397, !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_6398(w_eco6398, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6399(w_eco6399, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6400(w_eco6400, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6401(w_eco6401, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6402(w_eco6402, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_6403(w_eco6403, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6404(w_eco6404, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6405(w_eco6405, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6406(w_eco6406, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6407(w_eco6407, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6408(w_eco6408, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6409(w_eco6409, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6410(w_eco6410, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6411(w_eco6411, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6412(w_eco6412, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6413(w_eco6413, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6414(w_eco6414, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6415(w_eco6415, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6416(w_eco6416, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6417(w_eco6417, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6418(w_eco6418, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6419(w_eco6419, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6420(w_eco6420, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6421(w_eco6421, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6422(w_eco6422, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6423(w_eco6423, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6424(w_eco6424, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6425(w_eco6425, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6426(w_eco6426, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6427(w_eco6427, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6428(w_eco6428, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6429(w_eco6429, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6430(w_eco6430, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6431(w_eco6431, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6432(w_eco6432, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6433(w_eco6433, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6434(w_eco6434, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6435(w_eco6435, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6436(w_eco6436, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6437(w_eco6437, !prev_cnt[14], prev_cnt[1], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_6438(w_eco6438, !prev_cnt[14], prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_6439(w_eco6439, prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_6440(w_eco6440, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_6441(w_eco6441, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6442(w_eco6442, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6443(w_eco6443, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6444(w_eco6444, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6445(w_eco6445, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6446(w_eco6446, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6447(w_eco6447, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6448(w_eco6448, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6449(w_eco6449, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6450(w_eco6450, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6451(w_eco6451, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6452(w_eco6452, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6453(w_eco6453, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6454(w_eco6454, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6455(w_eco6455, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6456(w_eco6456, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6457(w_eco6457, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6458(w_eco6458, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6459(w_eco6459, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6460(w_eco6460, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6461(w_eco6461, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6462(w_eco6462, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6463(w_eco6463, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6464(w_eco6464, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6465(w_eco6465, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6466(w_eco6466, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6467(w_eco6467, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6468(w_eco6468, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6469(w_eco6469, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6470(w_eco6470, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6471(w_eco6471, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6472(w_eco6472, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6473(w_eco6473, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6474(w_eco6474, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6475(w_eco6475, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6476(w_eco6476, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6477(w_eco6477, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6478(w_eco6478, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6479(w_eco6479, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6480(w_eco6480, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6481(w_eco6481, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6482(w_eco6482, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6483(w_eco6483, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6484(w_eco6484, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6485(w_eco6485, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6486(w_eco6486, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6487(w_eco6487, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6488(w_eco6488, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6489(w_eco6489, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6490(w_eco6490, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6491(w_eco6491, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6492(w_eco6492, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6493(w_eco6493, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6494(w_eco6494, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6495(w_eco6495, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6496(w_eco6496, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6497(w_eco6497, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6498(w_eco6498, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6499(w_eco6499, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6500(w_eco6500, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6501(w_eco6501, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6502(w_eco6502, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6503(w_eco6503, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6504(w_eco6504, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6505(w_eco6505, !Tsync[4], Tsync[3], !prev_cnt[4], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6506(w_eco6506, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6507(w_eco6507, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6508(w_eco6508, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6509(w_eco6509, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6510(w_eco6510, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6511(w_eco6511, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6512(w_eco6512, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6513(w_eco6513, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6514(w_eco6514, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6515(w_eco6515, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6516(w_eco6516, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6517(w_eco6517, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6518(w_eco6518, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6519(w_eco6519, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6520(w_eco6520, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6521(w_eco6521, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6522(w_eco6522, Tsync[4], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6523(w_eco6523, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6524(w_eco6524, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6525(w_eco6525, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6526(w_eco6526, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6527(w_eco6527, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6528(w_eco6528, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6529(w_eco6529, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6530(w_eco6530, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6531(w_eco6531, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6532(w_eco6532, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6533(w_eco6533, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6534(w_eco6534, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6535(w_eco6535, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6536(w_eco6536, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6537(w_eco6537, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6538(w_eco6538, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6539(w_eco6539, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6540(w_eco6540, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6541(w_eco6541, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6542(w_eco6542, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6543(w_eco6543, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6544(w_eco6544, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6545(w_eco6545, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6546(w_eco6546, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6547(w_eco6547, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6548(w_eco6548, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6549(w_eco6549, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6550(w_eco6550, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6551(w_eco6551, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6552(w_eco6552, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6553(w_eco6553, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6554(w_eco6554, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6555(w_eco6555, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6556(w_eco6556, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6557(w_eco6557, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6558(w_eco6558, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6559(w_eco6559, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6560(w_eco6560, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6561(w_eco6561, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6562(w_eco6562, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6563(w_eco6563, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6564(w_eco6564, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6565(w_eco6565, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6566(w_eco6566, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6567(w_eco6567, !prev_cnt[14], prev_cnt[2], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_6568(w_eco6568, !prev_cnt[14], prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_6569(w_eco6569, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_6570(w_eco6570, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6571(w_eco6571, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6572(w_eco6572, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6573(w_eco6573, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6574(w_eco6574, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6575(w_eco6575, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6576(w_eco6576, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6577(w_eco6577, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6578(w_eco6578, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6579(w_eco6579, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6580(w_eco6580, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6581(w_eco6581, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6582(w_eco6582, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6583(w_eco6583, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6584(w_eco6584, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6585(w_eco6585, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6586(w_eco6586, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6587(w_eco6587, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6588(w_eco6588, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6589(w_eco6589, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6590(w_eco6590, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6591(w_eco6591, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6592(w_eco6592, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6593(w_eco6593, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6594(w_eco6594, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6595(w_eco6595, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6596(w_eco6596, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6597(w_eco6597, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6598(w_eco6598, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6599(w_eco6599, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6600(w_eco6600, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6601(w_eco6601, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6602(w_eco6602, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6603(w_eco6603, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6604(w_eco6604, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6605(w_eco6605, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6606(w_eco6606, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6607(w_eco6607, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6608(w_eco6608, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6609(w_eco6609, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6610(w_eco6610, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6611(w_eco6611, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6612(w_eco6612, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6613(w_eco6613, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6614(w_eco6614, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6615(w_eco6615, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6616(w_eco6616, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6617(w_eco6617, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6618(w_eco6618, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6619(w_eco6619, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6620(w_eco6620, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6621(w_eco6621, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6622(w_eco6622, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6623(w_eco6623, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6624(w_eco6624, !Tsync[4], Tsync[3], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6625(w_eco6625, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6626(w_eco6626, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6627(w_eco6627, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6628(w_eco6628, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6629(w_eco6629, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6630(w_eco6630, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6631(w_eco6631, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6632(w_eco6632, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6633(w_eco6633, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6634(w_eco6634, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6635(w_eco6635, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6636(w_eco6636, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6637(w_eco6637, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6638(w_eco6638, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6639(w_eco6639, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6640(w_eco6640, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6641(w_eco6641, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6642(w_eco6642, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6643(w_eco6643, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6644(w_eco6644, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6645(w_eco6645, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6646(w_eco6646, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6647(w_eco6647, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6648(w_eco6648, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6649(w_eco6649, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6650(w_eco6650, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6651(w_eco6651, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6652(w_eco6652, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6653(w_eco6653, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6654(w_eco6654, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6655(w_eco6655, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6656(w_eco6656, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6657(w_eco6657, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6658(w_eco6658, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6659(w_eco6659, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6660(w_eco6660, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6661(w_eco6661, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6662(w_eco6662, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6663(w_eco6663, !Tsync[4], Tsync[3], !prev_cnt[4], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6664(w_eco6664, !Tsync[4], Tsync[3], !prev_cnt[4], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6665(w_eco6665, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6666(w_eco6666, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[1], !prev_cnt[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6667(w_eco6667, Tsync[4], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6668(w_eco6668, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6669(w_eco6669, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6670(w_eco6670, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6671(w_eco6671, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6672(w_eco6672, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6673(w_eco6673, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6674(w_eco6674, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6675(w_eco6675, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6676(w_eco6676, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6677(w_eco6677, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6678(w_eco6678, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6679(w_eco6679, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6680(w_eco6680, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6681(w_eco6681, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6682(w_eco6682, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6683(w_eco6683, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6684(w_eco6684, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6685(w_eco6685, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6686(w_eco6686, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6687(w_eco6687, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6688(w_eco6688, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6689(w_eco6689, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6690(w_eco6690, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6691(w_eco6691, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6692(w_eco6692, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6693(w_eco6693, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6694(w_eco6694, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6695(w_eco6695, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6696(w_eco6696, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6697(w_eco6697, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6698(w_eco6698, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6699(w_eco6699, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6700(w_eco6700, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6701(w_eco6701, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6702(w_eco6702, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6703(w_eco6703, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6704(w_eco6704, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6705(w_eco6705, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6706(w_eco6706, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6707(w_eco6707, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6708(w_eco6708, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6709(w_eco6709, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6710(w_eco6710, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6711(w_eco6711, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6712(w_eco6712, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6713(w_eco6713, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6714(w_eco6714, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6715(w_eco6715, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6716(w_eco6716, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6717(w_eco6717, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6718(w_eco6718, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6719(w_eco6719, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6720(w_eco6720, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6721(w_eco6721, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6722(w_eco6722, !prev_cnt[14], prev_cnt[0], prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_6723(w_eco6723, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_6724(w_eco6724, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6725(w_eco6725, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6726(w_eco6726, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6727(w_eco6727, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6728(w_eco6728, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6729(w_eco6729, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6730(w_eco6730, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6731(w_eco6731, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6732(w_eco6732, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6733(w_eco6733, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6734(w_eco6734, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6735(w_eco6735, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6736(w_eco6736, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6737(w_eco6737, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6738(w_eco6738, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6739(w_eco6739, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6740(w_eco6740, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6741(w_eco6741, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6742(w_eco6742, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6743(w_eco6743, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6744(w_eco6744, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6745(w_eco6745, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6746(w_eco6746, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6747(w_eco6747, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6748(w_eco6748, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6749(w_eco6749, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6750(w_eco6750, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6751(w_eco6751, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6752(w_eco6752, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6753(w_eco6753, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6754(w_eco6754, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6755(w_eco6755, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6756(w_eco6756, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6757(w_eco6757, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6758(w_eco6758, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6759(w_eco6759, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6760(w_eco6760, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6761(w_eco6761, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6762(w_eco6762, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6763(w_eco6763, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6764(w_eco6764, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6765(w_eco6765, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6766(w_eco6766, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6767(w_eco6767, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6768(w_eco6768, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6769(w_eco6769, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6770(w_eco6770, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6771(w_eco6771, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6772(w_eco6772, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6773(w_eco6773, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6774(w_eco6774, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6775(w_eco6775, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6776(w_eco6776, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6777(w_eco6777, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6778(w_eco6778, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6779(w_eco6779, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6780(w_eco6780, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6781(w_eco6781, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6782(w_eco6782, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6783(w_eco6783, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6784(w_eco6784, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6785(w_eco6785, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6786(w_eco6786, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6787(w_eco6787, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6788(w_eco6788, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6789(w_eco6789, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6790(w_eco6790, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6791(w_eco6791, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6792(w_eco6792, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6793(w_eco6793, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6794(w_eco6794, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6795(w_eco6795, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6796(w_eco6796, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6797(w_eco6797, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6798(w_eco6798, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6799(w_eco6799, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6800(w_eco6800, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6801(w_eco6801, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6802(w_eco6802, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6803(w_eco6803, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6804(w_eco6804, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6805(w_eco6805, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6806(w_eco6806, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6807(w_eco6807, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6808(w_eco6808, !Tsync[4], Tsync[3], !prev_cnt[4], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6809(w_eco6809, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6810(w_eco6810, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6811(w_eco6811, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6812(w_eco6812, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6813(w_eco6813, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6814(w_eco6814, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6815(w_eco6815, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6816(w_eco6816, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6817(w_eco6817, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6818(w_eco6818, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6819(w_eco6819, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6820(w_eco6820, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6821(w_eco6821, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6822(w_eco6822, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6823(w_eco6823, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6824(w_eco6824, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6825(w_eco6825, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6826(w_eco6826, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6827(w_eco6827, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6828(w_eco6828, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6829(w_eco6829, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6830(w_eco6830, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6831(w_eco6831, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[2], !prev_cnt[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6832(w_eco6832, Tsync[4], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6833(w_eco6833, Tsync[4], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_6834(w_eco6834, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6835(w_eco6835, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6836(w_eco6836, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6837(w_eco6837, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6838(w_eco6838, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6839(w_eco6839, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6840(w_eco6840, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6841(w_eco6841, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6842(w_eco6842, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6843(w_eco6843, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6844(w_eco6844, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6845(w_eco6845, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6846(w_eco6846, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6847(w_eco6847, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6848(w_eco6848, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6849(w_eco6849, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6850(w_eco6850, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6851(w_eco6851, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6852(w_eco6852, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6853(w_eco6853, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6854(w_eco6854, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6855(w_eco6855, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6856(w_eco6856, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6857(w_eco6857, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6858(w_eco6858, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6859(w_eco6859, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6860(w_eco6860, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6861(w_eco6861, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6862(w_eco6862, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6863(w_eco6863, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6864(w_eco6864, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6865(w_eco6865, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6866(w_eco6866, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6867(w_eco6867, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6868(w_eco6868, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6869(w_eco6869, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6870(w_eco6870, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6871(w_eco6871, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6872(w_eco6872, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6873(w_eco6873, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6874(w_eco6874, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6875(w_eco6875, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6876(w_eco6876, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6877(w_eco6877, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6878(w_eco6878, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6879(w_eco6879, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6880(w_eco6880, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6881(w_eco6881, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6882(w_eco6882, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6883(w_eco6883, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6884(w_eco6884, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6885(w_eco6885, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6886(w_eco6886, Tsync[3], !prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6887(w_eco6887, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6888(w_eco6888, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6889(w_eco6889, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6890(w_eco6890, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6891(w_eco6891, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_6892(w_eco6892, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6893(w_eco6893, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6894(w_eco6894, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_6895(w_eco6895, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6896(w_eco6896, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6897(w_eco6897, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_6898(w_eco6898, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6899(w_eco6899, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6900(w_eco6900, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6901(w_eco6901, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6902(w_eco6902, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6903(w_eco6903, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6904(w_eco6904, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6905(w_eco6905, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6906(w_eco6906, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6907(w_eco6907, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6908(w_eco6908, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6909(w_eco6909, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6910(w_eco6910, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6911(w_eco6911, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6912(w_eco6912, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6913(w_eco6913, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6914(w_eco6914, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6915(w_eco6915, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6916(w_eco6916, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6917(w_eco6917, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6918(w_eco6918, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6919(w_eco6919, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6920(w_eco6920, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6921(w_eco6921, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6922(w_eco6922, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6923(w_eco6923, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6924(w_eco6924, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6925(w_eco6925, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6926(w_eco6926, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6927(w_eco6927, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6928(w_eco6928, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6929(w_eco6929, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6930(w_eco6930, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6931(w_eco6931, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6932(w_eco6932, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6933(w_eco6933, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6934(w_eco6934, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6935(w_eco6935, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6936(w_eco6936, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6937(w_eco6937, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6938(w_eco6938, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6939(w_eco6939, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6940(w_eco6940, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6941(w_eco6941, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6942(w_eco6942, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6943(w_eco6943, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6944(w_eco6944, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6945(w_eco6945, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6946(w_eco6946, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6947(w_eco6947, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6948(w_eco6948, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6949(w_eco6949, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6950(w_eco6950, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6951(w_eco6951, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6952(w_eco6952, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6953(w_eco6953, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6954(w_eco6954, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6955(w_eco6955, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6956(w_eco6956, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6957(w_eco6957, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6958(w_eco6958, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6959(w_eco6959, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6960(w_eco6960, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6961(w_eco6961, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6962(w_eco6962, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6963(w_eco6963, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6964(w_eco6964, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6965(w_eco6965, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6966(w_eco6966, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6967(w_eco6967, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6968(w_eco6968, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_6969(w_eco6969, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6970(w_eco6970, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6971(w_eco6971, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6972(w_eco6972, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6973(w_eco6973, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6974(w_eco6974, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6975(w_eco6975, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6976(w_eco6976, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6977(w_eco6977, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6978(w_eco6978, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6979(w_eco6979, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6980(w_eco6980, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6981(w_eco6981, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6982(w_eco6982, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6983(w_eco6983, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6984(w_eco6984, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6985(w_eco6985, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6986(w_eco6986, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6987(w_eco6987, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6988(w_eco6988, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6989(w_eco6989, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6990(w_eco6990, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6991(w_eco6991, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6992(w_eco6992, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_6993(w_eco6993, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6994(w_eco6994, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6995(w_eco6995, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6996(w_eco6996, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6997(w_eco6997, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_6998(w_eco6998, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_6999(w_eco6999, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7000(w_eco7000, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7001(w_eco7001, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7002(w_eco7002, !Tsync[4], Tsync[3], !prev_cnt[4], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7003(w_eco7003, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7004(w_eco7004, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7005(w_eco7005, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7006(w_eco7006, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7007(w_eco7007, Tsync[4], !Tgate[3], !Tgdel[3], !Tsync[3], prev_cnt[0], !prev_cnt[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7008(w_eco7008, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7009(w_eco7009, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7010(w_eco7010, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7011(w_eco7011, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7012(w_eco7012, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7013(w_eco7013, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7014(w_eco7014, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7015(w_eco7015, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7016(w_eco7016, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7017(w_eco7017, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7018(w_eco7018, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7019(w_eco7019, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7020(w_eco7020, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7021(w_eco7021, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7022(w_eco7022, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7023(w_eco7023, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7024(w_eco7024, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7025(w_eco7025, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7026(w_eco7026, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7027(w_eco7027, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7028(w_eco7028, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7029(w_eco7029, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7030(w_eco7030, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7031(w_eco7031, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7032(w_eco7032, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7033(w_eco7033, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7034(w_eco7034, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7035(w_eco7035, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7036(w_eco7036, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7037(w_eco7037, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7038(w_eco7038, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7039(w_eco7039, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7040(w_eco7040, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7041(w_eco7041, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7042(w_eco7042, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7043(w_eco7043, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7044(w_eco7044, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7045(w_eco7045, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7046(w_eco7046, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7047(w_eco7047, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7048(w_eco7048, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7049(w_eco7049, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7050(w_eco7050, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7051(w_eco7051, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7052(w_eco7052, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7053(w_eco7053, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7054(w_eco7054, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7055(w_eco7055, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7056(w_eco7056, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7057(w_eco7057, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7058(w_eco7058, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7059(w_eco7059, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7060(w_eco7060, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7061(w_eco7061, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7062(w_eco7062, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7063(w_eco7063, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7064(w_eco7064, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7065(w_eco7065, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7066(w_eco7066, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7067(w_eco7067, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7068(w_eco7068, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7069(w_eco7069, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7070(w_eco7070, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7071(w_eco7071, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7072(w_eco7072, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7073(w_eco7073, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7074(w_eco7074, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7075(w_eco7075, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7076(w_eco7076, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7077(w_eco7077, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7078(w_eco7078, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7079(w_eco7079, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7080(w_eco7080, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7081(w_eco7081, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7082(w_eco7082, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7083(w_eco7083, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7084(w_eco7084, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7085(w_eco7085, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7086(w_eco7086, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7087(w_eco7087, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7088(w_eco7088, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7089(w_eco7089, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7090(w_eco7090, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7091(w_eco7091, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7092(w_eco7092, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7093(w_eco7093, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7094(w_eco7094, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7095(w_eco7095, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7096(w_eco7096, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7097(w_eco7097, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7098(w_eco7098, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7099(w_eco7099, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7100(w_eco7100, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7101(w_eco7101, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7102(w_eco7102, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7103(w_eco7103, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7104(w_eco7104, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7105(w_eco7105, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7106(w_eco7106, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7107(w_eco7107, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7108(w_eco7108, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7109(w_eco7109, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7110(w_eco7110, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7111(w_eco7111, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7112(w_eco7112, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7113(w_eco7113, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7114(w_eco7114, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7115(w_eco7115, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7116(w_eco7116, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7117(w_eco7117, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7118(w_eco7118, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7119(w_eco7119, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7120(w_eco7120, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7121(w_eco7121, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7122(w_eco7122, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7123(w_eco7123, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7124(w_eco7124, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7125(w_eco7125, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7126(w_eco7126, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7127(w_eco7127, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7128(w_eco7128, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7129(w_eco7129, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7130(w_eco7130, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7131(w_eco7131, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7132(w_eco7132, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7133(w_eco7133, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7134(w_eco7134, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7135(w_eco7135, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7136(w_eco7136, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7137(w_eco7137, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7138(w_eco7138, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7139(w_eco7139, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7140(w_eco7140, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7141(w_eco7141, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7142(w_eco7142, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7143(w_eco7143, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7144(w_eco7144, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7145(w_eco7145, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7146(w_eco7146, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7147(w_eco7147, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7148(w_eco7148, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7149(w_eco7149, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7150(w_eco7150, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7151(w_eco7151, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7152(w_eco7152, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7153(w_eco7153, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7154(w_eco7154, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7155(w_eco7155, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7156(w_eco7156, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7157(w_eco7157, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7158(w_eco7158, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7159(w_eco7159, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7160(w_eco7160, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7161(w_eco7161, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7162(w_eco7162, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7163(w_eco7163, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7164(w_eco7164, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7165(w_eco7165, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7166(w_eco7166, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7167(w_eco7167, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7168(w_eco7168, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7169(w_eco7169, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7170(w_eco7170, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7171(w_eco7171, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7172(w_eco7172, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7173(w_eco7173, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7174(w_eco7174, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7175(w_eco7175, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7176(w_eco7176, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7177(w_eco7177, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7178(w_eco7178, Tsync[4], !Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7179(w_eco7179, Tsync[4], !Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7180(w_eco7180, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7181(w_eco7181, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7182(w_eco7182, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7183(w_eco7183, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7184(w_eco7184, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7185(w_eco7185, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7186(w_eco7186, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7187(w_eco7187, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7188(w_eco7188, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7189(w_eco7189, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7190(w_eco7190, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7191(w_eco7191, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7192(w_eco7192, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7193(w_eco7193, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7194(w_eco7194, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7195(w_eco7195, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7196(w_eco7196, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7197(w_eco7197, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7198(w_eco7198, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7199(w_eco7199, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7200(w_eco7200, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7201(w_eco7201, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7202(w_eco7202, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7203(w_eco7203, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7204(w_eco7204, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7205(w_eco7205, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7206(w_eco7206, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7207(w_eco7207, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7208(w_eco7208, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7209(w_eco7209, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7210(w_eco7210, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7211(w_eco7211, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7212(w_eco7212, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7213(w_eco7213, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7214(w_eco7214, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7215(w_eco7215, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7216(w_eco7216, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7217(w_eco7217, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7218(w_eco7218, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7219(w_eco7219, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7220(w_eco7220, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7221(w_eco7221, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7222(w_eco7222, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7223(w_eco7223, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7224(w_eco7224, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7225(w_eco7225, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7226(w_eco7226, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7227(w_eco7227, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7228(w_eco7228, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7229(w_eco7229, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7230(w_eco7230, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7231(w_eco7231, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7232(w_eco7232, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7233(w_eco7233, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7234(w_eco7234, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7235(w_eco7235, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7236(w_eco7236, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7237(w_eco7237, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7238(w_eco7238, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7239(w_eco7239, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7240(w_eco7240, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7241(w_eco7241, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7242(w_eco7242, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7243(w_eco7243, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7244(w_eco7244, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7245(w_eco7245, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7246(w_eco7246, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7247(w_eco7247, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7248(w_eco7248, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7249(w_eco7249, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7250(w_eco7250, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7251(w_eco7251, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7252(w_eco7252, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7253(w_eco7253, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7254(w_eco7254, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7255(w_eco7255, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7256(w_eco7256, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7257(w_eco7257, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7258(w_eco7258, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7259(w_eco7259, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7260(w_eco7260, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7261(w_eco7261, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7262(w_eco7262, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7263(w_eco7263, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7264(w_eco7264, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7265(w_eco7265, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7266(w_eco7266, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7267(w_eco7267, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7268(w_eco7268, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7269(w_eco7269, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7270(w_eco7270, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7271(w_eco7271, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7272(w_eco7272, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7273(w_eco7273, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7274(w_eco7274, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7275(w_eco7275, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7276(w_eco7276, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7277(w_eco7277, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7278(w_eco7278, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7279(w_eco7279, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7280(w_eco7280, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7281(w_eco7281, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7282(w_eco7282, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7283(w_eco7283, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7284(w_eco7284, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7285(w_eco7285, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7286(w_eco7286, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7287(w_eco7287, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7288(w_eco7288, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7289(w_eco7289, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7290(w_eco7290, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7291(w_eco7291, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7292(w_eco7292, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7293(w_eco7293, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7294(w_eco7294, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7295(w_eco7295, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7296(w_eco7296, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7297(w_eco7297, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7298(w_eco7298, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7299(w_eco7299, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7300(w_eco7300, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7301(w_eco7301, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7302(w_eco7302, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7303(w_eco7303, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7304(w_eco7304, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7305(w_eco7305, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7306(w_eco7306, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7307(w_eco7307, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7308(w_eco7308, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7309(w_eco7309, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7310(w_eco7310, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7311(w_eco7311, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7312(w_eco7312, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7313(w_eco7313, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7314(w_eco7314, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7315(w_eco7315, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7316(w_eco7316, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7317(w_eco7317, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7318(w_eco7318, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7319(w_eco7319, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7320(w_eco7320, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7321(w_eco7321, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7322(w_eco7322, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7323(w_eco7323, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7324(w_eco7324, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7325(w_eco7325, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7326(w_eco7326, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7327(w_eco7327, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7328(w_eco7328, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7329(w_eco7329, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7330(w_eco7330, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7331(w_eco7331, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7332(w_eco7332, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7333(w_eco7333, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7334(w_eco7334, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7335(w_eco7335, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7336(w_eco7336, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7337(w_eco7337, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7338(w_eco7338, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7339(w_eco7339, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7340(w_eco7340, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7341(w_eco7341, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7342(w_eco7342, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7343(w_eco7343, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7344(w_eco7344, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7345(w_eco7345, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7346(w_eco7346, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7347(w_eco7347, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7348(w_eco7348, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7349(w_eco7349, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7350(w_eco7350, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7351(w_eco7351, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7352(w_eco7352, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7353(w_eco7353, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7354(w_eco7354, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7355(w_eco7355, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7356(w_eco7356, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7357(w_eco7357, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7358(w_eco7358, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7359(w_eco7359, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7360(w_eco7360, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7361(w_eco7361, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7362(w_eco7362, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7363(w_eco7363, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7364(w_eco7364, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7365(w_eco7365, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7366(w_eco7366, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7367(w_eco7367, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7368(w_eco7368, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7369(w_eco7369, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7370(w_eco7370, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7371(w_eco7371, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7372(w_eco7372, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7373(w_eco7373, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7374(w_eco7374, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7375(w_eco7375, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7376(w_eco7376, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7377(w_eco7377, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7378(w_eco7378, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7379(w_eco7379, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7380(w_eco7380, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7381(w_eco7381, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7382(w_eco7382, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7383(w_eco7383, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7384(w_eco7384, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7385(w_eco7385, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7386(w_eco7386, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7387(w_eco7387, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7388(w_eco7388, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7389(w_eco7389, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7390(w_eco7390, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7391(w_eco7391, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7392(w_eco7392, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7393(w_eco7393, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7394(w_eco7394, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7395(w_eco7395, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7396(w_eco7396, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7397(w_eco7397, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7398(w_eco7398, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7399(w_eco7399, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7400(w_eco7400, prev_cnt[1], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7401(w_eco7401, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7402(w_eco7402, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7403(w_eco7403, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7404(w_eco7404, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7405(w_eco7405, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7406(w_eco7406, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7407(w_eco7407, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7408(w_eco7408, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7409(w_eco7409, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7410(w_eco7410, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7411(w_eco7411, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7412(w_eco7412, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7413(w_eco7413, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7414(w_eco7414, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7415(w_eco7415, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7416(w_eco7416, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7417(w_eco7417, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7418(w_eco7418, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7419(w_eco7419, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7420(w_eco7420, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7421(w_eco7421, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7422(w_eco7422, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7423(w_eco7423, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7424(w_eco7424, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7425(w_eco7425, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7426(w_eco7426, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7427(w_eco7427, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7428(w_eco7428, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7429(w_eco7429, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7430(w_eco7430, Tsync[4], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7431(w_eco7431, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7432(w_eco7432, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7433(w_eco7433, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7434(w_eco7434, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7435(w_eco7435, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7436(w_eco7436, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7437(w_eco7437, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7438(w_eco7438, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7439(w_eco7439, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7440(w_eco7440, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7441(w_eco7441, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7442(w_eco7442, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7443(w_eco7443, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7444(w_eco7444, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7445(w_eco7445, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7446(w_eco7446, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7447(w_eco7447, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7448(w_eco7448, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7449(w_eco7449, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7450(w_eco7450, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7451(w_eco7451, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7452(w_eco7452, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7453(w_eco7453, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7454(w_eco7454, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7455(w_eco7455, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7456(w_eco7456, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_7457(w_eco7457, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7458(w_eco7458, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7459(w_eco7459, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7460(w_eco7460, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7461(w_eco7461, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7462(w_eco7462, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7463(w_eco7463, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7464(w_eco7464, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7465(w_eco7465, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7466(w_eco7466, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7467(w_eco7467, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7468(w_eco7468, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7469(w_eco7469, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7470(w_eco7470, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7471(w_eco7471, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7472(w_eco7472, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7473(w_eco7473, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7474(w_eco7474, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7475(w_eco7475, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7476(w_eco7476, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7477(w_eco7477, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7478(w_eco7478, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7479(w_eco7479, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7480(w_eco7480, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7481(w_eco7481, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7482(w_eco7482, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7483(w_eco7483, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7484(w_eco7484, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7485(w_eco7485, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7486(w_eco7486, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7487(w_eco7487, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7488(w_eco7488, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7489(w_eco7489, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7490(w_eco7490, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7491(w_eco7491, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7492(w_eco7492, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7493(w_eco7493, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7494(w_eco7494, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7495(w_eco7495, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7496(w_eco7496, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7497(w_eco7497, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7498(w_eco7498, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7499(w_eco7499, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7500(w_eco7500, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7501(w_eco7501, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7502(w_eco7502, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7503(w_eco7503, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7504(w_eco7504, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7505(w_eco7505, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7506(w_eco7506, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7507(w_eco7507, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7508(w_eco7508, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7509(w_eco7509, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7510(w_eco7510, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7511(w_eco7511, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7512(w_eco7512, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7513(w_eco7513, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7514(w_eco7514, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7515(w_eco7515, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7516(w_eco7516, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7517(w_eco7517, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7518(w_eco7518, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7519(w_eco7519, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7520(w_eco7520, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7521(w_eco7521, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7522(w_eco7522, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7523(w_eco7523, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7524(w_eco7524, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7525(w_eco7525, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7526(w_eco7526, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7527(w_eco7527, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7528(w_eco7528, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7529(w_eco7529, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7530(w_eco7530, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7531(w_eco7531, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7532(w_eco7532, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7533(w_eco7533, prev_cnt[2], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7534(w_eco7534, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7535(w_eco7535, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7536(w_eco7536, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7537(w_eco7537, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7538(w_eco7538, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7539(w_eco7539, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7540(w_eco7540, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7541(w_eco7541, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7542(w_eco7542, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7543(w_eco7543, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7544(w_eco7544, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7545(w_eco7545, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7546(w_eco7546, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7547(w_eco7547, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7548(w_eco7548, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7549(w_eco7549, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7550(w_eco7550, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7551(w_eco7551, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7552(w_eco7552, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7553(w_eco7553, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7554(w_eco7554, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7555(w_eco7555, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7556(w_eco7556, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7557(w_eco7557, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7558(w_eco7558, Tsync[4], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7559(w_eco7559, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7560(w_eco7560, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7561(w_eco7561, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7562(w_eco7562, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7563(w_eco7563, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7564(w_eco7564, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7565(w_eco7565, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7566(w_eco7566, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7567(w_eco7567, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7568(w_eco7568, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7569(w_eco7569, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7570(w_eco7570, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7571(w_eco7571, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7572(w_eco7572, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7573(w_eco7573, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7574(w_eco7574, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7575(w_eco7575, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7576(w_eco7576, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7577(w_eco7577, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7578(w_eco7578, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7579(w_eco7579, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7580(w_eco7580, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7581(w_eco7581, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7582(w_eco7582, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7583(w_eco7583, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7584(w_eco7584, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7585(w_eco7585, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7586(w_eco7586, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7587(w_eco7587, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7588(w_eco7588, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7589(w_eco7589, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7590(w_eco7590, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7591(w_eco7591, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7592(w_eco7592, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7593(w_eco7593, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7594(w_eco7594, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7595(w_eco7595, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7596(w_eco7596, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7597(w_eco7597, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7598(w_eco7598, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7599(w_eco7599, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7600(w_eco7600, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7601(w_eco7601, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7602(w_eco7602, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7603(w_eco7603, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7604(w_eco7604, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7605(w_eco7605, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7606(w_eco7606, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7607(w_eco7607, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7608(w_eco7608, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7609(w_eco7609, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7610(w_eco7610, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7611(w_eco7611, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7612(w_eco7612, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7613(w_eco7613, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7614(w_eco7614, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7615(w_eco7615, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7616(w_eco7616, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7617(w_eco7617, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7618(w_eco7618, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7619(w_eco7619, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7620(w_eco7620, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7621(w_eco7621, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7622(w_eco7622, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7623(w_eco7623, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7624(w_eco7624, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7625(w_eco7625, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7626(w_eco7626, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7627(w_eco7627, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7628(w_eco7628, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7629(w_eco7629, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7630(w_eco7630, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7631(w_eco7631, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7632(w_eco7632, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7633(w_eco7633, prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7634(w_eco7634, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7635(w_eco7635, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7636(w_eco7636, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7637(w_eco7637, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7638(w_eco7638, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7639(w_eco7639, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7640(w_eco7640, prev_cnt[0], prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7641(w_eco7641, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7642(w_eco7642, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7643(w_eco7643, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7644(w_eco7644, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7645(w_eco7645, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7646(w_eco7646, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7647(w_eco7647, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7648(w_eco7648, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7649(w_eco7649, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7650(w_eco7650, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7651(w_eco7651, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7652(w_eco7652, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7653(w_eco7653, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7654(w_eco7654, Tsync[4], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7655(w_eco7655, Tsync[4], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7656(w_eco7656, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7657(w_eco7657, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7658(w_eco7658, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7659(w_eco7659, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7660(w_eco7660, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7661(w_eco7661, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7662(w_eco7662, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7663(w_eco7663, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7664(w_eco7664, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7665(w_eco7665, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7666(w_eco7666, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7667(w_eco7667, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7668(w_eco7668, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7669(w_eco7669, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7670(w_eco7670, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7671(w_eco7671, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7672(w_eco7672, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7673(w_eco7673, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7674(w_eco7674, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7675(w_eco7675, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7676(w_eco7676, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7677(w_eco7677, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7678(w_eco7678, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7679(w_eco7679, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7680(w_eco7680, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7681(w_eco7681, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7682(w_eco7682, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7683(w_eco7683, Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7684(w_eco7684, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7685(w_eco7685, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7686(w_eco7686, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7687(w_eco7687, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7688(w_eco7688, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7689(w_eco7689, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7690(w_eco7690, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7691(w_eco7691, !Tgate[3], !Tsync[3], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7692(w_eco7692, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7693(w_eco7693, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7694(w_eco7694, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7695(w_eco7695, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7696(w_eco7696, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7697(w_eco7697, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7698(w_eco7698, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7699(w_eco7699, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7700(w_eco7700, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7701(w_eco7701, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7702(w_eco7702, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7703(w_eco7703, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7704(w_eco7704, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7705(w_eco7705, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7706(w_eco7706, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7707(w_eco7707, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7708(w_eco7708, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7709(w_eco7709, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7710(w_eco7710, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7711(w_eco7711, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7712(w_eco7712, !Tgate[3], !Tgdel[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7713(w_eco7713, prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7714(w_eco7714, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7715(w_eco7715, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7716(w_eco7716, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7717(w_eco7717, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7718(w_eco7718, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7719(w_eco7719, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7720(w_eco7720, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7721(w_eco7721, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7722(w_eco7722, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7723(w_eco7723, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7724(w_eco7724, Tsync[4], !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7725(w_eco7725, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7726(w_eco7726, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7727(w_eco7727, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7728(w_eco7728, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7729(w_eco7729, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7730(w_eco7730, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7731(w_eco7731, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7732(w_eco7732, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7733(w_eco7733, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7734(w_eco7734, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7735(w_eco7735, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7736(w_eco7736, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7737(w_eco7737, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7738(w_eco7738, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7739(w_eco7739, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7740(w_eco7740, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7741(w_eco7741, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7742(w_eco7742, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7743(w_eco7743, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7744(w_eco7744, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7745(w_eco7745, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[1], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7746(w_eco7746, Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7747(w_eco7747, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7748(w_eco7748, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7749(w_eco7749, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7750(w_eco7750, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7751(w_eco7751, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7752(w_eco7752, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7753(w_eco7753, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7754(w_eco7754, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7755(w_eco7755, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7756(w_eco7756, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7757(w_eco7757, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7758(w_eco7758, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7759(w_eco7759, !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7760(w_eco7760, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7761(w_eco7761, !Tgate[3], !Tgdel[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7762(w_eco7762, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7763(w_eco7763, prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7764(w_eco7764, Tsync[4], Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7765(w_eco7765, Tsync[4], Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7766(w_eco7766, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7767(w_eco7767, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7768(w_eco7768, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7769(w_eco7769, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7770(w_eco7770, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7771(w_eco7771, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7772(w_eco7772, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7773(w_eco7773, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7774(w_eco7774, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_7775(w_eco7775, Tsync[3], !prev_cnt[14], prev_cnt[1], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7776(w_eco7776, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7777(w_eco7777, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[2], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7778(w_eco7778, Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7779(w_eco7779, Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7780(w_eco7780, !Tgate[3], !Tsync[3], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_7781(w_eco7781, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7782(w_eco7782, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7783(w_eco7783, !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7784(w_eco7784, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7785(w_eco7785, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7786(w_eco7786, !Tgate[3], !Tgdel[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7787(w_eco7787, !Tgate[3], !Tgdel[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7788(w_eco7788, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7789(w_eco7789, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7790(w_eco7790, Tsync[3], !prev_cnt[14], prev_cnt[2], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7791(w_eco7791, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7792(w_eco7792, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7793(w_eco7793, !Tgate[3], !Tgdel[3], Tsync[3], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7794(w_eco7794, !Tgate[3], !Tgdel[3], Tsync[3], prev_cnt[0], !prev_cnt[3], prev_cnt[4], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7795(w_eco7795, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7796(w_eco7796, !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7797(w_eco7797, Tsync[3], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_7798(w_eco7798, Tsync[3], !prev_cnt[14], prev_cnt[0], !prev_cnt[3], prev_cnt[4], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_7799(w_eco7799, w_eco5481, w_eco5482, w_eco5483, w_eco5484, w_eco5485, w_eco5486, w_eco5487, w_eco5488, w_eco5489, w_eco5490, w_eco5491, w_eco5492, w_eco5493, w_eco5494, w_eco5495, w_eco5496, w_eco5497, w_eco5498, w_eco5499, w_eco5500, w_eco5501, w_eco5502, w_eco5503, w_eco5504, w_eco5505, w_eco5506, w_eco5507, w_eco5508, w_eco5509, w_eco5510, w_eco5511, w_eco5512, w_eco5513, w_eco5514, w_eco5515, w_eco5516, w_eco5517, w_eco5518, w_eco5519, w_eco5520, w_eco5521, w_eco5522, w_eco5523, w_eco5524, w_eco5525, w_eco5526, w_eco5527, w_eco5528, w_eco5529, w_eco5530, w_eco5531, w_eco5532, w_eco5533, w_eco5534, w_eco5535, w_eco5536, w_eco5537, w_eco5538, w_eco5539, w_eco5540, w_eco5541, w_eco5542, w_eco5543, w_eco5544, w_eco5545, w_eco5546, w_eco5547, w_eco5548, w_eco5549, w_eco5550, w_eco5551, w_eco5552, w_eco5553, w_eco5554, w_eco5555, w_eco5556, w_eco5557, w_eco5558, w_eco5559, w_eco5560, w_eco5561, w_eco5562, w_eco5563, w_eco5564, w_eco5565, w_eco5566, w_eco5567, w_eco5568, w_eco5569, w_eco5570, w_eco5571, w_eco5572, w_eco5573, w_eco5574, w_eco5575, w_eco5576, w_eco5577, w_eco5578, w_eco5579, w_eco5580, w_eco5581, w_eco5582, w_eco5583, w_eco5584, w_eco5585, w_eco5586, w_eco5587, w_eco5588, w_eco5589, w_eco5590, w_eco5591, w_eco5592, w_eco5593, w_eco5594, w_eco5595, w_eco5596, w_eco5597, w_eco5598, w_eco5599, w_eco5600, w_eco5601, w_eco5602, w_eco5603, w_eco5604, w_eco5605, w_eco5606, w_eco5607, w_eco5608, w_eco5609, w_eco5610, w_eco5611, w_eco5612, w_eco5613, w_eco5614, w_eco5615, w_eco5616, w_eco5617, w_eco5618, w_eco5619, w_eco5620, w_eco5621, w_eco5622, w_eco5623, w_eco5624, w_eco5625, w_eco5626, w_eco5627, w_eco5628, w_eco5629, w_eco5630, w_eco5631, w_eco5632, w_eco5633, w_eco5634, w_eco5635, w_eco5636, w_eco5637, w_eco5638, w_eco5639, w_eco5640, w_eco5641, w_eco5642, w_eco5643, w_eco5644, w_eco5645, w_eco5646, w_eco5647, w_eco5648, w_eco5649, w_eco5650, w_eco5651, w_eco5652, w_eco5653, w_eco5654, w_eco5655, w_eco5656, w_eco5657, w_eco5658, w_eco5659, w_eco5660, w_eco5661, w_eco5662, w_eco5663, w_eco5664, w_eco5665, w_eco5666, w_eco5667, w_eco5668, w_eco5669, w_eco5670, w_eco5671, w_eco5672, w_eco5673, w_eco5674, w_eco5675, w_eco5676, w_eco5677, w_eco5678, w_eco5679, w_eco5680, w_eco5681, w_eco5682, w_eco5683, w_eco5684, w_eco5685, w_eco5686, w_eco5687, w_eco5688, w_eco5689, w_eco5690, w_eco5691, w_eco5692, w_eco5693, w_eco5694, w_eco5695, w_eco5696, w_eco5697, w_eco5698, w_eco5699, w_eco5700, w_eco5701, w_eco5702, w_eco5703, w_eco5704, w_eco5705, w_eco5706, w_eco5707, w_eco5708, w_eco5709, w_eco5710, w_eco5711, w_eco5712, w_eco5713, w_eco5714, w_eco5715, w_eco5716, w_eco5717, w_eco5718, w_eco5719, w_eco5720, w_eco5721, w_eco5722, w_eco5723, w_eco5724, w_eco5725, w_eco5726, w_eco5727, w_eco5728, w_eco5729, w_eco5730, w_eco5731, w_eco5732, w_eco5733, w_eco5734, w_eco5735, w_eco5736, w_eco5737, w_eco5738, w_eco5739, w_eco5740, w_eco5741, w_eco5742, w_eco5743, w_eco5744, w_eco5745, w_eco5746, w_eco5747, w_eco5748, w_eco5749, w_eco5750, w_eco5751, w_eco5752, w_eco5753, w_eco5754, w_eco5755, w_eco5756, w_eco5757, w_eco5758, w_eco5759, w_eco5760, w_eco5761, w_eco5762, w_eco5763, w_eco5764, w_eco5765, w_eco5766, w_eco5767, w_eco5768, w_eco5769, w_eco5770, w_eco5771, w_eco5772, w_eco5773, w_eco5774, w_eco5775, w_eco5776, w_eco5777, w_eco5778, w_eco5779, w_eco5780, w_eco5781, w_eco5782, w_eco5783, w_eco5784, w_eco5785, w_eco5786, w_eco5787, w_eco5788, w_eco5789, w_eco5790, w_eco5791, w_eco5792, w_eco5793, w_eco5794, w_eco5795, w_eco5796, w_eco5797, w_eco5798, w_eco5799, w_eco5800, w_eco5801, w_eco5802, w_eco5803, w_eco5804, w_eco5805, w_eco5806, w_eco5807, w_eco5808, w_eco5809, w_eco5810, w_eco5811, w_eco5812, w_eco5813, w_eco5814, w_eco5815, w_eco5816, w_eco5817, w_eco5818, w_eco5819, w_eco5820, w_eco5821, w_eco5822, w_eco5823, w_eco5824, w_eco5825, w_eco5826, w_eco5827, w_eco5828, w_eco5829, w_eco5830, w_eco5831, w_eco5832, w_eco5833, w_eco5834, w_eco5835, w_eco5836, w_eco5837, w_eco5838, w_eco5839, w_eco5840, w_eco5841, w_eco5842, w_eco5843, w_eco5844, w_eco5845, w_eco5846, w_eco5847, w_eco5848, w_eco5849, w_eco5850, w_eco5851, w_eco5852, w_eco5853, w_eco5854, w_eco5855, w_eco5856, w_eco5857, w_eco5858, w_eco5859, w_eco5860, w_eco5861, w_eco5862, w_eco5863, w_eco5864, w_eco5865, w_eco5866, w_eco5867, w_eco5868, w_eco5869, w_eco5870, w_eco5871, w_eco5872, w_eco5873, w_eco5874, w_eco5875, w_eco5876, w_eco5877, w_eco5878, w_eco5879, w_eco5880, w_eco5881, w_eco5882, w_eco5883, w_eco5884, w_eco5885, w_eco5886, w_eco5887, w_eco5888, w_eco5889, w_eco5890, w_eco5891, w_eco5892, w_eco5893, w_eco5894, w_eco5895, w_eco5896, w_eco5897, w_eco5898, w_eco5899, w_eco5900, w_eco5901, w_eco5902, w_eco5903, w_eco5904, w_eco5905, w_eco5906, w_eco5907, w_eco5908, w_eco5909, w_eco5910, w_eco5911, w_eco5912, w_eco5913, w_eco5914, w_eco5915, w_eco5916, w_eco5917, w_eco5918, w_eco5919, w_eco5920, w_eco5921, w_eco5922, w_eco5923, w_eco5924, w_eco5925, w_eco5926, w_eco5927, w_eco5928, w_eco5929, w_eco5930, w_eco5931, w_eco5932, w_eco5933, w_eco5934, w_eco5935, w_eco5936, w_eco5937, w_eco5938, w_eco5939, w_eco5940, w_eco5941, w_eco5942, w_eco5943, w_eco5944, w_eco5945, w_eco5946, w_eco5947, w_eco5948, w_eco5949, w_eco5950, w_eco5951, w_eco5952, w_eco5953, w_eco5954, w_eco5955, w_eco5956, w_eco5957, w_eco5958, w_eco5959, w_eco5960, w_eco5961, w_eco5962, w_eco5963, w_eco5964, w_eco5965, w_eco5966, w_eco5967, w_eco5968, w_eco5969, w_eco5970, w_eco5971, w_eco5972, w_eco5973, w_eco5974, w_eco5975, w_eco5976, w_eco5977, w_eco5978, w_eco5979, w_eco5980, w_eco5981, w_eco5982, w_eco5983, w_eco5984, w_eco5985, w_eco5986, w_eco5987, w_eco5988, w_eco5989, w_eco5990, w_eco5991, w_eco5992, w_eco5993, w_eco5994, w_eco5995, w_eco5996, w_eco5997, w_eco5998, w_eco5999, w_eco6000, w_eco6001, w_eco6002, w_eco6003, w_eco6004, w_eco6005, w_eco6006, w_eco6007, w_eco6008, w_eco6009, w_eco6010, w_eco6011, w_eco6012, w_eco6013, w_eco6014, w_eco6015, w_eco6016, w_eco6017, w_eco6018, w_eco6019, w_eco6020, w_eco6021, w_eco6022, w_eco6023, w_eco6024, w_eco6025, w_eco6026, w_eco6027, w_eco6028, w_eco6029, w_eco6030, w_eco6031, w_eco6032, w_eco6033, w_eco6034, w_eco6035, w_eco6036, w_eco6037, w_eco6038, w_eco6039, w_eco6040, w_eco6041, w_eco6042, w_eco6043, w_eco6044, w_eco6045, w_eco6046, w_eco6047, w_eco6048, w_eco6049, w_eco6050, w_eco6051, w_eco6052, w_eco6053, w_eco6054, w_eco6055, w_eco6056, w_eco6057, w_eco6058, w_eco6059, w_eco6060, w_eco6061, w_eco6062, w_eco6063, w_eco6064, w_eco6065, w_eco6066, w_eco6067, w_eco6068, w_eco6069, w_eco6070, w_eco6071, w_eco6072, w_eco6073, w_eco6074, w_eco6075, w_eco6076, w_eco6077, w_eco6078, w_eco6079, w_eco6080, w_eco6081, w_eco6082, w_eco6083, w_eco6084, w_eco6085, w_eco6086, w_eco6087, w_eco6088, w_eco6089, w_eco6090, w_eco6091, w_eco6092, w_eco6093, w_eco6094, w_eco6095, w_eco6096, w_eco6097, w_eco6098, w_eco6099, w_eco6100, w_eco6101, w_eco6102, w_eco6103, w_eco6104, w_eco6105, w_eco6106, w_eco6107, w_eco6108, w_eco6109, w_eco6110, w_eco6111, w_eco6112, w_eco6113, w_eco6114, w_eco6115, w_eco6116, w_eco6117, w_eco6118, w_eco6119, w_eco6120, w_eco6121, w_eco6122, w_eco6123, w_eco6124, w_eco6125, w_eco6126, w_eco6127, w_eco6128, w_eco6129, w_eco6130, w_eco6131, w_eco6132, w_eco6133, w_eco6134, w_eco6135, w_eco6136, w_eco6137, w_eco6138, w_eco6139, w_eco6140, w_eco6141, w_eco6142, w_eco6143, w_eco6144, w_eco6145, w_eco6146, w_eco6147, w_eco6148, w_eco6149, w_eco6150, w_eco6151, w_eco6152, w_eco6153, w_eco6154, w_eco6155, w_eco6156, w_eco6157, w_eco6158, w_eco6159, w_eco6160, w_eco6161, w_eco6162, w_eco6163, w_eco6164, w_eco6165, w_eco6166, w_eco6167, w_eco6168, w_eco6169, w_eco6170, w_eco6171, w_eco6172, w_eco6173, w_eco6174, w_eco6175, w_eco6176, w_eco6177, w_eco6178, w_eco6179, w_eco6180, w_eco6181, w_eco6182, w_eco6183, w_eco6184, w_eco6185, w_eco6186, w_eco6187, w_eco6188, w_eco6189, w_eco6190, w_eco6191, w_eco6192, w_eco6193, w_eco6194, w_eco6195, w_eco6196, w_eco6197, w_eco6198, w_eco6199, w_eco6200, w_eco6201, w_eco6202, w_eco6203, w_eco6204, w_eco6205, w_eco6206, w_eco6207, w_eco6208, w_eco6209, w_eco6210, w_eco6211, w_eco6212, w_eco6213, w_eco6214, w_eco6215, w_eco6216, w_eco6217, w_eco6218, w_eco6219, w_eco6220, w_eco6221, w_eco6222, w_eco6223, w_eco6224, w_eco6225, w_eco6226, w_eco6227, w_eco6228, w_eco6229, w_eco6230, w_eco6231, w_eco6232, w_eco6233, w_eco6234, w_eco6235, w_eco6236, w_eco6237, w_eco6238, w_eco6239, w_eco6240, w_eco6241, w_eco6242, w_eco6243, w_eco6244, w_eco6245, w_eco6246, w_eco6247, w_eco6248, w_eco6249, w_eco6250, w_eco6251, w_eco6252, w_eco6253, w_eco6254, w_eco6255, w_eco6256, w_eco6257, w_eco6258, w_eco6259, w_eco6260, w_eco6261, w_eco6262, w_eco6263, w_eco6264, w_eco6265, w_eco6266, w_eco6267, w_eco6268, w_eco6269, w_eco6270, w_eco6271, w_eco6272, w_eco6273, w_eco6274, w_eco6275, w_eco6276, w_eco6277, w_eco6278, w_eco6279, w_eco6280, w_eco6281, w_eco6282, w_eco6283, w_eco6284, w_eco6285, w_eco6286, w_eco6287, w_eco6288, w_eco6289, w_eco6290, w_eco6291, w_eco6292, w_eco6293, w_eco6294, w_eco6295, w_eco6296, w_eco6297, w_eco6298, w_eco6299, w_eco6300, w_eco6301, w_eco6302, w_eco6303, w_eco6304, w_eco6305, w_eco6306, w_eco6307, w_eco6308, w_eco6309, w_eco6310, w_eco6311, w_eco6312, w_eco6313, w_eco6314, w_eco6315, w_eco6316, w_eco6317, w_eco6318, w_eco6319, w_eco6320, w_eco6321, w_eco6322, w_eco6323, w_eco6324, w_eco6325, w_eco6326, w_eco6327, w_eco6328, w_eco6329, w_eco6330, w_eco6331, w_eco6332, w_eco6333, w_eco6334, w_eco6335, w_eco6336, w_eco6337, w_eco6338, w_eco6339, w_eco6340, w_eco6341, w_eco6342, w_eco6343, w_eco6344, w_eco6345, w_eco6346, w_eco6347, w_eco6348, w_eco6349, w_eco6350, w_eco6351, w_eco6352, w_eco6353, w_eco6354, w_eco6355, w_eco6356, w_eco6357, w_eco6358, w_eco6359, w_eco6360, w_eco6361, w_eco6362, w_eco6363, w_eco6364, w_eco6365, w_eco6366, w_eco6367, w_eco6368, w_eco6369, w_eco6370, w_eco6371, w_eco6372, w_eco6373, w_eco6374, w_eco6375, w_eco6376, w_eco6377, w_eco6378, w_eco6379, w_eco6380, w_eco6381, w_eco6382, w_eco6383, w_eco6384, w_eco6385, w_eco6386, w_eco6387, w_eco6388, w_eco6389, w_eco6390, w_eco6391, w_eco6392, w_eco6393, w_eco6394, w_eco6395, w_eco6396, w_eco6397, w_eco6398, w_eco6399, w_eco6400, w_eco6401, w_eco6402, w_eco6403, w_eco6404, w_eco6405, w_eco6406, w_eco6407, w_eco6408, w_eco6409, w_eco6410, w_eco6411, w_eco6412, w_eco6413, w_eco6414, w_eco6415, w_eco6416, w_eco6417, w_eco6418, w_eco6419, w_eco6420, w_eco6421, w_eco6422, w_eco6423, w_eco6424, w_eco6425, w_eco6426, w_eco6427, w_eco6428, w_eco6429, w_eco6430, w_eco6431, w_eco6432, w_eco6433, w_eco6434, w_eco6435, w_eco6436, w_eco6437, w_eco6438, w_eco6439, w_eco6440, w_eco6441, w_eco6442, w_eco6443, w_eco6444, w_eco6445, w_eco6446, w_eco6447, w_eco6448, w_eco6449, w_eco6450, w_eco6451, w_eco6452, w_eco6453, w_eco6454, w_eco6455, w_eco6456, w_eco6457, w_eco6458, w_eco6459, w_eco6460, w_eco6461, w_eco6462, w_eco6463, w_eco6464, w_eco6465, w_eco6466, w_eco6467, w_eco6468, w_eco6469, w_eco6470, w_eco6471, w_eco6472, w_eco6473, w_eco6474, w_eco6475, w_eco6476, w_eco6477, w_eco6478, w_eco6479, w_eco6480, w_eco6481, w_eco6482, w_eco6483, w_eco6484, w_eco6485, w_eco6486, w_eco6487, w_eco6488, w_eco6489, w_eco6490, w_eco6491, w_eco6492, w_eco6493, w_eco6494, w_eco6495, w_eco6496, w_eco6497, w_eco6498, w_eco6499, w_eco6500, w_eco6501, w_eco6502, w_eco6503, w_eco6504, w_eco6505, w_eco6506, w_eco6507, w_eco6508, w_eco6509, w_eco6510, w_eco6511, w_eco6512, w_eco6513, w_eco6514, w_eco6515, w_eco6516, w_eco6517, w_eco6518, w_eco6519, w_eco6520, w_eco6521, w_eco6522, w_eco6523, w_eco6524, w_eco6525, w_eco6526, w_eco6527, w_eco6528, w_eco6529, w_eco6530, w_eco6531, w_eco6532, w_eco6533, w_eco6534, w_eco6535, w_eco6536, w_eco6537, w_eco6538, w_eco6539, w_eco6540, w_eco6541, w_eco6542, w_eco6543, w_eco6544, w_eco6545, w_eco6546, w_eco6547, w_eco6548, w_eco6549, w_eco6550, w_eco6551, w_eco6552, w_eco6553, w_eco6554, w_eco6555, w_eco6556, w_eco6557, w_eco6558, w_eco6559, w_eco6560, w_eco6561, w_eco6562, w_eco6563, w_eco6564, w_eco6565, w_eco6566, w_eco6567, w_eco6568, w_eco6569, w_eco6570, w_eco6571, w_eco6572, w_eco6573, w_eco6574, w_eco6575, w_eco6576, w_eco6577, w_eco6578, w_eco6579, w_eco6580, w_eco6581, w_eco6582, w_eco6583, w_eco6584, w_eco6585, w_eco6586, w_eco6587, w_eco6588, w_eco6589, w_eco6590, w_eco6591, w_eco6592, w_eco6593, w_eco6594, w_eco6595, w_eco6596, w_eco6597, w_eco6598, w_eco6599, w_eco6600, w_eco6601, w_eco6602, w_eco6603, w_eco6604, w_eco6605, w_eco6606, w_eco6607, w_eco6608, w_eco6609, w_eco6610, w_eco6611, w_eco6612, w_eco6613, w_eco6614, w_eco6615, w_eco6616, w_eco6617, w_eco6618, w_eco6619, w_eco6620, w_eco6621, w_eco6622, w_eco6623, w_eco6624, w_eco6625, w_eco6626, w_eco6627, w_eco6628, w_eco6629, w_eco6630, w_eco6631, w_eco6632, w_eco6633, w_eco6634, w_eco6635, w_eco6636, w_eco6637, w_eco6638, w_eco6639, w_eco6640, w_eco6641, w_eco6642, w_eco6643, w_eco6644, w_eco6645, w_eco6646, w_eco6647, w_eco6648, w_eco6649, w_eco6650, w_eco6651, w_eco6652, w_eco6653, w_eco6654, w_eco6655, w_eco6656, w_eco6657, w_eco6658, w_eco6659, w_eco6660, w_eco6661, w_eco6662, w_eco6663, w_eco6664, w_eco6665, w_eco6666, w_eco6667, w_eco6668, w_eco6669, w_eco6670, w_eco6671, w_eco6672, w_eco6673, w_eco6674, w_eco6675, w_eco6676, w_eco6677, w_eco6678, w_eco6679, w_eco6680, w_eco6681, w_eco6682, w_eco6683, w_eco6684, w_eco6685, w_eco6686, w_eco6687, w_eco6688, w_eco6689, w_eco6690, w_eco6691, w_eco6692, w_eco6693, w_eco6694, w_eco6695, w_eco6696, w_eco6697, w_eco6698, w_eco6699, w_eco6700, w_eco6701, w_eco6702, w_eco6703, w_eco6704, w_eco6705, w_eco6706, w_eco6707, w_eco6708, w_eco6709, w_eco6710, w_eco6711, w_eco6712, w_eco6713, w_eco6714, w_eco6715, w_eco6716, w_eco6717, w_eco6718, w_eco6719, w_eco6720, w_eco6721, w_eco6722, w_eco6723, w_eco6724, w_eco6725, w_eco6726, w_eco6727, w_eco6728, w_eco6729, w_eco6730, w_eco6731, w_eco6732, w_eco6733, w_eco6734, w_eco6735, w_eco6736, w_eco6737, w_eco6738, w_eco6739, w_eco6740, w_eco6741, w_eco6742, w_eco6743, w_eco6744, w_eco6745, w_eco6746, w_eco6747, w_eco6748, w_eco6749, w_eco6750, w_eco6751, w_eco6752, w_eco6753, w_eco6754, w_eco6755, w_eco6756, w_eco6757, w_eco6758, w_eco6759, w_eco6760, w_eco6761, w_eco6762, w_eco6763, w_eco6764, w_eco6765, w_eco6766, w_eco6767, w_eco6768, w_eco6769, w_eco6770, w_eco6771, w_eco6772, w_eco6773, w_eco6774, w_eco6775, w_eco6776, w_eco6777, w_eco6778, w_eco6779, w_eco6780, w_eco6781, w_eco6782, w_eco6783, w_eco6784, w_eco6785, w_eco6786, w_eco6787, w_eco6788, w_eco6789, w_eco6790, w_eco6791, w_eco6792, w_eco6793, w_eco6794, w_eco6795, w_eco6796, w_eco6797, w_eco6798, w_eco6799, w_eco6800, w_eco6801, w_eco6802, w_eco6803, w_eco6804, w_eco6805, w_eco6806, w_eco6807, w_eco6808, w_eco6809, w_eco6810, w_eco6811, w_eco6812, w_eco6813, w_eco6814, w_eco6815, w_eco6816, w_eco6817, w_eco6818, w_eco6819, w_eco6820, w_eco6821, w_eco6822, w_eco6823, w_eco6824, w_eco6825, w_eco6826, w_eco6827, w_eco6828, w_eco6829, w_eco6830, w_eco6831, w_eco6832, w_eco6833, w_eco6834, w_eco6835, w_eco6836, w_eco6837, w_eco6838, w_eco6839, w_eco6840, w_eco6841, w_eco6842, w_eco6843, w_eco6844, w_eco6845, w_eco6846, w_eco6847, w_eco6848, w_eco6849, w_eco6850, w_eco6851, w_eco6852, w_eco6853, w_eco6854, w_eco6855, w_eco6856, w_eco6857, w_eco6858, w_eco6859, w_eco6860, w_eco6861, w_eco6862, w_eco6863, w_eco6864, w_eco6865, w_eco6866, w_eco6867, w_eco6868, w_eco6869, w_eco6870, w_eco6871, w_eco6872, w_eco6873, w_eco6874, w_eco6875, w_eco6876, w_eco6877, w_eco6878, w_eco6879, w_eco6880, w_eco6881, w_eco6882, w_eco6883, w_eco6884, w_eco6885, w_eco6886, w_eco6887, w_eco6888, w_eco6889, w_eco6890, w_eco6891, w_eco6892, w_eco6893, w_eco6894, w_eco6895, w_eco6896, w_eco6897, w_eco6898, w_eco6899, w_eco6900, w_eco6901, w_eco6902, w_eco6903, w_eco6904, w_eco6905, w_eco6906, w_eco6907, w_eco6908, w_eco6909, w_eco6910, w_eco6911, w_eco6912, w_eco6913, w_eco6914, w_eco6915, w_eco6916, w_eco6917, w_eco6918, w_eco6919, w_eco6920, w_eco6921, w_eco6922, w_eco6923, w_eco6924, w_eco6925, w_eco6926, w_eco6927, w_eco6928, w_eco6929, w_eco6930, w_eco6931, w_eco6932, w_eco6933, w_eco6934, w_eco6935, w_eco6936, w_eco6937, w_eco6938, w_eco6939, w_eco6940, w_eco6941, w_eco6942, w_eco6943, w_eco6944, w_eco6945, w_eco6946, w_eco6947, w_eco6948, w_eco6949, w_eco6950, w_eco6951, w_eco6952, w_eco6953, w_eco6954, w_eco6955, w_eco6956, w_eco6957, w_eco6958, w_eco6959, w_eco6960, w_eco6961, w_eco6962, w_eco6963, w_eco6964, w_eco6965, w_eco6966, w_eco6967, w_eco6968, w_eco6969, w_eco6970, w_eco6971, w_eco6972, w_eco6973, w_eco6974, w_eco6975, w_eco6976, w_eco6977, w_eco6978, w_eco6979, w_eco6980, w_eco6981, w_eco6982, w_eco6983, w_eco6984, w_eco6985, w_eco6986, w_eco6987, w_eco6988, w_eco6989, w_eco6990, w_eco6991, w_eco6992, w_eco6993, w_eco6994, w_eco6995, w_eco6996, w_eco6997, w_eco6998, w_eco6999, w_eco7000, w_eco7001, w_eco7002, w_eco7003, w_eco7004, w_eco7005, w_eco7006, w_eco7007, w_eco7008, w_eco7009, w_eco7010, w_eco7011, w_eco7012, w_eco7013, w_eco7014, w_eco7015, w_eco7016, w_eco7017, w_eco7018, w_eco7019, w_eco7020, w_eco7021, w_eco7022, w_eco7023, w_eco7024, w_eco7025, w_eco7026, w_eco7027, w_eco7028, w_eco7029, w_eco7030, w_eco7031, w_eco7032, w_eco7033, w_eco7034, w_eco7035, w_eco7036, w_eco7037, w_eco7038, w_eco7039, w_eco7040, w_eco7041, w_eco7042, w_eco7043, w_eco7044, w_eco7045, w_eco7046, w_eco7047, w_eco7048, w_eco7049, w_eco7050, w_eco7051, w_eco7052, w_eco7053, w_eco7054, w_eco7055, w_eco7056, w_eco7057, w_eco7058, w_eco7059, w_eco7060, w_eco7061, w_eco7062, w_eco7063, w_eco7064, w_eco7065, w_eco7066, w_eco7067, w_eco7068, w_eco7069, w_eco7070, w_eco7071, w_eco7072, w_eco7073, w_eco7074, w_eco7075, w_eco7076, w_eco7077, w_eco7078, w_eco7079, w_eco7080, w_eco7081, w_eco7082, w_eco7083, w_eco7084, w_eco7085, w_eco7086, w_eco7087, w_eco7088, w_eco7089, w_eco7090, w_eco7091, w_eco7092, w_eco7093, w_eco7094, w_eco7095, w_eco7096, w_eco7097, w_eco7098, w_eco7099, w_eco7100, w_eco7101, w_eco7102, w_eco7103, w_eco7104, w_eco7105, w_eco7106, w_eco7107, w_eco7108, w_eco7109, w_eco7110, w_eco7111, w_eco7112, w_eco7113, w_eco7114, w_eco7115, w_eco7116, w_eco7117, w_eco7118, w_eco7119, w_eco7120, w_eco7121, w_eco7122, w_eco7123, w_eco7124, w_eco7125, w_eco7126, w_eco7127, w_eco7128, w_eco7129, w_eco7130, w_eco7131, w_eco7132, w_eco7133, w_eco7134, w_eco7135, w_eco7136, w_eco7137, w_eco7138, w_eco7139, w_eco7140, w_eco7141, w_eco7142, w_eco7143, w_eco7144, w_eco7145, w_eco7146, w_eco7147, w_eco7148, w_eco7149, w_eco7150, w_eco7151, w_eco7152, w_eco7153, w_eco7154, w_eco7155, w_eco7156, w_eco7157, w_eco7158, w_eco7159, w_eco7160, w_eco7161, w_eco7162, w_eco7163, w_eco7164, w_eco7165, w_eco7166, w_eco7167, w_eco7168, w_eco7169, w_eco7170, w_eco7171, w_eco7172, w_eco7173, w_eco7174, w_eco7175, w_eco7176, w_eco7177, w_eco7178, w_eco7179, w_eco7180, w_eco7181, w_eco7182, w_eco7183, w_eco7184, w_eco7185, w_eco7186, w_eco7187, w_eco7188, w_eco7189, w_eco7190, w_eco7191, w_eco7192, w_eco7193, w_eco7194, w_eco7195, w_eco7196, w_eco7197, w_eco7198, w_eco7199, w_eco7200, w_eco7201, w_eco7202, w_eco7203, w_eco7204, w_eco7205, w_eco7206, w_eco7207, w_eco7208, w_eco7209, w_eco7210, w_eco7211, w_eco7212, w_eco7213, w_eco7214, w_eco7215, w_eco7216, w_eco7217, w_eco7218, w_eco7219, w_eco7220, w_eco7221, w_eco7222, w_eco7223, w_eco7224, w_eco7225, w_eco7226, w_eco7227, w_eco7228, w_eco7229, w_eco7230, w_eco7231, w_eco7232, w_eco7233, w_eco7234, w_eco7235, w_eco7236, w_eco7237, w_eco7238, w_eco7239, w_eco7240, w_eco7241, w_eco7242, w_eco7243, w_eco7244, w_eco7245, w_eco7246, w_eco7247, w_eco7248, w_eco7249, w_eco7250, w_eco7251, w_eco7252, w_eco7253, w_eco7254, w_eco7255, w_eco7256, w_eco7257, w_eco7258, w_eco7259, w_eco7260, w_eco7261, w_eco7262, w_eco7263, w_eco7264, w_eco7265, w_eco7266, w_eco7267, w_eco7268, w_eco7269, w_eco7270, w_eco7271, w_eco7272, w_eco7273, w_eco7274, w_eco7275, w_eco7276, w_eco7277, w_eco7278, w_eco7279, w_eco7280, w_eco7281, w_eco7282, w_eco7283, w_eco7284, w_eco7285, w_eco7286, w_eco7287, w_eco7288, w_eco7289, w_eco7290, w_eco7291, w_eco7292, w_eco7293, w_eco7294, w_eco7295, w_eco7296, w_eco7297, w_eco7298, w_eco7299, w_eco7300, w_eco7301, w_eco7302, w_eco7303, w_eco7304, w_eco7305, w_eco7306, w_eco7307, w_eco7308, w_eco7309, w_eco7310, w_eco7311, w_eco7312, w_eco7313, w_eco7314, w_eco7315, w_eco7316, w_eco7317, w_eco7318, w_eco7319, w_eco7320, w_eco7321, w_eco7322, w_eco7323, w_eco7324, w_eco7325, w_eco7326, w_eco7327, w_eco7328, w_eco7329, w_eco7330, w_eco7331, w_eco7332, w_eco7333, w_eco7334, w_eco7335, w_eco7336, w_eco7337, w_eco7338, w_eco7339, w_eco7340, w_eco7341, w_eco7342, w_eco7343, w_eco7344, w_eco7345, w_eco7346, w_eco7347, w_eco7348, w_eco7349, w_eco7350, w_eco7351, w_eco7352, w_eco7353, w_eco7354, w_eco7355, w_eco7356, w_eco7357, w_eco7358, w_eco7359, w_eco7360, w_eco7361, w_eco7362, w_eco7363, w_eco7364, w_eco7365, w_eco7366, w_eco7367, w_eco7368, w_eco7369, w_eco7370, w_eco7371, w_eco7372, w_eco7373, w_eco7374, w_eco7375, w_eco7376, w_eco7377, w_eco7378, w_eco7379, w_eco7380, w_eco7381, w_eco7382, w_eco7383, w_eco7384, w_eco7385, w_eco7386, w_eco7387, w_eco7388, w_eco7389, w_eco7390, w_eco7391, w_eco7392, w_eco7393, w_eco7394, w_eco7395, w_eco7396, w_eco7397, w_eco7398, w_eco7399, w_eco7400, w_eco7401, w_eco7402, w_eco7403, w_eco7404, w_eco7405, w_eco7406, w_eco7407, w_eco7408, w_eco7409, w_eco7410, w_eco7411, w_eco7412, w_eco7413, w_eco7414, w_eco7415, w_eco7416, w_eco7417, w_eco7418, w_eco7419, w_eco7420, w_eco7421, w_eco7422, w_eco7423, w_eco7424, w_eco7425, w_eco7426, w_eco7427, w_eco7428, w_eco7429, w_eco7430, w_eco7431, w_eco7432, w_eco7433, w_eco7434, w_eco7435, w_eco7436, w_eco7437, w_eco7438, w_eco7439, w_eco7440, w_eco7441, w_eco7442, w_eco7443, w_eco7444, w_eco7445, w_eco7446, w_eco7447, w_eco7448, w_eco7449, w_eco7450, w_eco7451, w_eco7452, w_eco7453, w_eco7454, w_eco7455, w_eco7456, w_eco7457, w_eco7458, w_eco7459, w_eco7460, w_eco7461, w_eco7462, w_eco7463, w_eco7464, w_eco7465, w_eco7466, w_eco7467, w_eco7468, w_eco7469, w_eco7470, w_eco7471, w_eco7472, w_eco7473, w_eco7474, w_eco7475, w_eco7476, w_eco7477, w_eco7478, w_eco7479, w_eco7480, w_eco7481, w_eco7482, w_eco7483, w_eco7484, w_eco7485, w_eco7486, w_eco7487, w_eco7488, w_eco7489, w_eco7490, w_eco7491, w_eco7492, w_eco7493, w_eco7494, w_eco7495, w_eco7496, w_eco7497, w_eco7498, w_eco7499, w_eco7500, w_eco7501, w_eco7502, w_eco7503, w_eco7504, w_eco7505, w_eco7506, w_eco7507, w_eco7508, w_eco7509, w_eco7510, w_eco7511, w_eco7512, w_eco7513, w_eco7514, w_eco7515, w_eco7516, w_eco7517, w_eco7518, w_eco7519, w_eco7520, w_eco7521, w_eco7522, w_eco7523, w_eco7524, w_eco7525, w_eco7526, w_eco7527, w_eco7528, w_eco7529, w_eco7530, w_eco7531, w_eco7532, w_eco7533, w_eco7534, w_eco7535, w_eco7536, w_eco7537, w_eco7538, w_eco7539, w_eco7540, w_eco7541, w_eco7542, w_eco7543, w_eco7544, w_eco7545, w_eco7546, w_eco7547, w_eco7548, w_eco7549, w_eco7550, w_eco7551, w_eco7552, w_eco7553, w_eco7554, w_eco7555, w_eco7556, w_eco7557, w_eco7558, w_eco7559, w_eco7560, w_eco7561, w_eco7562, w_eco7563, w_eco7564, w_eco7565, w_eco7566, w_eco7567, w_eco7568, w_eco7569, w_eco7570, w_eco7571, w_eco7572, w_eco7573, w_eco7574, w_eco7575, w_eco7576, w_eco7577, w_eco7578, w_eco7579, w_eco7580, w_eco7581, w_eco7582, w_eco7583, w_eco7584, w_eco7585, w_eco7586, w_eco7587, w_eco7588, w_eco7589, w_eco7590, w_eco7591, w_eco7592, w_eco7593, w_eco7594, w_eco7595, w_eco7596, w_eco7597, w_eco7598, w_eco7599, w_eco7600, w_eco7601, w_eco7602, w_eco7603, w_eco7604, w_eco7605, w_eco7606, w_eco7607, w_eco7608, w_eco7609, w_eco7610, w_eco7611, w_eco7612, w_eco7613, w_eco7614, w_eco7615, w_eco7616, w_eco7617, w_eco7618, w_eco7619, w_eco7620, w_eco7621, w_eco7622, w_eco7623, w_eco7624, w_eco7625, w_eco7626, w_eco7627, w_eco7628, w_eco7629, w_eco7630, w_eco7631, w_eco7632, w_eco7633, w_eco7634, w_eco7635, w_eco7636, w_eco7637, w_eco7638, w_eco7639, w_eco7640, w_eco7641, w_eco7642, w_eco7643, w_eco7644, w_eco7645, w_eco7646, w_eco7647, w_eco7648, w_eco7649, w_eco7650, w_eco7651, w_eco7652, w_eco7653, w_eco7654, w_eco7655, w_eco7656, w_eco7657, w_eco7658, w_eco7659, w_eco7660, w_eco7661, w_eco7662, w_eco7663, w_eco7664, w_eco7665, w_eco7666, w_eco7667, w_eco7668, w_eco7669, w_eco7670, w_eco7671, w_eco7672, w_eco7673, w_eco7674, w_eco7675, w_eco7676, w_eco7677, w_eco7678, w_eco7679, w_eco7680, w_eco7681, w_eco7682, w_eco7683, w_eco7684, w_eco7685, w_eco7686, w_eco7687, w_eco7688, w_eco7689, w_eco7690, w_eco7691, w_eco7692, w_eco7693, w_eco7694, w_eco7695, w_eco7696, w_eco7697, w_eco7698, w_eco7699, w_eco7700, w_eco7701, w_eco7702, w_eco7703, w_eco7704, w_eco7705, w_eco7706, w_eco7707, w_eco7708, w_eco7709, w_eco7710, w_eco7711, w_eco7712, w_eco7713, w_eco7714, w_eco7715, w_eco7716, w_eco7717, w_eco7718, w_eco7719, w_eco7720, w_eco7721, w_eco7722, w_eco7723, w_eco7724, w_eco7725, w_eco7726, w_eco7727, w_eco7728, w_eco7729, w_eco7730, w_eco7731, w_eco7732, w_eco7733, w_eco7734, w_eco7735, w_eco7736, w_eco7737, w_eco7738, w_eco7739, w_eco7740, w_eco7741, w_eco7742, w_eco7743, w_eco7744, w_eco7745, w_eco7746, w_eco7747, w_eco7748, w_eco7749, w_eco7750, w_eco7751, w_eco7752, w_eco7753, w_eco7754, w_eco7755, w_eco7756, w_eco7757, w_eco7758, w_eco7759, w_eco7760, w_eco7761, w_eco7762, w_eco7763, w_eco7764, w_eco7765, w_eco7766, w_eco7767, w_eco7768, w_eco7769, w_eco7770, w_eco7771, w_eco7772, w_eco7773, w_eco7774, w_eco7775, w_eco7776, w_eco7777, w_eco7778, w_eco7779, w_eco7780, w_eco7781, w_eco7782, w_eco7783, w_eco7784, w_eco7785, w_eco7786, w_eco7787, w_eco7788, w_eco7789, w_eco7790, w_eco7791, w_eco7792, w_eco7793, w_eco7794, w_eco7795, w_eco7796, w_eco7797, w_eco7798);
	xor _ECO_out5(cnt[3], sub_wire5, w_eco7799);
	assign w_eco7800 = rst;
	and _ECO_7801(w_eco7801, Tsync[2], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_7802(w_eco7802, Tsync[2], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7803(w_eco7803, Tsync[2], !prev_cnt[5], ena, !prev_state[0]);
	and _ECO_7804(w_eco7804, !Tsync[5], Tsync[2], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_7805(w_eco7805, Tsync[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1]);
	and _ECO_7806(w_eco7806, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_state[1]);
	and _ECO_7807(w_eco7807, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], !ena);
	and _ECO_7808(w_eco7808, Tgate[2], prev_cnt[1], prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7809(w_eco7809, Tgate[2], prev_cnt[1], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7810(w_eco7810, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_state[3], !prev_state[2]);
	and _ECO_7811(w_eco7811, Tgate[2], prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1]);
	and _ECO_7812(w_eco7812, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_7813(w_eco7813, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_state[4], !prev_state[2]);
	and _ECO_7814(w_eco7814, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], !ena);
	and _ECO_7815(w_eco7815, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], !ena);
	and _ECO_7816(w_eco7816, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], !ena);
	and _ECO_7817(w_eco7817, !Tsync[5], Tgate[2], prev_cnt[1], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_7818(w_eco7818, !Tsync[5], prev_cnt[1], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7819(w_eco7819, Tgate[2], prev_cnt[0], prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7820(w_eco7820, Tgate[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7821(w_eco7821, prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7822(w_eco7822, Tgate[2], prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0]);
	and _ECO_7823(w_eco7823, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7824(w_eco7824, !Tsync[5], prev_cnt[1], prev_cnt[2], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_7825(w_eco7825, Tgate[2], prev_cnt[0], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7826(w_eco7826, Tgate[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7827(w_eco7827, prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7828(w_eco7828, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7829(w_eco7829, !Tsync[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7830(w_eco7830, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_7831(w_eco7831, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], prev_state[1]);
	and _ECO_7832(w_eco7832, Tgate[2], prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1]);
	and _ECO_7833(w_eco7833, Tgate[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1]);
	and _ECO_7834(w_eco7834, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_7835(w_eco7835, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_7836(w_eco7836, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_7837(w_eco7837, !Tsync[5], prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[0]);
	and _ECO_7838(w_eco7838, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_7839(w_eco7839, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], !ena);
	and _ECO_7840(w_eco7840, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], !ena);
	and _ECO_7841(w_eco7841, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7842(w_eco7842, !Tsync[5], Tgate[2], prev_cnt[0], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_7843(w_eco7843, !Tsync[5], Tgate[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_7844(w_eco7844, !Tsync[5], prev_cnt[0], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7845(w_eco7845, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_7846(w_eco7846, prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7847(w_eco7847, prev_cnt[0], prev_cnt[2], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7848(w_eco7848, Tgate[2], prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0]);
	and _ECO_7849(w_eco7849, Tgate[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0]);
	and _ECO_7850(w_eco7850, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7851(w_eco7851, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7852(w_eco7852, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7853(w_eco7853, !Tsync[5], prev_cnt[0], prev_cnt[2], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_7854(w_eco7854, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_7855(w_eco7855, prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7856(w_eco7856, prev_cnt[0], prev_cnt[2], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7857(w_eco7857, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7858(w_eco7858, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7859(w_eco7859, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_7860(w_eco7860, !Tsync[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7861(w_eco7861, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_7862(w_eco7862, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_7863(w_eco7863, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], prev_state[1]);
	and _ECO_7864(w_eco7864, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], prev_state[1]);
	and _ECO_7865(w_eco7865, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], prev_state[1]);
	and _ECO_7866(w_eco7866, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7867(w_eco7867, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_7868(w_eco7868, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_7869(w_eco7869, !Tsync[5], prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[0]);
	and _ECO_7870(w_eco7870, !Tsync[5], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[0]);
	and _ECO_7871(w_eco7871, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_7872(w_eco7872, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_7873(w_eco7873, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], !ena);
	and _ECO_7874(w_eco7874, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7875(w_eco7875, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7876(w_eco7876, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7877(w_eco7877, prev_cnt[0], prev_cnt[2], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7878(w_eco7878, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7879(w_eco7879, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7880(w_eco7880, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7881(w_eco7881, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7882(w_eco7882, prev_cnt[0], prev_cnt[2], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7883(w_eco7883, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7884(w_eco7884, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_7885(w_eco7885, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_7886(w_eco7886, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_7887(w_eco7887, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_7888(w_eco7888, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7889(w_eco7889, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], prev_state[1]);
	and _ECO_7890(w_eco7890, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], prev_state[1]);
	and _ECO_7891(w_eco7891, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_7892(w_eco7892, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7893(w_eco7893, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7894(w_eco7894, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7895(w_eco7895, !Tgate[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7896(w_eco7896, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], !ena);
	and _ECO_7897(w_eco7897, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], !ena);
	and _ECO_7898(w_eco7898, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], !ena);
	and _ECO_7899(w_eco7899, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7900(w_eco7900, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7901(w_eco7901, Tgdel[2], prev_cnt[1], prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7902(w_eco7902, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7903(w_eco7903, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7904(w_eco7904, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7905(w_eco7905, Tgdel[2], prev_cnt[1], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7906(w_eco7906, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7907(w_eco7907, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_7908(w_eco7908, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_7909(w_eco7909, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_7910(w_eco7910, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_7911(w_eco7911, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_7912(w_eco7912, !Tsync[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7913(w_eco7913, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7914(w_eco7914, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7915(w_eco7915, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7916(w_eco7916, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], prev_state[1]);
	and _ECO_7917(w_eco7917, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_7918(w_eco7918, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_7919(w_eco7919, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_7920(w_eco7920, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7921(w_eco7921, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7922(w_eco7922, !Tgate[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7923(w_eco7923, !Tgate[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_7924(w_eco7924, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], !ena);
	and _ECO_7925(w_eco7925, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], !ena);
	and _ECO_7926(w_eco7926, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], !ena);
	and _ECO_7927(w_eco7927, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7928(w_eco7928, prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7929(w_eco7929, Tgdel[2], prev_cnt[0], prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7930(w_eco7930, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7931(w_eco7931, prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7932(w_eco7932, Tgdel[2], prev_cnt[0], prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7933(w_eco7933, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_7934(w_eco7934, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_7935(w_eco7935, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_7936(w_eco7936, !Tsync[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7937(w_eco7937, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7938(w_eco7938, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7939(w_eco7939, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], prev_state[1]);
	and _ECO_7940(w_eco7940, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], prev_state[1]);
	and _ECO_7941(w_eco7941, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], prev_state[1]);
	and _ECO_7942(w_eco7942, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_7943(w_eco7943, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_7944(w_eco7944, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7945(w_eco7945, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7946(w_eco7946, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], !ena);
	and _ECO_7947(w_eco7947, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], !ena);
	and _ECO_7948(w_eco7948, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], !ena);
	and _ECO_7949(w_eco7949, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7950(w_eco7950, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7951(w_eco7951, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7952(w_eco7952, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7953(w_eco7953, prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7954(w_eco7954, prev_cnt[0], prev_cnt[2], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7955(w_eco7955, Tgdel[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7956(w_eco7956, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7957(w_eco7957, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7958(w_eco7958, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7959(w_eco7959, prev_cnt[14], prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7960(w_eco7960, prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7961(w_eco7961, prev_cnt[0], prev_cnt[2], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7962(w_eco7962, Tgdel[2], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7963(w_eco7963, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_7964(w_eco7964, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_7965(w_eco7965, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_7966(w_eco7966, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_7967(w_eco7967, !Tsync[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7968(w_eco7968, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7969(w_eco7969, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], prev_state[1]);
	and _ECO_7970(w_eco7970, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], prev_state[1]);
	and _ECO_7971(w_eco7971, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], prev_state[1]);
	and _ECO_7972(w_eco7972, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_7973(w_eco7973, prev_cnt[14], prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7974(w_eco7974, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7975(w_eco7975, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7976(w_eco7976, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7977(w_eco7977, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_7978(w_eco7978, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_7979(w_eco7979, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7980(w_eco7980, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7981(w_eco7981, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], !ena);
	and _ECO_7982(w_eco7982, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], !ena);
	and _ECO_7983(w_eco7983, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], !ena);
	and _ECO_7984(w_eco7984, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], !ena);
	and _ECO_7985(w_eco7985, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7986(w_eco7986, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7987(w_eco7987, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_7988(w_eco7988, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_7989(w_eco7989, Tgate[2], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7990(w_eco7990, prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7991(w_eco7991, prev_cnt[0], prev_cnt[2], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7992(w_eco7992, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7993(w_eco7993, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7994(w_eco7994, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7995(w_eco7995, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_7996(w_eco7996, Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_7997(w_eco7997, prev_cnt[14], prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7998(w_eco7998, Tgate[2], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_7999(w_eco7999, prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8000(w_eco8000, prev_cnt[0], prev_cnt[2], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8001(w_eco8001, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8002(w_eco8002, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_8003(w_eco8003, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_8004(w_eco8004, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_8005(w_eco8005, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_8006(w_eco8006, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_8007(w_eco8007, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_8008(w_eco8008, !Tsync[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8009(w_eco8009, prev_cnt[14], prev_cnt[1], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8010(w_eco8010, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8011(w_eco8011, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8012(w_eco8012, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8013(w_eco8013, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8014(w_eco8014, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], prev_state[1]);
	and _ECO_8015(w_eco8015, Tgate[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_8016(w_eco8016, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], prev_state[1]);
	and _ECO_8017(w_eco8017, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], prev_state[1]);
	and _ECO_8018(w_eco8018, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_8019(w_eco8019, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_8020(w_eco8020, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_8021(w_eco8021, Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8022(w_eco8022, prev_cnt[14], prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8023(w_eco8023, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8024(w_eco8024, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8025(w_eco8025, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8026(w_eco8026, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8027(w_eco8027, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_8028(w_eco8028, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_8029(w_eco8029, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8030(w_eco8030, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], !ena);
	and _ECO_8031(w_eco8031, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], !ena);
	and _ECO_8032(w_eco8032, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], !ena);
	and _ECO_8033(w_eco8033, !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], !ena);
	and _ECO_8034(w_eco8034, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], !ena);
	and _ECO_8035(w_eco8035, Tsync[5], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8036(w_eco8036, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8037(w_eco8037, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8038(w_eco8038, !Tsync[5], Tgate[2], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_8039(w_eco8039, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8040(w_eco8040, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8041(w_eco8041, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8042(w_eco8042, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8043(w_eco8043, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8044(w_eco8044, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8045(w_eco8045, prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8046(w_eco8046, prev_cnt[0], prev_cnt[2], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8047(w_eco8047, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8048(w_eco8048, Tgate[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_8049(w_eco8049, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8050(w_eco8050, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8051(w_eco8051, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8052(w_eco8052, !Tsync[5], Tgate[2], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_8053(w_eco8053, prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8054(w_eco8054, Tgdel[2], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_8055(w_eco8055, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8056(w_eco8056, prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8057(w_eco8057, prev_cnt[0], prev_cnt[2], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8058(w_eco8058, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8059(w_eco8059, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_8060(w_eco8060, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_8061(w_eco8061, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_8062(w_eco8062, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_8063(w_eco8063, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_8064(w_eco8064, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_8065(w_eco8065, !Tsync[2], !prev_cnt[14], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8066(w_eco8066, !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8067(w_eco8067, Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8068(w_eco8068, prev_cnt[14], prev_cnt[0], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8069(w_eco8069, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8070(w_eco8070, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8071(w_eco8071, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8072(w_eco8072, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8073(w_eco8073, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], prev_state[1]);
	and _ECO_8074(w_eco8074, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], prev_state[1]);
	and _ECO_8075(w_eco8075, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], prev_state[1]);
	and _ECO_8076(w_eco8076, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_state[1]);
	and _ECO_8077(w_eco8077, Tgdel[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_8078(w_eco8078, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_8079(w_eco8079, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_8080(w_eco8080, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_8081(w_eco8081, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8082(w_eco8082, prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8083(w_eco8083, Tgdel[2], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8084(w_eco8084, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8085(w_eco8085, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8086(w_eco8086, Tgate[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_8087(w_eco8087, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8088(w_eco8088, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8089(w_eco8089, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8090(w_eco8090, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8091(w_eco8091, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8092(w_eco8092, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8093(w_eco8093, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8094(w_eco8094, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8095(w_eco8095, !Tsync[5], Tgate[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_8096(w_eco8096, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8097(w_eco8097, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_8098(w_eco8098, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_8099(w_eco8099, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8100(w_eco8100, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], !ena);
	and _ECO_8101(w_eco8101, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], !ena);
	and _ECO_8102(w_eco8102, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8103(w_eco8103, Tsync[5], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8104(w_eco8104, Tsync[5], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8105(w_eco8105, Tsync[5], !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8106(w_eco8106, !Tsync[5], Tgdel[2], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_8107(w_eco8107, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8108(w_eco8108, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8109(w_eco8109, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8110(w_eco8110, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8111(w_eco8111, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8112(w_eco8112, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8113(w_eco8113, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8114(w_eco8114, Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8115(w_eco8115, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8116(w_eco8116, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8117(w_eco8117, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8118(w_eco8118, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8119(w_eco8119, !Tsync[5], Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_8120(w_eco8120, Tgdel[2], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_8121(w_eco8121, prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8122(w_eco8122, Tgdel[2], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_8123(w_eco8123, !prev_cnt[14], prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8124(w_eco8124, prev_cnt[0], prev_cnt[2], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8125(w_eco8125, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8126(w_eco8126, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8127(w_eco8127, Tgdel[2], prev_cnt[14], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8128(w_eco8128, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_8129(w_eco8129, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_8130(w_eco8130, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_8131(w_eco8131, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_state[3], prev_state[0]);
	and _ECO_8132(w_eco8132, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_8133(w_eco8133, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_8134(w_eco8134, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_8135(w_eco8135, !Tsync[2], !prev_cnt[14], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8136(w_eco8136, prev_cnt[1], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8137(w_eco8137, !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8138(w_eco8138, Tgdel[2], prev_cnt[14], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8139(w_eco8139, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8140(w_eco8140, Tgdel[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_8141(w_eco8141, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8142(w_eco8142, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8143(w_eco8143, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8144(w_eco8144, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8145(w_eco8145, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8146(w_eco8146, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8147(w_eco8147, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8148(w_eco8148, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8149(w_eco8149, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8150(w_eco8150, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], prev_state[1]);
	and _ECO_8151(w_eco8151, Tgate[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_8152(w_eco8152, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], prev_state[1]);
	and _ECO_8153(w_eco8153, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], prev_state[1]);
	and _ECO_8154(w_eco8154, !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_state[1]);
	and _ECO_8155(w_eco8155, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_state[1]);
	and _ECO_8156(w_eco8156, !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_8157(w_eco8157, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_8158(w_eco8158, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_8159(w_eco8159, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8160(w_eco8160, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8161(w_eco8161, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8162(w_eco8162, Tgdel[2], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8163(w_eco8163, prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8164(w_eco8164, Tgdel[2], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8165(w_eco8165, !prev_cnt[14], prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8166(w_eco8166, prev_cnt[0], prev_cnt[2], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8167(w_eco8167, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8168(w_eco8168, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8169(w_eco8169, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8170(w_eco8170, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8171(w_eco8171, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8172(w_eco8172, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8173(w_eco8173, Tgdel[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_8174(w_eco8174, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8175(w_eco8175, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8176(w_eco8176, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8177(w_eco8177, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8178(w_eco8178, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8179(w_eco8179, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8180(w_eco8180, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8181(w_eco8181, !Tsync[5], Tgdel[2], prev_cnt[14], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_8182(w_eco8182, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8183(w_eco8183, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_8184(w_eco8184, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_8185(w_eco8185, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8186(w_eco8186, Tsync[5], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8187(w_eco8187, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8188(w_eco8188, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8189(w_eco8189, Tsync[5], !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8190(w_eco8190, Tsync[5], !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8191(w_eco8191, !Tsync[5], Tgate[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_8192(w_eco8192, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8193(w_eco8193, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8194(w_eco8194, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8195(w_eco8195, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8196(w_eco8196, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8197(w_eco8197, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8198(w_eco8198, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8199(w_eco8199, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8200(w_eco8200, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8201(w_eco8201, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8202(w_eco8202, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8203(w_eco8203, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8204(w_eco8204, Tgate[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_8205(w_eco8205, Tgdel[2], prev_cnt[14], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8206(w_eco8206, Tgdel[2], prev_cnt[14], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8207(w_eco8207, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8208(w_eco8208, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8209(w_eco8209, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8210(w_eco8210, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8211(w_eco8211, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8212(w_eco8212, !Tsync[5], Tgate[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_8213(w_eco8213, Tgdel[2], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_8214(w_eco8214, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8215(w_eco8215, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8216(w_eco8216, Tgdel[2], prev_cnt[14], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8217(w_eco8217, Tgdel[2], prev_cnt[14], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8218(w_eco8218, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_8219(w_eco8219, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_8220(w_eco8220, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_8221(w_eco8221, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_state[3], prev_state[0]);
	and _ECO_8222(w_eco8222, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_state[3], prev_state[0]);
	and _ECO_8223(w_eco8223, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_8224(w_eco8224, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_8225(w_eco8225, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_8226(w_eco8226, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_state[4], !prev_state[2]);
	and _ECO_8227(w_eco8227, Tgdel[2], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8228(w_eco8228, prev_cnt[0], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8229(w_eco8229, !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8230(w_eco8230, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8231(w_eco8231, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8232(w_eco8232, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8233(w_eco8233, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8234(w_eco8234, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8235(w_eco8235, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8236(w_eco8236, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8237(w_eco8237, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8238(w_eco8238, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8239(w_eco8239, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8240(w_eco8240, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8241(w_eco8241, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8242(w_eco8242, Tgate[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8243(w_eco8243, !prev_cnt[14], prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8244(w_eco8244, !prev_cnt[14], prev_cnt[0], prev_cnt[2], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8245(w_eco8245, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8246(w_eco8246, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], prev_state[1]);
	and _ECO_8247(w_eco8247, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], prev_state[1]);
	and _ECO_8248(w_eco8248, Tgdel[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_8249(w_eco8249, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_8250(w_eco8250, !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_8251(w_eco8251, !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_8252(w_eco8252, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_state[3], prev_state[0]);
	and _ECO_8253(w_eco8253, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8254(w_eco8254, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8255(w_eco8255, Tgdel[2], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8256(w_eco8256, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8257(w_eco8257, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8258(w_eco8258, !Tgate[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_8259(w_eco8259, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8260(w_eco8260, Tgate[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_8261(w_eco8261, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8262(w_eco8262, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8263(w_eco8263, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8264(w_eco8264, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8265(w_eco8265, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8266(w_eco8266, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8267(w_eco8267, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8268(w_eco8268, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8269(w_eco8269, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8270(w_eco8270, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8271(w_eco8271, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8272(w_eco8272, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8273(w_eco8273, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8274(w_eco8274, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8275(w_eco8275, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8276(w_eco8276, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8277(w_eco8277, Tgdel[2], prev_cnt[14], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8278(w_eco8278, !Tsync[5], Tgate[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_8279(w_eco8279, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8280(w_eco8280, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_8281(w_eco8281, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_8282(w_eco8282, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8283(w_eco8283, Tsync[5], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8284(w_eco8284, Tsync[5], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8285(w_eco8285, !Tsync[5], Tgdel[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_8286(w_eco8286, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8287(w_eco8287, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8288(w_eco8288, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8289(w_eco8289, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8290(w_eco8290, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8291(w_eco8291, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8292(w_eco8292, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8293(w_eco8293, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8294(w_eco8294, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8295(w_eco8295, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8296(w_eco8296, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8297(w_eco8297, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8298(w_eco8298, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8299(w_eco8299, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8300(w_eco8300, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8301(w_eco8301, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8302(w_eco8302, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8303(w_eco8303, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8304(w_eco8304, Tgdel[2], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8305(w_eco8305, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8306(w_eco8306, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_8307(w_eco8307, !Tsync[5], Tgdel[2], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_8308(w_eco8308, !Tsync[5], Tgdel[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_8309(w_eco8309, Tgdel[2], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_8310(w_eco8310, !prev_cnt[14], prev_cnt[0], prev_cnt[2], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8311(w_eco8311, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8312(w_eco8312, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8313(w_eco8313, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8314(w_eco8314, Tgate[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8315(w_eco8315, !prev_cnt[14], prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8316(w_eco8316, !prev_cnt[14], prev_cnt[0], prev_cnt[2], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8317(w_eco8317, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8318(w_eco8318, Tgdel[2], prev_cnt[1], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8319(w_eco8319, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_8320(w_eco8320, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_8321(w_eco8321, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_8322(w_eco8322, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_8323(w_eco8323, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_8324(w_eco8324, !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], !prev_state[4], !prev_state[2]);
	and _ECO_8325(w_eco8325, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], !prev_state[4], !prev_state[2]);
	and _ECO_8326(w_eco8326, Tgdel[2], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8327(w_eco8327, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[3], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8328(w_eco8328, Tgdel[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_8329(w_eco8329, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8330(w_eco8330, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8331(w_eco8331, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8332(w_eco8332, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8333(w_eco8333, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8334(w_eco8334, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8335(w_eco8335, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8336(w_eco8336, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8337(w_eco8337, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8338(w_eco8338, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8339(w_eco8339, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8340(w_eco8340, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8341(w_eco8341, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8342(w_eco8342, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8343(w_eco8343, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8344(w_eco8344, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8345(w_eco8345, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8346(w_eco8346, !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_8347(w_eco8347, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_8348(w_eco8348, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_8349(w_eco8349, !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], !prev_state[3], prev_state[0]);
	and _ECO_8350(w_eco8350, !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], !prev_state[3], prev_state[0]);
	and _ECO_8351(w_eco8351, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8352(w_eco8352, Tgdel[2], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8353(w_eco8353, !prev_cnt[14], prev_cnt[0], prev_cnt[2], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8354(w_eco8354, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8355(w_eco8355, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8356(w_eco8356, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_8357(w_eco8357, !Tgate[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_8358(w_eco8358, !Tgate[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_8359(w_eco8359, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8360(w_eco8360, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8361(w_eco8361, Tgdel[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_8362(w_eco8362, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8363(w_eco8363, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8364(w_eco8364, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8365(w_eco8365, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8366(w_eco8366, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8367(w_eco8367, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8368(w_eco8368, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8369(w_eco8369, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8370(w_eco8370, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8371(w_eco8371, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8372(w_eco8372, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8373(w_eco8373, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8374(w_eco8374, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8375(w_eco8375, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8376(w_eco8376, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8377(w_eco8377, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8378(w_eco8378, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8379(w_eco8379, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8380(w_eco8380, !Tsync[5], Tgdel[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_8381(w_eco8381, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8382(w_eco8382, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_8383(w_eco8383, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_8384(w_eco8384, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_8385(w_eco8385, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8386(w_eco8386, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8387(w_eco8387, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8388(w_eco8388, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8389(w_eco8389, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8390(w_eco8390, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8391(w_eco8391, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8392(w_eco8392, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8393(w_eco8393, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8394(w_eco8394, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8395(w_eco8395, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8396(w_eco8396, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8397(w_eco8397, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8398(w_eco8398, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8399(w_eco8399, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8400(w_eco8400, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8401(w_eco8401, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8402(w_eco8402, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8403(w_eco8403, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8404(w_eco8404, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8405(w_eco8405, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8406(w_eco8406, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8407(w_eco8407, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8408(w_eco8408, Tgdel[2], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8409(w_eco8409, Tgdel[2], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_8410(w_eco8410, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8411(w_eco8411, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8412(w_eco8412, Tgdel[2], prev_cnt[2], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8413(w_eco8413, Tgdel[2], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_8414(w_eco8414, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_8415(w_eco8415, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_8416(w_eco8416, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8417(w_eco8417, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8418(w_eco8418, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_8419(w_eco8419, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8420(w_eco8420, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8421(w_eco8421, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8422(w_eco8422, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8423(w_eco8423, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8424(w_eco8424, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8425(w_eco8425, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8426(w_eco8426, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8427(w_eco8427, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8428(w_eco8428, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8429(w_eco8429, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8430(w_eco8430, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8431(w_eco8431, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8432(w_eco8432, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8433(w_eco8433, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8434(w_eco8434, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8435(w_eco8435, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8436(w_eco8436, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8437(w_eco8437, !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_8438(w_eco8438, !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_8439(w_eco8439, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8440(w_eco8440, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8441(w_eco8441, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8442(w_eco8442, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8443(w_eco8443, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8444(w_eco8444, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8445(w_eco8445, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8446(w_eco8446, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8447(w_eco8447, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8448(w_eco8448, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8449(w_eco8449, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8450(w_eco8450, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8451(w_eco8451, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8452(w_eco8452, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8453(w_eco8453, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8454(w_eco8454, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8455(w_eco8455, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8456(w_eco8456, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8457(w_eco8457, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8458(w_eco8458, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8459(w_eco8459, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8460(w_eco8460, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8461(w_eco8461, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8462(w_eco8462, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8463(w_eco8463, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8464(w_eco8464, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8465(w_eco8465, Tgdel[2], prev_cnt[0], !prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_8466(w_eco8466, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8467(w_eco8467, prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_8468(w_eco8468, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_8469(w_eco8469, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_8470(w_eco8470, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8471(w_eco8471, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8472(w_eco8472, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8473(w_eco8473, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8474(w_eco8474, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8475(w_eco8475, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8476(w_eco8476, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8477(w_eco8477, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8478(w_eco8478, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8479(w_eco8479, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8480(w_eco8480, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8481(w_eco8481, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8482(w_eco8482, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8483(w_eco8483, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8484(w_eco8484, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8485(w_eco8485, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8486(w_eco8486, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8487(w_eco8487, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8488(w_eco8488, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8489(w_eco8489, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8490(w_eco8490, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8491(w_eco8491, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8492(w_eco8492, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8493(w_eco8493, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8494(w_eco8494, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8495(w_eco8495, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8496(w_eco8496, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8497(w_eco8497, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8498(w_eco8498, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_8499(w_eco8499, !Tsync[5], Tgdel[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_8500(w_eco8500, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_8501(w_eco8501, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_8502(w_eco8502, !prev_cnt[14], prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_8503(w_eco8503, prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_8504(w_eco8504, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_8505(w_eco8505, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8506(w_eco8506, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8507(w_eco8507, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8508(w_eco8508, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8509(w_eco8509, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8510(w_eco8510, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8511(w_eco8511, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8512(w_eco8512, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8513(w_eco8513, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8514(w_eco8514, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8515(w_eco8515, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8516(w_eco8516, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8517(w_eco8517, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8518(w_eco8518, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8519(w_eco8519, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8520(w_eco8520, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8521(w_eco8521, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8522(w_eco8522, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8523(w_eco8523, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8524(w_eco8524, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8525(w_eco8525, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8526(w_eco8526, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8527(w_eco8527, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8528(w_eco8528, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8529(w_eco8529, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8530(w_eco8530, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8531(w_eco8531, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8532(w_eco8532, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8533(w_eco8533, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8534(w_eco8534, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8535(w_eco8535, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8536(w_eco8536, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8537(w_eco8537, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8538(w_eco8538, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8539(w_eco8539, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8540(w_eco8540, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8541(w_eco8541, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8542(w_eco8542, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8543(w_eco8543, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8544(w_eco8544, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8545(w_eco8545, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8546(w_eco8546, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8547(w_eco8547, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8548(w_eco8548, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8549(w_eco8549, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8550(w_eco8550, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8551(w_eco8551, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8552(w_eco8552, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8553(w_eco8553, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8554(w_eco8554, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8555(w_eco8555, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8556(w_eco8556, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8557(w_eco8557, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8558(w_eco8558, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8559(w_eco8559, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8560(w_eco8560, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8561(w_eco8561, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8562(w_eco8562, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8563(w_eco8563, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8564(w_eco8564, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_8565(w_eco8565, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8566(w_eco8566, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8567(w_eco8567, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8568(w_eco8568, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8569(w_eco8569, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8570(w_eco8570, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8571(w_eco8571, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8572(w_eco8572, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8573(w_eco8573, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8574(w_eco8574, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8575(w_eco8575, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8576(w_eco8576, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8577(w_eco8577, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8578(w_eco8578, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8579(w_eco8579, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8580(w_eco8580, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8581(w_eco8581, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8582(w_eco8582, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8583(w_eco8583, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8584(w_eco8584, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8585(w_eco8585, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8586(w_eco8586, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8587(w_eco8587, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8588(w_eco8588, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8589(w_eco8589, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8590(w_eco8590, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8591(w_eco8591, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8592(w_eco8592, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8593(w_eco8593, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8594(w_eco8594, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8595(w_eco8595, !prev_cnt[14], prev_cnt[1], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_8596(w_eco8596, !prev_cnt[14], prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_8597(w_eco8597, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_8598(w_eco8598, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8599(w_eco8599, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8600(w_eco8600, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8601(w_eco8601, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8602(w_eco8602, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8603(w_eco8603, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8604(w_eco8604, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8605(w_eco8605, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8606(w_eco8606, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8607(w_eco8607, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8608(w_eco8608, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8609(w_eco8609, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8610(w_eco8610, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8611(w_eco8611, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8612(w_eco8612, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8613(w_eco8613, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8614(w_eco8614, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8615(w_eco8615, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8616(w_eco8616, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8617(w_eco8617, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8618(w_eco8618, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8619(w_eco8619, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8620(w_eco8620, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8621(w_eco8621, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8622(w_eco8622, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8623(w_eco8623, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8624(w_eco8624, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8625(w_eco8625, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8626(w_eco8626, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8627(w_eco8627, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8628(w_eco8628, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8629(w_eco8629, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8630(w_eco8630, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8631(w_eco8631, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8632(w_eco8632, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8633(w_eco8633, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8634(w_eco8634, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8635(w_eco8635, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8636(w_eco8636, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8637(w_eco8637, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8638(w_eco8638, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8639(w_eco8639, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8640(w_eco8640, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8641(w_eco8641, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8642(w_eco8642, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8643(w_eco8643, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8644(w_eco8644, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8645(w_eco8645, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8646(w_eco8646, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8647(w_eco8647, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8648(w_eco8648, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8649(w_eco8649, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8650(w_eco8650, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8651(w_eco8651, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8652(w_eco8652, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8653(w_eco8653, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8654(w_eco8654, !Tsync[5], Tsync[2], !prev_cnt[5], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8655(w_eco8655, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8656(w_eco8656, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8657(w_eco8657, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8658(w_eco8658, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8659(w_eco8659, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8660(w_eco8660, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8661(w_eco8661, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8662(w_eco8662, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8663(w_eco8663, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8664(w_eco8664, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8665(w_eco8665, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8666(w_eco8666, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8667(w_eco8667, Tsync[5], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8668(w_eco8668, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8669(w_eco8669, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8670(w_eco8670, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8671(w_eco8671, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8672(w_eco8672, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8673(w_eco8673, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8674(w_eco8674, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8675(w_eco8675, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8676(w_eco8676, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8677(w_eco8677, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8678(w_eco8678, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8679(w_eco8679, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8680(w_eco8680, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8681(w_eco8681, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8682(w_eco8682, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8683(w_eco8683, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8684(w_eco8684, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8685(w_eco8685, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8686(w_eco8686, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8687(w_eco8687, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8688(w_eco8688, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8689(w_eco8689, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8690(w_eco8690, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8691(w_eco8691, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8692(w_eco8692, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8693(w_eco8693, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8694(w_eco8694, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8695(w_eco8695, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8696(w_eco8696, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8697(w_eco8697, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8698(w_eco8698, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8699(w_eco8699, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8700(w_eco8700, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8701(w_eco8701, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8702(w_eco8702, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8703(w_eco8703, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8704(w_eco8704, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8705(w_eco8705, !prev_cnt[14], prev_cnt[0], prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_8706(w_eco8706, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_8707(w_eco8707, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8708(w_eco8708, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8709(w_eco8709, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8710(w_eco8710, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8711(w_eco8711, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8712(w_eco8712, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8713(w_eco8713, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8714(w_eco8714, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8715(w_eco8715, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8716(w_eco8716, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8717(w_eco8717, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8718(w_eco8718, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8719(w_eco8719, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8720(w_eco8720, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8721(w_eco8721, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8722(w_eco8722, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8723(w_eco8723, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8724(w_eco8724, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8725(w_eco8725, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8726(w_eco8726, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8727(w_eco8727, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8728(w_eco8728, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8729(w_eco8729, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8730(w_eco8730, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8731(w_eco8731, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8732(w_eco8732, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8733(w_eco8733, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8734(w_eco8734, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8735(w_eco8735, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8736(w_eco8736, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8737(w_eco8737, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8738(w_eco8738, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8739(w_eco8739, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8740(w_eco8740, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8741(w_eco8741, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8742(w_eco8742, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8743(w_eco8743, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8744(w_eco8744, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8745(w_eco8745, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8746(w_eco8746, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8747(w_eco8747, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8748(w_eco8748, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8749(w_eco8749, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8750(w_eco8750, !Tsync[5], Tsync[2], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8751(w_eco8751, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8752(w_eco8752, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8753(w_eco8753, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8754(w_eco8754, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8755(w_eco8755, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8756(w_eco8756, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8757(w_eco8757, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8758(w_eco8758, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8759(w_eco8759, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8760(w_eco8760, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8761(w_eco8761, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8762(w_eco8762, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8763(w_eco8763, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8764(w_eco8764, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8765(w_eco8765, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8766(w_eco8766, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8767(w_eco8767, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8768(w_eco8768, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8769(w_eco8769, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8770(w_eco8770, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8771(w_eco8771, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8772(w_eco8772, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8773(w_eco8773, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8774(w_eco8774, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8775(w_eco8775, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8776(w_eco8776, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8777(w_eco8777, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8778(w_eco8778, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8779(w_eco8779, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8780(w_eco8780, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8781(w_eco8781, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8782(w_eco8782, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8783(w_eco8783, !Tsync[5], Tsync[2], !prev_cnt[5], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8784(w_eco8784, !Tsync[5], Tsync[2], !prev_cnt[5], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8785(w_eco8785, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8786(w_eco8786, Tsync[5], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8787(w_eco8787, Tsync[5], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8788(w_eco8788, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[1], !prev_cnt[2], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8789(w_eco8789, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8790(w_eco8790, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8791(w_eco8791, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8792(w_eco8792, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8793(w_eco8793, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8794(w_eco8794, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8795(w_eco8795, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8796(w_eco8796, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8797(w_eco8797, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8798(w_eco8798, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8799(w_eco8799, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8800(w_eco8800, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8801(w_eco8801, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8802(w_eco8802, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8803(w_eco8803, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8804(w_eco8804, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8805(w_eco8805, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8806(w_eco8806, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8807(w_eco8807, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8808(w_eco8808, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8809(w_eco8809, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8810(w_eco8810, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8811(w_eco8811, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8812(w_eco8812, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8813(w_eco8813, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8814(w_eco8814, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8815(w_eco8815, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8816(w_eco8816, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8817(w_eco8817, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8818(w_eco8818, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8819(w_eco8819, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8820(w_eco8820, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8821(w_eco8821, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8822(w_eco8822, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8823(w_eco8823, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8824(w_eco8824, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8825(w_eco8825, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8826(w_eco8826, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8827(w_eco8827, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8828(w_eco8828, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8829(w_eco8829, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8830(w_eco8830, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8831(w_eco8831, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8832(w_eco8832, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8833(w_eco8833, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_8834(w_eco8834, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8835(w_eco8835, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8836(w_eco8836, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8837(w_eco8837, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8838(w_eco8838, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8839(w_eco8839, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8840(w_eco8840, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8841(w_eco8841, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8842(w_eco8842, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8843(w_eco8843, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8844(w_eco8844, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8845(w_eco8845, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8846(w_eco8846, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8847(w_eco8847, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8848(w_eco8848, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8849(w_eco8849, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8850(w_eco8850, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8851(w_eco8851, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8852(w_eco8852, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8853(w_eco8853, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8854(w_eco8854, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8855(w_eco8855, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8856(w_eco8856, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8857(w_eco8857, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8858(w_eco8858, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8859(w_eco8859, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8860(w_eco8860, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8861(w_eco8861, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8862(w_eco8862, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8863(w_eco8863, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8864(w_eco8864, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8865(w_eco8865, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8866(w_eco8866, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8867(w_eco8867, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8868(w_eco8868, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8869(w_eco8869, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8870(w_eco8870, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8871(w_eco8871, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8872(w_eco8872, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8873(w_eco8873, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8874(w_eco8874, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8875(w_eco8875, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8876(w_eco8876, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8877(w_eco8877, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8878(w_eco8878, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8879(w_eco8879, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8880(w_eco8880, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8881(w_eco8881, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8882(w_eco8882, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8883(w_eco8883, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8884(w_eco8884, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8885(w_eco8885, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8886(w_eco8886, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8887(w_eco8887, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8888(w_eco8888, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8889(w_eco8889, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8890(w_eco8890, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8891(w_eco8891, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8892(w_eco8892, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8893(w_eco8893, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8894(w_eco8894, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8895(w_eco8895, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8896(w_eco8896, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8897(w_eco8897, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8898(w_eco8898, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8899(w_eco8899, !Tsync[5], Tsync[2], !prev_cnt[5], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8900(w_eco8900, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8901(w_eco8901, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8902(w_eco8902, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8903(w_eco8903, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8904(w_eco8904, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8905(w_eco8905, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8906(w_eco8906, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8907(w_eco8907, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8908(w_eco8908, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8909(w_eco8909, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8910(w_eco8910, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8911(w_eco8911, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8912(w_eco8912, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8913(w_eco8913, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8914(w_eco8914, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8915(w_eco8915, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8916(w_eco8916, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8917(w_eco8917, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8918(w_eco8918, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8919(w_eco8919, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8920(w_eco8920, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8921(w_eco8921, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8922(w_eco8922, Tsync[5], !Tgate[2], !Tgdel[2], !Tsync[2], prev_cnt[0], !prev_cnt[2], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_8923(w_eco8923, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8924(w_eco8924, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8925(w_eco8925, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8926(w_eco8926, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8927(w_eco8927, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8928(w_eco8928, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8929(w_eco8929, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8930(w_eco8930, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8931(w_eco8931, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8932(w_eco8932, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8933(w_eco8933, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8934(w_eco8934, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8935(w_eco8935, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8936(w_eco8936, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8937(w_eco8937, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8938(w_eco8938, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8939(w_eco8939, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8940(w_eco8940, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8941(w_eco8941, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8942(w_eco8942, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8943(w_eco8943, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8944(w_eco8944, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8945(w_eco8945, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8946(w_eco8946, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8947(w_eco8947, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8948(w_eco8948, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8949(w_eco8949, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8950(w_eco8950, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8951(w_eco8951, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8952(w_eco8952, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8953(w_eco8953, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8954(w_eco8954, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8955(w_eco8955, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8956(w_eco8956, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_8957(w_eco8957, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8958(w_eco8958, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8959(w_eco8959, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8960(w_eco8960, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8961(w_eco8961, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8962(w_eco8962, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8963(w_eco8963, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8964(w_eco8964, Tsync[2], !prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8965(w_eco8965, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8966(w_eco8966, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8967(w_eco8967, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8968(w_eco8968, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8969(w_eco8969, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8970(w_eco8970, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_8971(w_eco8971, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8972(w_eco8972, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_8973(w_eco8973, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8974(w_eco8974, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8975(w_eco8975, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8976(w_eco8976, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8977(w_eco8977, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8978(w_eco8978, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8979(w_eco8979, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8980(w_eco8980, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8981(w_eco8981, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8982(w_eco8982, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8983(w_eco8983, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8984(w_eco8984, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8985(w_eco8985, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8986(w_eco8986, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8987(w_eco8987, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8988(w_eco8988, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8989(w_eco8989, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_8990(w_eco8990, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8991(w_eco8991, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8992(w_eco8992, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8993(w_eco8993, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8994(w_eco8994, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8995(w_eco8995, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_8996(w_eco8996, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8997(w_eco8997, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8998(w_eco8998, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_8999(w_eco8999, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9000(w_eco9000, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9001(w_eco9001, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9002(w_eco9002, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9003(w_eco9003, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9004(w_eco9004, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9005(w_eco9005, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9006(w_eco9006, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9007(w_eco9007, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9008(w_eco9008, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9009(w_eco9009, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9010(w_eco9010, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9011(w_eco9011, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9012(w_eco9012, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9013(w_eco9013, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9014(w_eco9014, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9015(w_eco9015, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9016(w_eco9016, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9017(w_eco9017, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9018(w_eco9018, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9019(w_eco9019, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9020(w_eco9020, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9021(w_eco9021, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9022(w_eco9022, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9023(w_eco9023, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9024(w_eco9024, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9025(w_eco9025, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9026(w_eco9026, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9027(w_eco9027, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9028(w_eco9028, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9029(w_eco9029, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9030(w_eco9030, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9031(w_eco9031, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9032(w_eco9032, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9033(w_eco9033, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9034(w_eco9034, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9035(w_eco9035, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9036(w_eco9036, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9037(w_eco9037, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9038(w_eco9038, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9039(w_eco9039, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9040(w_eco9040, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9041(w_eco9041, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9042(w_eco9042, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9043(w_eco9043, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9044(w_eco9044, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9045(w_eco9045, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9046(w_eco9046, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9047(w_eco9047, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9048(w_eco9048, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9049(w_eco9049, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9050(w_eco9050, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9051(w_eco9051, !Tsync[5], Tsync[2], !prev_cnt[5], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9052(w_eco9052, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_9053(w_eco9053, Tsync[5], !Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9054(w_eco9054, Tsync[5], !Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9055(w_eco9055, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9056(w_eco9056, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9057(w_eco9057, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9058(w_eco9058, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9059(w_eco9059, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9060(w_eco9060, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9061(w_eco9061, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9062(w_eco9062, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9063(w_eco9063, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9064(w_eco9064, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9065(w_eco9065, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9066(w_eco9066, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9067(w_eco9067, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9068(w_eco9068, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9069(w_eco9069, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9070(w_eco9070, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9071(w_eco9071, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9072(w_eco9072, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9073(w_eco9073, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9074(w_eco9074, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9075(w_eco9075, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9076(w_eco9076, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9077(w_eco9077, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9078(w_eco9078, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9079(w_eco9079, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9080(w_eco9080, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9081(w_eco9081, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9082(w_eco9082, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9083(w_eco9083, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9084(w_eco9084, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9085(w_eco9085, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9086(w_eco9086, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9087(w_eco9087, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9088(w_eco9088, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9089(w_eco9089, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9090(w_eco9090, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9091(w_eco9091, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9092(w_eco9092, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9093(w_eco9093, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9094(w_eco9094, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9095(w_eco9095, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9096(w_eco9096, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9097(w_eco9097, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9098(w_eco9098, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9099(w_eco9099, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9100(w_eco9100, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9101(w_eco9101, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9102(w_eco9102, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9103(w_eco9103, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9104(w_eco9104, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9105(w_eco9105, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9106(w_eco9106, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9107(w_eco9107, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9108(w_eco9108, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9109(w_eco9109, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9110(w_eco9110, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9111(w_eco9111, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9112(w_eco9112, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9113(w_eco9113, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9114(w_eco9114, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9115(w_eco9115, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9116(w_eco9116, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9117(w_eco9117, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9118(w_eco9118, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9119(w_eco9119, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9120(w_eco9120, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9121(w_eco9121, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9122(w_eco9122, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9123(w_eco9123, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9124(w_eco9124, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9125(w_eco9125, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9126(w_eco9126, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9127(w_eco9127, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9128(w_eco9128, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9129(w_eco9129, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9130(w_eco9130, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9131(w_eco9131, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9132(w_eco9132, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9133(w_eco9133, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9134(w_eco9134, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9135(w_eco9135, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9136(w_eco9136, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9137(w_eco9137, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9138(w_eco9138, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9139(w_eco9139, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9140(w_eco9140, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9141(w_eco9141, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9142(w_eco9142, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9143(w_eco9143, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9144(w_eco9144, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9145(w_eco9145, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9146(w_eco9146, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9147(w_eco9147, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9148(w_eco9148, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9149(w_eco9149, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9150(w_eco9150, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9151(w_eco9151, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9152(w_eco9152, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9153(w_eco9153, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9154(w_eco9154, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9155(w_eco9155, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9156(w_eco9156, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9157(w_eco9157, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9158(w_eco9158, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9159(w_eco9159, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9160(w_eco9160, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9161(w_eco9161, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9162(w_eco9162, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9163(w_eco9163, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9164(w_eco9164, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9165(w_eco9165, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9166(w_eco9166, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9167(w_eco9167, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9168(w_eco9168, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9169(w_eco9169, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9170(w_eco9170, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9171(w_eco9171, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9172(w_eco9172, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9173(w_eco9173, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9174(w_eco9174, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9175(w_eco9175, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9176(w_eco9176, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9177(w_eco9177, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9178(w_eco9178, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9179(w_eco9179, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9180(w_eco9180, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9181(w_eco9181, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9182(w_eco9182, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9183(w_eco9183, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9184(w_eco9184, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9185(w_eco9185, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9186(w_eco9186, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9187(w_eco9187, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9188(w_eco9188, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9189(w_eco9189, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9190(w_eco9190, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9191(w_eco9191, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9192(w_eco9192, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9193(w_eco9193, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9194(w_eco9194, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9195(w_eco9195, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9196(w_eco9196, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9197(w_eco9197, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9198(w_eco9198, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9199(w_eco9199, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9200(w_eco9200, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9201(w_eco9201, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9202(w_eco9202, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9203(w_eco9203, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9204(w_eco9204, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9205(w_eco9205, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9206(w_eco9206, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9207(w_eco9207, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9208(w_eco9208, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9209(w_eco9209, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9210(w_eco9210, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9211(w_eco9211, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9212(w_eco9212, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9213(w_eco9213, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9214(w_eco9214, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9215(w_eco9215, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9216(w_eco9216, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9217(w_eco9217, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9218(w_eco9218, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9219(w_eco9219, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9220(w_eco9220, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9221(w_eco9221, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9222(w_eco9222, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9223(w_eco9223, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9224(w_eco9224, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9225(w_eco9225, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9226(w_eco9226, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9227(w_eco9227, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9228(w_eco9228, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9229(w_eco9229, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9230(w_eco9230, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9231(w_eco9231, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9232(w_eco9232, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9233(w_eco9233, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9234(w_eco9234, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9235(w_eco9235, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9236(w_eco9236, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9237(w_eco9237, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9238(w_eco9238, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9239(w_eco9239, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9240(w_eco9240, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9241(w_eco9241, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9242(w_eco9242, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9243(w_eco9243, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9244(w_eco9244, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9245(w_eco9245, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9246(w_eco9246, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9247(w_eco9247, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9248(w_eco9248, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9249(w_eco9249, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9250(w_eco9250, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9251(w_eco9251, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9252(w_eco9252, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9253(w_eco9253, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9254(w_eco9254, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9255(w_eco9255, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9256(w_eco9256, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9257(w_eco9257, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9258(w_eco9258, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9259(w_eco9259, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9260(w_eco9260, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9261(w_eco9261, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9262(w_eco9262, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9263(w_eco9263, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9264(w_eco9264, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9265(w_eco9265, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9266(w_eco9266, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9267(w_eco9267, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9268(w_eco9268, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9269(w_eco9269, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9270(w_eco9270, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9271(w_eco9271, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9272(w_eco9272, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9273(w_eco9273, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9274(w_eco9274, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9275(w_eco9275, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9276(w_eco9276, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9277(w_eco9277, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9278(w_eco9278, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9279(w_eco9279, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9280(w_eco9280, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9281(w_eco9281, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9282(w_eco9282, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9283(w_eco9283, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9284(w_eco9284, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9285(w_eco9285, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9286(w_eco9286, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9287(w_eco9287, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9288(w_eco9288, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9289(w_eco9289, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9290(w_eco9290, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9291(w_eco9291, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9292(w_eco9292, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9293(w_eco9293, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9294(w_eco9294, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9295(w_eco9295, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9296(w_eco9296, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9297(w_eco9297, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9298(w_eco9298, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9299(w_eco9299, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9300(w_eco9300, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9301(w_eco9301, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9302(w_eco9302, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9303(w_eco9303, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9304(w_eco9304, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9305(w_eco9305, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9306(w_eco9306, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9307(w_eco9307, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9308(w_eco9308, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9309(w_eco9309, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9310(w_eco9310, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9311(w_eco9311, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9312(w_eco9312, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9313(w_eco9313, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9314(w_eco9314, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9315(w_eco9315, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9316(w_eco9316, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9317(w_eco9317, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9318(w_eco9318, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9319(w_eco9319, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9320(w_eco9320, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9321(w_eco9321, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9322(w_eco9322, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9323(w_eco9323, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9324(w_eco9324, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9325(w_eco9325, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9326(w_eco9326, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9327(w_eco9327, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9328(w_eco9328, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9329(w_eco9329, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9330(w_eco9330, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9331(w_eco9331, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9332(w_eco9332, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9333(w_eco9333, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9334(w_eco9334, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9335(w_eco9335, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9336(w_eco9336, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9337(w_eco9337, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9338(w_eco9338, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9339(w_eco9339, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9340(w_eco9340, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9341(w_eco9341, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9342(w_eco9342, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9343(w_eco9343, prev_cnt[1], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9344(w_eco9344, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9345(w_eco9345, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9346(w_eco9346, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9347(w_eco9347, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9348(w_eco9348, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9349(w_eco9349, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9350(w_eco9350, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9351(w_eco9351, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9352(w_eco9352, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9353(w_eco9353, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9354(w_eco9354, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9355(w_eco9355, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9356(w_eco9356, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9357(w_eco9357, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9358(w_eco9358, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9359(w_eco9359, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9360(w_eco9360, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9361(w_eco9361, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9362(w_eco9362, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9363(w_eco9363, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9364(w_eco9364, Tsync[5], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9365(w_eco9365, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9366(w_eco9366, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9367(w_eco9367, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9368(w_eco9368, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9369(w_eco9369, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9370(w_eco9370, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9371(w_eco9371, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9372(w_eco9372, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9373(w_eco9373, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9374(w_eco9374, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9375(w_eco9375, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9376(w_eco9376, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9377(w_eco9377, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9378(w_eco9378, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9379(w_eco9379, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9380(w_eco9380, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9381(w_eco9381, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9382(w_eco9382, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9383(w_eco9383, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9384(w_eco9384, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9385(w_eco9385, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9386(w_eco9386, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9387(w_eco9387, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9388(w_eco9388, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9389(w_eco9389, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9390(w_eco9390, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9391(w_eco9391, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9392(w_eco9392, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9393(w_eco9393, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9394(w_eco9394, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9395(w_eco9395, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9396(w_eco9396, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9397(w_eco9397, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9398(w_eco9398, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9399(w_eco9399, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9400(w_eco9400, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9401(w_eco9401, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9402(w_eco9402, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9403(w_eco9403, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9404(w_eco9404, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9405(w_eco9405, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9406(w_eco9406, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9407(w_eco9407, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9408(w_eco9408, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9409(w_eco9409, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9410(w_eco9410, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9411(w_eco9411, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9412(w_eco9412, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9413(w_eco9413, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9414(w_eco9414, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9415(w_eco9415, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9416(w_eco9416, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9417(w_eco9417, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9418(w_eco9418, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9419(w_eco9419, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9420(w_eco9420, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9421(w_eco9421, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9422(w_eco9422, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9423(w_eco9423, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9424(w_eco9424, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9425(w_eco9425, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9426(w_eco9426, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9427(w_eco9427, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9428(w_eco9428, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9429(w_eco9429, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9430(w_eco9430, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9431(w_eco9431, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9432(w_eco9432, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9433(w_eco9433, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9434(w_eco9434, prev_cnt[0], prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9435(w_eco9435, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9436(w_eco9436, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9437(w_eco9437, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9438(w_eco9438, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9439(w_eco9439, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9440(w_eco9440, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9441(w_eco9441, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9442(w_eco9442, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9443(w_eco9443, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9444(w_eco9444, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9445(w_eco9445, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9446(w_eco9446, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9447(w_eco9447, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9448(w_eco9448, Tsync[5], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9449(w_eco9449, Tsync[5], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9450(w_eco9450, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9451(w_eco9451, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9452(w_eco9452, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9453(w_eco9453, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9454(w_eco9454, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9455(w_eco9455, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9456(w_eco9456, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9457(w_eco9457, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9458(w_eco9458, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9459(w_eco9459, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9460(w_eco9460, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9461(w_eco9461, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9462(w_eco9462, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9463(w_eco9463, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9464(w_eco9464, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9465(w_eco9465, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9466(w_eco9466, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9467(w_eco9467, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9468(w_eco9468, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9469(w_eco9469, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9470(w_eco9470, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9471(w_eco9471, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9472(w_eco9472, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9473(w_eco9473, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9474(w_eco9474, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9475(w_eco9475, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9476(w_eco9476, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9477(w_eco9477, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9478(w_eco9478, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9479(w_eco9479, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9480(w_eco9480, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9481(w_eco9481, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9482(w_eco9482, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9483(w_eco9483, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9484(w_eco9484, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9485(w_eco9485, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9486(w_eco9486, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9487(w_eco9487, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9488(w_eco9488, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9489(w_eco9489, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9490(w_eco9490, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9491(w_eco9491, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9492(w_eco9492, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9493(w_eco9493, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9494(w_eco9494, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9495(w_eco9495, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9496(w_eco9496, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9497(w_eco9497, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9498(w_eco9498, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9499(w_eco9499, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9500(w_eco9500, prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9501(w_eco9501, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9502(w_eco9502, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9503(w_eco9503, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[5], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9504(w_eco9504, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9505(w_eco9505, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9506(w_eco9506, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9507(w_eco9507, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9508(w_eco9508, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9509(w_eco9509, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9510(w_eco9510, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9511(w_eco9511, Tsync[5], !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9512(w_eco9512, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9513(w_eco9513, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9514(w_eco9514, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9515(w_eco9515, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9516(w_eco9516, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9517(w_eco9517, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9518(w_eco9518, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9519(w_eco9519, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9520(w_eco9520, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9521(w_eco9521, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9522(w_eco9522, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9523(w_eco9523, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9524(w_eco9524, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9525(w_eco9525, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9526(w_eco9526, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9527(w_eco9527, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9528(w_eco9528, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9529(w_eco9529, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9530(w_eco9530, Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9531(w_eco9531, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9532(w_eco9532, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9533(w_eco9533, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9534(w_eco9534, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9535(w_eco9535, !Tgate[2], !Tsync[2], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9536(w_eco9536, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9537(w_eco9537, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9538(w_eco9538, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9539(w_eco9539, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9540(w_eco9540, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9541(w_eco9541, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9542(w_eco9542, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9543(w_eco9543, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9544(w_eco9544, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9545(w_eco9545, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9546(w_eco9546, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9547(w_eco9547, prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9548(w_eco9548, !Tgate[2], !Tgdel[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9549(w_eco9549, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9550(w_eco9550, Tsync[5], Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9551(w_eco9551, Tsync[5], Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9552(w_eco9552, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9553(w_eco9553, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9554(w_eco9554, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9555(w_eco9555, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9556(w_eco9556, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9557(w_eco9557, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9558(w_eco9558, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9559(w_eco9559, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9560(w_eco9560, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9561(w_eco9561, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9562(w_eco9562, Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9563(w_eco9563, Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9564(w_eco9564, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[1], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9565(w_eco9565, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9566(w_eco9566, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9567(w_eco9567, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9568(w_eco9568, !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9569(w_eco9569, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9570(w_eco9570, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9571(w_eco9571, !Tgate[2], !Tgdel[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9572(w_eco9572, !Tgate[2], !Tgdel[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9573(w_eco9573, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9574(w_eco9574, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9575(w_eco9575, Tsync[2], !prev_cnt[14], prev_cnt[1], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9576(w_eco9576, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9577(w_eco9577, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9578(w_eco9578, !Tgate[2], !Tgdel[2], Tsync[2], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9579(w_eco9579, !Tgate[2], !Tgdel[2], Tsync[2], prev_cnt[0], !prev_cnt[2], prev_cnt[5], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9580(w_eco9580, !Tgate[2], !Tsync[2], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9581(w_eco9581, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9582(w_eco9582, !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9583(w_eco9583, Tsync[2], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9584(w_eco9584, Tsync[2], !prev_cnt[14], prev_cnt[0], !prev_cnt[2], prev_cnt[5], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_9585(w_eco9585, w_eco7800, w_eco7801, w_eco7802, w_eco7803, w_eco7804, w_eco7805, w_eco7806, w_eco7807, w_eco7808, w_eco7809, w_eco7810, w_eco7811, w_eco7812, w_eco7813, w_eco7814, w_eco7815, w_eco7816, w_eco7817, w_eco7818, w_eco7819, w_eco7820, w_eco7821, w_eco7822, w_eco7823, w_eco7824, w_eco7825, w_eco7826, w_eco7827, w_eco7828, w_eco7829, w_eco7830, w_eco7831, w_eco7832, w_eco7833, w_eco7834, w_eco7835, w_eco7836, w_eco7837, w_eco7838, w_eco7839, w_eco7840, w_eco7841, w_eco7842, w_eco7843, w_eco7844, w_eco7845, w_eco7846, w_eco7847, w_eco7848, w_eco7849, w_eco7850, w_eco7851, w_eco7852, w_eco7853, w_eco7854, w_eco7855, w_eco7856, w_eco7857, w_eco7858, w_eco7859, w_eco7860, w_eco7861, w_eco7862, w_eco7863, w_eco7864, w_eco7865, w_eco7866, w_eco7867, w_eco7868, w_eco7869, w_eco7870, w_eco7871, w_eco7872, w_eco7873, w_eco7874, w_eco7875, w_eco7876, w_eco7877, w_eco7878, w_eco7879, w_eco7880, w_eco7881, w_eco7882, w_eco7883, w_eco7884, w_eco7885, w_eco7886, w_eco7887, w_eco7888, w_eco7889, w_eco7890, w_eco7891, w_eco7892, w_eco7893, w_eco7894, w_eco7895, w_eco7896, w_eco7897, w_eco7898, w_eco7899, w_eco7900, w_eco7901, w_eco7902, w_eco7903, w_eco7904, w_eco7905, w_eco7906, w_eco7907, w_eco7908, w_eco7909, w_eco7910, w_eco7911, w_eco7912, w_eco7913, w_eco7914, w_eco7915, w_eco7916, w_eco7917, w_eco7918, w_eco7919, w_eco7920, w_eco7921, w_eco7922, w_eco7923, w_eco7924, w_eco7925, w_eco7926, w_eco7927, w_eco7928, w_eco7929, w_eco7930, w_eco7931, w_eco7932, w_eco7933, w_eco7934, w_eco7935, w_eco7936, w_eco7937, w_eco7938, w_eco7939, w_eco7940, w_eco7941, w_eco7942, w_eco7943, w_eco7944, w_eco7945, w_eco7946, w_eco7947, w_eco7948, w_eco7949, w_eco7950, w_eco7951, w_eco7952, w_eco7953, w_eco7954, w_eco7955, w_eco7956, w_eco7957, w_eco7958, w_eco7959, w_eco7960, w_eco7961, w_eco7962, w_eco7963, w_eco7964, w_eco7965, w_eco7966, w_eco7967, w_eco7968, w_eco7969, w_eco7970, w_eco7971, w_eco7972, w_eco7973, w_eco7974, w_eco7975, w_eco7976, w_eco7977, w_eco7978, w_eco7979, w_eco7980, w_eco7981, w_eco7982, w_eco7983, w_eco7984, w_eco7985, w_eco7986, w_eco7987, w_eco7988, w_eco7989, w_eco7990, w_eco7991, w_eco7992, w_eco7993, w_eco7994, w_eco7995, w_eco7996, w_eco7997, w_eco7998, w_eco7999, w_eco8000, w_eco8001, w_eco8002, w_eco8003, w_eco8004, w_eco8005, w_eco8006, w_eco8007, w_eco8008, w_eco8009, w_eco8010, w_eco8011, w_eco8012, w_eco8013, w_eco8014, w_eco8015, w_eco8016, w_eco8017, w_eco8018, w_eco8019, w_eco8020, w_eco8021, w_eco8022, w_eco8023, w_eco8024, w_eco8025, w_eco8026, w_eco8027, w_eco8028, w_eco8029, w_eco8030, w_eco8031, w_eco8032, w_eco8033, w_eco8034, w_eco8035, w_eco8036, w_eco8037, w_eco8038, w_eco8039, w_eco8040, w_eco8041, w_eco8042, w_eco8043, w_eco8044, w_eco8045, w_eco8046, w_eco8047, w_eco8048, w_eco8049, w_eco8050, w_eco8051, w_eco8052, w_eco8053, w_eco8054, w_eco8055, w_eco8056, w_eco8057, w_eco8058, w_eco8059, w_eco8060, w_eco8061, w_eco8062, w_eco8063, w_eco8064, w_eco8065, w_eco8066, w_eco8067, w_eco8068, w_eco8069, w_eco8070, w_eco8071, w_eco8072, w_eco8073, w_eco8074, w_eco8075, w_eco8076, w_eco8077, w_eco8078, w_eco8079, w_eco8080, w_eco8081, w_eco8082, w_eco8083, w_eco8084, w_eco8085, w_eco8086, w_eco8087, w_eco8088, w_eco8089, w_eco8090, w_eco8091, w_eco8092, w_eco8093, w_eco8094, w_eco8095, w_eco8096, w_eco8097, w_eco8098, w_eco8099, w_eco8100, w_eco8101, w_eco8102, w_eco8103, w_eco8104, w_eco8105, w_eco8106, w_eco8107, w_eco8108, w_eco8109, w_eco8110, w_eco8111, w_eco8112, w_eco8113, w_eco8114, w_eco8115, w_eco8116, w_eco8117, w_eco8118, w_eco8119, w_eco8120, w_eco8121, w_eco8122, w_eco8123, w_eco8124, w_eco8125, w_eco8126, w_eco8127, w_eco8128, w_eco8129, w_eco8130, w_eco8131, w_eco8132, w_eco8133, w_eco8134, w_eco8135, w_eco8136, w_eco8137, w_eco8138, w_eco8139, w_eco8140, w_eco8141, w_eco8142, w_eco8143, w_eco8144, w_eco8145, w_eco8146, w_eco8147, w_eco8148, w_eco8149, w_eco8150, w_eco8151, w_eco8152, w_eco8153, w_eco8154, w_eco8155, w_eco8156, w_eco8157, w_eco8158, w_eco8159, w_eco8160, w_eco8161, w_eco8162, w_eco8163, w_eco8164, w_eco8165, w_eco8166, w_eco8167, w_eco8168, w_eco8169, w_eco8170, w_eco8171, w_eco8172, w_eco8173, w_eco8174, w_eco8175, w_eco8176, w_eco8177, w_eco8178, w_eco8179, w_eco8180, w_eco8181, w_eco8182, w_eco8183, w_eco8184, w_eco8185, w_eco8186, w_eco8187, w_eco8188, w_eco8189, w_eco8190, w_eco8191, w_eco8192, w_eco8193, w_eco8194, w_eco8195, w_eco8196, w_eco8197, w_eco8198, w_eco8199, w_eco8200, w_eco8201, w_eco8202, w_eco8203, w_eco8204, w_eco8205, w_eco8206, w_eco8207, w_eco8208, w_eco8209, w_eco8210, w_eco8211, w_eco8212, w_eco8213, w_eco8214, w_eco8215, w_eco8216, w_eco8217, w_eco8218, w_eco8219, w_eco8220, w_eco8221, w_eco8222, w_eco8223, w_eco8224, w_eco8225, w_eco8226, w_eco8227, w_eco8228, w_eco8229, w_eco8230, w_eco8231, w_eco8232, w_eco8233, w_eco8234, w_eco8235, w_eco8236, w_eco8237, w_eco8238, w_eco8239, w_eco8240, w_eco8241, w_eco8242, w_eco8243, w_eco8244, w_eco8245, w_eco8246, w_eco8247, w_eco8248, w_eco8249, w_eco8250, w_eco8251, w_eco8252, w_eco8253, w_eco8254, w_eco8255, w_eco8256, w_eco8257, w_eco8258, w_eco8259, w_eco8260, w_eco8261, w_eco8262, w_eco8263, w_eco8264, w_eco8265, w_eco8266, w_eco8267, w_eco8268, w_eco8269, w_eco8270, w_eco8271, w_eco8272, w_eco8273, w_eco8274, w_eco8275, w_eco8276, w_eco8277, w_eco8278, w_eco8279, w_eco8280, w_eco8281, w_eco8282, w_eco8283, w_eco8284, w_eco8285, w_eco8286, w_eco8287, w_eco8288, w_eco8289, w_eco8290, w_eco8291, w_eco8292, w_eco8293, w_eco8294, w_eco8295, w_eco8296, w_eco8297, w_eco8298, w_eco8299, w_eco8300, w_eco8301, w_eco8302, w_eco8303, w_eco8304, w_eco8305, w_eco8306, w_eco8307, w_eco8308, w_eco8309, w_eco8310, w_eco8311, w_eco8312, w_eco8313, w_eco8314, w_eco8315, w_eco8316, w_eco8317, w_eco8318, w_eco8319, w_eco8320, w_eco8321, w_eco8322, w_eco8323, w_eco8324, w_eco8325, w_eco8326, w_eco8327, w_eco8328, w_eco8329, w_eco8330, w_eco8331, w_eco8332, w_eco8333, w_eco8334, w_eco8335, w_eco8336, w_eco8337, w_eco8338, w_eco8339, w_eco8340, w_eco8341, w_eco8342, w_eco8343, w_eco8344, w_eco8345, w_eco8346, w_eco8347, w_eco8348, w_eco8349, w_eco8350, w_eco8351, w_eco8352, w_eco8353, w_eco8354, w_eco8355, w_eco8356, w_eco8357, w_eco8358, w_eco8359, w_eco8360, w_eco8361, w_eco8362, w_eco8363, w_eco8364, w_eco8365, w_eco8366, w_eco8367, w_eco8368, w_eco8369, w_eco8370, w_eco8371, w_eco8372, w_eco8373, w_eco8374, w_eco8375, w_eco8376, w_eco8377, w_eco8378, w_eco8379, w_eco8380, w_eco8381, w_eco8382, w_eco8383, w_eco8384, w_eco8385, w_eco8386, w_eco8387, w_eco8388, w_eco8389, w_eco8390, w_eco8391, w_eco8392, w_eco8393, w_eco8394, w_eco8395, w_eco8396, w_eco8397, w_eco8398, w_eco8399, w_eco8400, w_eco8401, w_eco8402, w_eco8403, w_eco8404, w_eco8405, w_eco8406, w_eco8407, w_eco8408, w_eco8409, w_eco8410, w_eco8411, w_eco8412, w_eco8413, w_eco8414, w_eco8415, w_eco8416, w_eco8417, w_eco8418, w_eco8419, w_eco8420, w_eco8421, w_eco8422, w_eco8423, w_eco8424, w_eco8425, w_eco8426, w_eco8427, w_eco8428, w_eco8429, w_eco8430, w_eco8431, w_eco8432, w_eco8433, w_eco8434, w_eco8435, w_eco8436, w_eco8437, w_eco8438, w_eco8439, w_eco8440, w_eco8441, w_eco8442, w_eco8443, w_eco8444, w_eco8445, w_eco8446, w_eco8447, w_eco8448, w_eco8449, w_eco8450, w_eco8451, w_eco8452, w_eco8453, w_eco8454, w_eco8455, w_eco8456, w_eco8457, w_eco8458, w_eco8459, w_eco8460, w_eco8461, w_eco8462, w_eco8463, w_eco8464, w_eco8465, w_eco8466, w_eco8467, w_eco8468, w_eco8469, w_eco8470, w_eco8471, w_eco8472, w_eco8473, w_eco8474, w_eco8475, w_eco8476, w_eco8477, w_eco8478, w_eco8479, w_eco8480, w_eco8481, w_eco8482, w_eco8483, w_eco8484, w_eco8485, w_eco8486, w_eco8487, w_eco8488, w_eco8489, w_eco8490, w_eco8491, w_eco8492, w_eco8493, w_eco8494, w_eco8495, w_eco8496, w_eco8497, w_eco8498, w_eco8499, w_eco8500, w_eco8501, w_eco8502, w_eco8503, w_eco8504, w_eco8505, w_eco8506, w_eco8507, w_eco8508, w_eco8509, w_eco8510, w_eco8511, w_eco8512, w_eco8513, w_eco8514, w_eco8515, w_eco8516, w_eco8517, w_eco8518, w_eco8519, w_eco8520, w_eco8521, w_eco8522, w_eco8523, w_eco8524, w_eco8525, w_eco8526, w_eco8527, w_eco8528, w_eco8529, w_eco8530, w_eco8531, w_eco8532, w_eco8533, w_eco8534, w_eco8535, w_eco8536, w_eco8537, w_eco8538, w_eco8539, w_eco8540, w_eco8541, w_eco8542, w_eco8543, w_eco8544, w_eco8545, w_eco8546, w_eco8547, w_eco8548, w_eco8549, w_eco8550, w_eco8551, w_eco8552, w_eco8553, w_eco8554, w_eco8555, w_eco8556, w_eco8557, w_eco8558, w_eco8559, w_eco8560, w_eco8561, w_eco8562, w_eco8563, w_eco8564, w_eco8565, w_eco8566, w_eco8567, w_eco8568, w_eco8569, w_eco8570, w_eco8571, w_eco8572, w_eco8573, w_eco8574, w_eco8575, w_eco8576, w_eco8577, w_eco8578, w_eco8579, w_eco8580, w_eco8581, w_eco8582, w_eco8583, w_eco8584, w_eco8585, w_eco8586, w_eco8587, w_eco8588, w_eco8589, w_eco8590, w_eco8591, w_eco8592, w_eco8593, w_eco8594, w_eco8595, w_eco8596, w_eco8597, w_eco8598, w_eco8599, w_eco8600, w_eco8601, w_eco8602, w_eco8603, w_eco8604, w_eco8605, w_eco8606, w_eco8607, w_eco8608, w_eco8609, w_eco8610, w_eco8611, w_eco8612, w_eco8613, w_eco8614, w_eco8615, w_eco8616, w_eco8617, w_eco8618, w_eco8619, w_eco8620, w_eco8621, w_eco8622, w_eco8623, w_eco8624, w_eco8625, w_eco8626, w_eco8627, w_eco8628, w_eco8629, w_eco8630, w_eco8631, w_eco8632, w_eco8633, w_eco8634, w_eco8635, w_eco8636, w_eco8637, w_eco8638, w_eco8639, w_eco8640, w_eco8641, w_eco8642, w_eco8643, w_eco8644, w_eco8645, w_eco8646, w_eco8647, w_eco8648, w_eco8649, w_eco8650, w_eco8651, w_eco8652, w_eco8653, w_eco8654, w_eco8655, w_eco8656, w_eco8657, w_eco8658, w_eco8659, w_eco8660, w_eco8661, w_eco8662, w_eco8663, w_eco8664, w_eco8665, w_eco8666, w_eco8667, w_eco8668, w_eco8669, w_eco8670, w_eco8671, w_eco8672, w_eco8673, w_eco8674, w_eco8675, w_eco8676, w_eco8677, w_eco8678, w_eco8679, w_eco8680, w_eco8681, w_eco8682, w_eco8683, w_eco8684, w_eco8685, w_eco8686, w_eco8687, w_eco8688, w_eco8689, w_eco8690, w_eco8691, w_eco8692, w_eco8693, w_eco8694, w_eco8695, w_eco8696, w_eco8697, w_eco8698, w_eco8699, w_eco8700, w_eco8701, w_eco8702, w_eco8703, w_eco8704, w_eco8705, w_eco8706, w_eco8707, w_eco8708, w_eco8709, w_eco8710, w_eco8711, w_eco8712, w_eco8713, w_eco8714, w_eco8715, w_eco8716, w_eco8717, w_eco8718, w_eco8719, w_eco8720, w_eco8721, w_eco8722, w_eco8723, w_eco8724, w_eco8725, w_eco8726, w_eco8727, w_eco8728, w_eco8729, w_eco8730, w_eco8731, w_eco8732, w_eco8733, w_eco8734, w_eco8735, w_eco8736, w_eco8737, w_eco8738, w_eco8739, w_eco8740, w_eco8741, w_eco8742, w_eco8743, w_eco8744, w_eco8745, w_eco8746, w_eco8747, w_eco8748, w_eco8749, w_eco8750, w_eco8751, w_eco8752, w_eco8753, w_eco8754, w_eco8755, w_eco8756, w_eco8757, w_eco8758, w_eco8759, w_eco8760, w_eco8761, w_eco8762, w_eco8763, w_eco8764, w_eco8765, w_eco8766, w_eco8767, w_eco8768, w_eco8769, w_eco8770, w_eco8771, w_eco8772, w_eco8773, w_eco8774, w_eco8775, w_eco8776, w_eco8777, w_eco8778, w_eco8779, w_eco8780, w_eco8781, w_eco8782, w_eco8783, w_eco8784, w_eco8785, w_eco8786, w_eco8787, w_eco8788, w_eco8789, w_eco8790, w_eco8791, w_eco8792, w_eco8793, w_eco8794, w_eco8795, w_eco8796, w_eco8797, w_eco8798, w_eco8799, w_eco8800, w_eco8801, w_eco8802, w_eco8803, w_eco8804, w_eco8805, w_eco8806, w_eco8807, w_eco8808, w_eco8809, w_eco8810, w_eco8811, w_eco8812, w_eco8813, w_eco8814, w_eco8815, w_eco8816, w_eco8817, w_eco8818, w_eco8819, w_eco8820, w_eco8821, w_eco8822, w_eco8823, w_eco8824, w_eco8825, w_eco8826, w_eco8827, w_eco8828, w_eco8829, w_eco8830, w_eco8831, w_eco8832, w_eco8833, w_eco8834, w_eco8835, w_eco8836, w_eco8837, w_eco8838, w_eco8839, w_eco8840, w_eco8841, w_eco8842, w_eco8843, w_eco8844, w_eco8845, w_eco8846, w_eco8847, w_eco8848, w_eco8849, w_eco8850, w_eco8851, w_eco8852, w_eco8853, w_eco8854, w_eco8855, w_eco8856, w_eco8857, w_eco8858, w_eco8859, w_eco8860, w_eco8861, w_eco8862, w_eco8863, w_eco8864, w_eco8865, w_eco8866, w_eco8867, w_eco8868, w_eco8869, w_eco8870, w_eco8871, w_eco8872, w_eco8873, w_eco8874, w_eco8875, w_eco8876, w_eco8877, w_eco8878, w_eco8879, w_eco8880, w_eco8881, w_eco8882, w_eco8883, w_eco8884, w_eco8885, w_eco8886, w_eco8887, w_eco8888, w_eco8889, w_eco8890, w_eco8891, w_eco8892, w_eco8893, w_eco8894, w_eco8895, w_eco8896, w_eco8897, w_eco8898, w_eco8899, w_eco8900, w_eco8901, w_eco8902, w_eco8903, w_eco8904, w_eco8905, w_eco8906, w_eco8907, w_eco8908, w_eco8909, w_eco8910, w_eco8911, w_eco8912, w_eco8913, w_eco8914, w_eco8915, w_eco8916, w_eco8917, w_eco8918, w_eco8919, w_eco8920, w_eco8921, w_eco8922, w_eco8923, w_eco8924, w_eco8925, w_eco8926, w_eco8927, w_eco8928, w_eco8929, w_eco8930, w_eco8931, w_eco8932, w_eco8933, w_eco8934, w_eco8935, w_eco8936, w_eco8937, w_eco8938, w_eco8939, w_eco8940, w_eco8941, w_eco8942, w_eco8943, w_eco8944, w_eco8945, w_eco8946, w_eco8947, w_eco8948, w_eco8949, w_eco8950, w_eco8951, w_eco8952, w_eco8953, w_eco8954, w_eco8955, w_eco8956, w_eco8957, w_eco8958, w_eco8959, w_eco8960, w_eco8961, w_eco8962, w_eco8963, w_eco8964, w_eco8965, w_eco8966, w_eco8967, w_eco8968, w_eco8969, w_eco8970, w_eco8971, w_eco8972, w_eco8973, w_eco8974, w_eco8975, w_eco8976, w_eco8977, w_eco8978, w_eco8979, w_eco8980, w_eco8981, w_eco8982, w_eco8983, w_eco8984, w_eco8985, w_eco8986, w_eco8987, w_eco8988, w_eco8989, w_eco8990, w_eco8991, w_eco8992, w_eco8993, w_eco8994, w_eco8995, w_eco8996, w_eco8997, w_eco8998, w_eco8999, w_eco9000, w_eco9001, w_eco9002, w_eco9003, w_eco9004, w_eco9005, w_eco9006, w_eco9007, w_eco9008, w_eco9009, w_eco9010, w_eco9011, w_eco9012, w_eco9013, w_eco9014, w_eco9015, w_eco9016, w_eco9017, w_eco9018, w_eco9019, w_eco9020, w_eco9021, w_eco9022, w_eco9023, w_eco9024, w_eco9025, w_eco9026, w_eco9027, w_eco9028, w_eco9029, w_eco9030, w_eco9031, w_eco9032, w_eco9033, w_eco9034, w_eco9035, w_eco9036, w_eco9037, w_eco9038, w_eco9039, w_eco9040, w_eco9041, w_eco9042, w_eco9043, w_eco9044, w_eco9045, w_eco9046, w_eco9047, w_eco9048, w_eco9049, w_eco9050, w_eco9051, w_eco9052, w_eco9053, w_eco9054, w_eco9055, w_eco9056, w_eco9057, w_eco9058, w_eco9059, w_eco9060, w_eco9061, w_eco9062, w_eco9063, w_eco9064, w_eco9065, w_eco9066, w_eco9067, w_eco9068, w_eco9069, w_eco9070, w_eco9071, w_eco9072, w_eco9073, w_eco9074, w_eco9075, w_eco9076, w_eco9077, w_eco9078, w_eco9079, w_eco9080, w_eco9081, w_eco9082, w_eco9083, w_eco9084, w_eco9085, w_eco9086, w_eco9087, w_eco9088, w_eco9089, w_eco9090, w_eco9091, w_eco9092, w_eco9093, w_eco9094, w_eco9095, w_eco9096, w_eco9097, w_eco9098, w_eco9099, w_eco9100, w_eco9101, w_eco9102, w_eco9103, w_eco9104, w_eco9105, w_eco9106, w_eco9107, w_eco9108, w_eco9109, w_eco9110, w_eco9111, w_eco9112, w_eco9113, w_eco9114, w_eco9115, w_eco9116, w_eco9117, w_eco9118, w_eco9119, w_eco9120, w_eco9121, w_eco9122, w_eco9123, w_eco9124, w_eco9125, w_eco9126, w_eco9127, w_eco9128, w_eco9129, w_eco9130, w_eco9131, w_eco9132, w_eco9133, w_eco9134, w_eco9135, w_eco9136, w_eco9137, w_eco9138, w_eco9139, w_eco9140, w_eco9141, w_eco9142, w_eco9143, w_eco9144, w_eco9145, w_eco9146, w_eco9147, w_eco9148, w_eco9149, w_eco9150, w_eco9151, w_eco9152, w_eco9153, w_eco9154, w_eco9155, w_eco9156, w_eco9157, w_eco9158, w_eco9159, w_eco9160, w_eco9161, w_eco9162, w_eco9163, w_eco9164, w_eco9165, w_eco9166, w_eco9167, w_eco9168, w_eco9169, w_eco9170, w_eco9171, w_eco9172, w_eco9173, w_eco9174, w_eco9175, w_eco9176, w_eco9177, w_eco9178, w_eco9179, w_eco9180, w_eco9181, w_eco9182, w_eco9183, w_eco9184, w_eco9185, w_eco9186, w_eco9187, w_eco9188, w_eco9189, w_eco9190, w_eco9191, w_eco9192, w_eco9193, w_eco9194, w_eco9195, w_eco9196, w_eco9197, w_eco9198, w_eco9199, w_eco9200, w_eco9201, w_eco9202, w_eco9203, w_eco9204, w_eco9205, w_eco9206, w_eco9207, w_eco9208, w_eco9209, w_eco9210, w_eco9211, w_eco9212, w_eco9213, w_eco9214, w_eco9215, w_eco9216, w_eco9217, w_eco9218, w_eco9219, w_eco9220, w_eco9221, w_eco9222, w_eco9223, w_eco9224, w_eco9225, w_eco9226, w_eco9227, w_eco9228, w_eco9229, w_eco9230, w_eco9231, w_eco9232, w_eco9233, w_eco9234, w_eco9235, w_eco9236, w_eco9237, w_eco9238, w_eco9239, w_eco9240, w_eco9241, w_eco9242, w_eco9243, w_eco9244, w_eco9245, w_eco9246, w_eco9247, w_eco9248, w_eco9249, w_eco9250, w_eco9251, w_eco9252, w_eco9253, w_eco9254, w_eco9255, w_eco9256, w_eco9257, w_eco9258, w_eco9259, w_eco9260, w_eco9261, w_eco9262, w_eco9263, w_eco9264, w_eco9265, w_eco9266, w_eco9267, w_eco9268, w_eco9269, w_eco9270, w_eco9271, w_eco9272, w_eco9273, w_eco9274, w_eco9275, w_eco9276, w_eco9277, w_eco9278, w_eco9279, w_eco9280, w_eco9281, w_eco9282, w_eco9283, w_eco9284, w_eco9285, w_eco9286, w_eco9287, w_eco9288, w_eco9289, w_eco9290, w_eco9291, w_eco9292, w_eco9293, w_eco9294, w_eco9295, w_eco9296, w_eco9297, w_eco9298, w_eco9299, w_eco9300, w_eco9301, w_eco9302, w_eco9303, w_eco9304, w_eco9305, w_eco9306, w_eco9307, w_eco9308, w_eco9309, w_eco9310, w_eco9311, w_eco9312, w_eco9313, w_eco9314, w_eco9315, w_eco9316, w_eco9317, w_eco9318, w_eco9319, w_eco9320, w_eco9321, w_eco9322, w_eco9323, w_eco9324, w_eco9325, w_eco9326, w_eco9327, w_eco9328, w_eco9329, w_eco9330, w_eco9331, w_eco9332, w_eco9333, w_eco9334, w_eco9335, w_eco9336, w_eco9337, w_eco9338, w_eco9339, w_eco9340, w_eco9341, w_eco9342, w_eco9343, w_eco9344, w_eco9345, w_eco9346, w_eco9347, w_eco9348, w_eco9349, w_eco9350, w_eco9351, w_eco9352, w_eco9353, w_eco9354, w_eco9355, w_eco9356, w_eco9357, w_eco9358, w_eco9359, w_eco9360, w_eco9361, w_eco9362, w_eco9363, w_eco9364, w_eco9365, w_eco9366, w_eco9367, w_eco9368, w_eco9369, w_eco9370, w_eco9371, w_eco9372, w_eco9373, w_eco9374, w_eco9375, w_eco9376, w_eco9377, w_eco9378, w_eco9379, w_eco9380, w_eco9381, w_eco9382, w_eco9383, w_eco9384, w_eco9385, w_eco9386, w_eco9387, w_eco9388, w_eco9389, w_eco9390, w_eco9391, w_eco9392, w_eco9393, w_eco9394, w_eco9395, w_eco9396, w_eco9397, w_eco9398, w_eco9399, w_eco9400, w_eco9401, w_eco9402, w_eco9403, w_eco9404, w_eco9405, w_eco9406, w_eco9407, w_eco9408, w_eco9409, w_eco9410, w_eco9411, w_eco9412, w_eco9413, w_eco9414, w_eco9415, w_eco9416, w_eco9417, w_eco9418, w_eco9419, w_eco9420, w_eco9421, w_eco9422, w_eco9423, w_eco9424, w_eco9425, w_eco9426, w_eco9427, w_eco9428, w_eco9429, w_eco9430, w_eco9431, w_eco9432, w_eco9433, w_eco9434, w_eco9435, w_eco9436, w_eco9437, w_eco9438, w_eco9439, w_eco9440, w_eco9441, w_eco9442, w_eco9443, w_eco9444, w_eco9445, w_eco9446, w_eco9447, w_eco9448, w_eco9449, w_eco9450, w_eco9451, w_eco9452, w_eco9453, w_eco9454, w_eco9455, w_eco9456, w_eco9457, w_eco9458, w_eco9459, w_eco9460, w_eco9461, w_eco9462, w_eco9463, w_eco9464, w_eco9465, w_eco9466, w_eco9467, w_eco9468, w_eco9469, w_eco9470, w_eco9471, w_eco9472, w_eco9473, w_eco9474, w_eco9475, w_eco9476, w_eco9477, w_eco9478, w_eco9479, w_eco9480, w_eco9481, w_eco9482, w_eco9483, w_eco9484, w_eco9485, w_eco9486, w_eco9487, w_eco9488, w_eco9489, w_eco9490, w_eco9491, w_eco9492, w_eco9493, w_eco9494, w_eco9495, w_eco9496, w_eco9497, w_eco9498, w_eco9499, w_eco9500, w_eco9501, w_eco9502, w_eco9503, w_eco9504, w_eco9505, w_eco9506, w_eco9507, w_eco9508, w_eco9509, w_eco9510, w_eco9511, w_eco9512, w_eco9513, w_eco9514, w_eco9515, w_eco9516, w_eco9517, w_eco9518, w_eco9519, w_eco9520, w_eco9521, w_eco9522, w_eco9523, w_eco9524, w_eco9525, w_eco9526, w_eco9527, w_eco9528, w_eco9529, w_eco9530, w_eco9531, w_eco9532, w_eco9533, w_eco9534, w_eco9535, w_eco9536, w_eco9537, w_eco9538, w_eco9539, w_eco9540, w_eco9541, w_eco9542, w_eco9543, w_eco9544, w_eco9545, w_eco9546, w_eco9547, w_eco9548, w_eco9549, w_eco9550, w_eco9551, w_eco9552, w_eco9553, w_eco9554, w_eco9555, w_eco9556, w_eco9557, w_eco9558, w_eco9559, w_eco9560, w_eco9561, w_eco9562, w_eco9563, w_eco9564, w_eco9565, w_eco9566, w_eco9567, w_eco9568, w_eco9569, w_eco9570, w_eco9571, w_eco9572, w_eco9573, w_eco9574, w_eco9575, w_eco9576, w_eco9577, w_eco9578, w_eco9579, w_eco9580, w_eco9581, w_eco9582, w_eco9583, w_eco9584);
	xor _ECO_out6(cnt[2], sub_wire6, w_eco9585);
	assign w_eco9586 = rst;
	and _ECO_9587(w_eco9587, Tsync[1], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9588(w_eco9588, Tsync[1], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_9589(w_eco9589, Tsync[1], !prev_cnt[6], ena, !prev_state[3], prev_state[1]);
	and _ECO_9590(w_eco9590, Tsync[1], !prev_cnt[6], ena, !prev_state[0]);
	and _ECO_9591(w_eco9591, !Tsync[6], Tsync[1], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_9592(w_eco9592, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_state[1]);
	and _ECO_9593(w_eco9593, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_state[3], !prev_state[2]);
	and _ECO_9594(w_eco9594, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_state[4], !prev_state[2]);
	and _ECO_9595(w_eco9595, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[11], !ena);
	and _ECO_9596(w_eco9596, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[11], !ena);
	and _ECO_9597(w_eco9597, Tgate[1], prev_cnt[0], prev_cnt[1], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9598(w_eco9598, Tgate[1], !prev_cnt[0], !prev_cnt[1], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9599(w_eco9599, Tgate[1], prev_cnt[0], prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9600(w_eco9600, Tgate[1], !prev_cnt[0], !prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9601(w_eco9601, Tgate[1], prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, !prev_state[3], prev_state[1]);
	and _ECO_9602(w_eco9602, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_9603(w_eco9603, Tgate[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, !prev_state[3], prev_state[1]);
	and _ECO_9604(w_eco9604, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_9605(w_eco9605, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[15], !ena);
	and _ECO_9606(w_eco9606, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[15], !ena);
	and _ECO_9607(w_eco9607, !Tsync[6], Tgate[1], prev_cnt[0], prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_9608(w_eco9608, !Tsync[6], prev_cnt[0], prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9609(w_eco9609, !Tsync[6], Tgate[1], !prev_cnt[0], !prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_9610(w_eco9610, !Tsync[6], !prev_cnt[0], !prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9611(w_eco9611, prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9612(w_eco9612, Tgate[1], prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_9613(w_eco9613, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_9614(w_eco9614, Tgate[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0]);
	and _ECO_9615(w_eco9615, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_9616(w_eco9616, !Tsync[6], prev_cnt[0], prev_cnt[1], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_9617(w_eco9617, !Tsync[6], !prev_cnt[0], !prev_cnt[1], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_9618(w_eco9618, prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9619(w_eco9619, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_9620(w_eco9620, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_9621(w_eco9621, !Tsync[1], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9622(w_eco9622, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_9623(w_eco9623, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_9624(w_eco9624, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[6], prev_state[1]);
	and _ECO_9625(w_eco9625, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[6], prev_state[1]);
	and _ECO_9626(w_eco9626, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9627(w_eco9627, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9628(w_eco9628, !Tsync[6], prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[0]);
	and _ECO_9629(w_eco9629, !Tsync[6], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[0]);
	and _ECO_9630(w_eco9630, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_9631(w_eco9631, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_9632(w_eco9632, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9633(w_eco9633, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9634(w_eco9634, prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9635(w_eco9635, !prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9636(w_eco9636, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9637(w_eco9637, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9638(w_eco9638, prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9639(w_eco9639, !prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9640(w_eco9640, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_9641(w_eco9641, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_9642(w_eco9642, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_9643(w_eco9643, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[6], !prev_state[4], !prev_state[2]);
	and _ECO_9644(w_eco9644, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9645(w_eco9645, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9646(w_eco9646, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9647(w_eco9647, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9648(w_eco9648, !prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9649(w_eco9649, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[9], !ena);
	and _ECO_9650(w_eco9650, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[9], !ena);
	and _ECO_9651(w_eco9651, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9652(w_eco9652, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9653(w_eco9653, !prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9654(w_eco9654, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_9655(w_eco9655, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[6], !prev_state[3], prev_state[0]);
	and _ECO_9656(w_eco9656, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9657(w_eco9657, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9658(w_eco9658, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_9659(w_eco9659, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_9660(w_eco9660, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9661(w_eco9661, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9662(w_eco9662, Tgdel[1], prev_cnt[0], prev_cnt[1], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9663(w_eco9663, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[6], !ena);
	and _ECO_9664(w_eco9664, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[6], !ena);
	and _ECO_9665(w_eco9665, Tgdel[1], prev_cnt[0], prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9666(w_eco9666, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9667(w_eco9667, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9668(w_eco9668, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[8], !ena);
	and _ECO_9669(w_eco9669, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[8], !ena);
	and _ECO_9670(w_eco9670, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9671(w_eco9671, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9672(w_eco9672, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9673(w_eco9673, prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9674(w_eco9674, Tgdel[1], !prev_cnt[0], !prev_cnt[1], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9675(w_eco9675, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9676(w_eco9676, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9677(w_eco9677, prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9678(w_eco9678, Tgdel[1], !prev_cnt[0], !prev_cnt[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9679(w_eco9679, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9680(w_eco9680, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_9681(w_eco9681, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_9682(w_eco9682, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9683(w_eco9683, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9684(w_eco9684, !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[10], !ena);
	and _ECO_9685(w_eco9685, !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[10], !ena);
	and _ECO_9686(w_eco9686, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9687(w_eco9687, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9688(w_eco9688, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[6], prev_state[0]);
	and _ECO_9689(w_eco9689, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[6], prev_state[0]);
	and _ECO_9690(w_eco9690, prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9691(w_eco9691, !prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9692(w_eco9692, prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9693(w_eco9693, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_9694(w_eco9694, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_9695(w_eco9695, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_9696(w_eco9696, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9697(w_eco9697, !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], !ena);
	and _ECO_9698(w_eco9698, !Tgate[1], !Tgdel[1], !Tsync[1], !prev_cnt[0], prev_cnt[1], !ena);
	and _ECO_9699(w_eco9699, !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], !ena);
	and _ECO_9700(w_eco9700, !Tgate[1], !Tgdel[1], !Tsync[1], prev_cnt[0], !prev_cnt[1], !ena);
	and _ECO_9701(w_eco9701, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9702(w_eco9702, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9703(w_eco9703, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9704(w_eco9704, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9705(w_eco9705, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9706(w_eco9706, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9707(w_eco9707, Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9708(w_eco9708, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9709(w_eco9709, !prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9710(w_eco9710, Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_9711(w_eco9711, Tgdel[1], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_9712(w_eco9712, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9713(w_eco9713, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9714(w_eco9714, prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9715(w_eco9715, !prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9716(w_eco9716, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_9717(w_eco9717, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_9718(w_eco9718, !Tsync[6], Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_9719(w_eco9719, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9720(w_eco9720, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_9721(w_eco9721, !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], !ena);
	and _ECO_9722(w_eco9722, !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], !ena);
	and _ECO_9723(w_eco9723, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9724(w_eco9724, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9725(w_eco9725, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9726(w_eco9726, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9727(w_eco9727, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9728(w_eco9728, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9729(w_eco9729, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9730(w_eco9730, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9731(w_eco9731, Tgdel[1], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_9732(w_eco9732, Tgdel[1], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_9733(w_eco9733, prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9734(w_eco9734, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9735(w_eco9735, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9736(w_eco9736, Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9737(w_eco9737, !prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9738(w_eco9738, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9739(w_eco9739, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9740(w_eco9740, prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9741(w_eco9741, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9742(w_eco9742, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_9743(w_eco9743, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_state[3], prev_state[0]);
	and _ECO_9744(w_eco9744, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_9745(w_eco9745, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_state[3], prev_state[0]);
	and _ECO_9746(w_eco9746, !Tsync[6], Tgdel[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_9747(w_eco9747, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9748(w_eco9748, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9749(w_eco9749, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9750(w_eco9750, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9751(w_eco9751, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9752(w_eco9752, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9753(w_eco9753, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9754(w_eco9754, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9755(w_eco9755, Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9756(w_eco9756, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9757(w_eco9757, Tgdel[1], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_9758(w_eco9758, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9759(w_eco9759, Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_9760(w_eco9760, Tgdel[1], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_9761(w_eco9761, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9762(w_eco9762, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9763(w_eco9763, Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_9764(w_eco9764, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9765(w_eco9765, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9766(w_eco9766, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9767(w_eco9767, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9768(w_eco9768, Tgdel[1], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_9769(w_eco9769, Tgdel[1], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_9770(w_eco9770, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9771(w_eco9771, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9772(w_eco9772, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_9773(w_eco9773, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9774(w_eco9774, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9775(w_eco9775, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9776(w_eco9776, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9777(w_eco9777, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9778(w_eco9778, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9779(w_eco9779, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9780(w_eco9780, Tgate[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9781(w_eco9781, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_9782(w_eco9782, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_9783(w_eco9783, !Tsync[6], Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_9784(w_eco9784, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9785(w_eco9785, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9786(w_eco9786, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9787(w_eco9787, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9788(w_eco9788, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9789(w_eco9789, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9790(w_eco9790, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9791(w_eco9791, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9792(w_eco9792, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9793(w_eco9793, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9794(w_eco9794, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9795(w_eco9795, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9796(w_eco9796, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9797(w_eco9797, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9798(w_eco9798, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9799(w_eco9799, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9800(w_eco9800, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9801(w_eco9801, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9802(w_eco9802, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9803(w_eco9803, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9804(w_eco9804, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9805(w_eco9805, Tgdel[1], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_9806(w_eco9806, Tgdel[1], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_9807(w_eco9807, !prev_cnt[0], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9808(w_eco9808, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9809(w_eco9809, Tgdel[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_9810(w_eco9810, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9811(w_eco9811, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9812(w_eco9812, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9813(w_eco9813, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9814(w_eco9814, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9815(w_eco9815, Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9816(w_eco9816, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9817(w_eco9817, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9818(w_eco9818, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9819(w_eco9819, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9820(w_eco9820, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9821(w_eco9821, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_9822(w_eco9822, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9823(w_eco9823, Tsync[6], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9824(w_eco9824, Tsync[6], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9825(w_eco9825, prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9826(w_eco9826, !prev_cnt[0], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9827(w_eco9827, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9828(w_eco9828, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9829(w_eco9829, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9830(w_eco9830, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9831(w_eco9831, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9832(w_eco9832, Tgdel[1], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9833(w_eco9833, !Tsync[6], Tgdel[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_9834(w_eco9834, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9835(w_eco9835, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9836(w_eco9836, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9837(w_eco9837, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9838(w_eco9838, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9839(w_eco9839, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9840(w_eco9840, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9841(w_eco9841, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9842(w_eco9842, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9843(w_eco9843, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_9844(w_eco9844, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9845(w_eco9845, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9846(w_eco9846, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9847(w_eco9847, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9848(w_eco9848, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9849(w_eco9849, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9850(w_eco9850, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9851(w_eco9851, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9852(w_eco9852, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9853(w_eco9853, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9854(w_eco9854, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9855(w_eco9855, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9856(w_eco9856, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9857(w_eco9857, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9858(w_eco9858, Tgdel[1], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_9859(w_eco9859, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9860(w_eco9860, !prev_cnt[0], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9861(w_eco9861, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9862(w_eco9862, Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_9863(w_eco9863, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9864(w_eco9864, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9865(w_eco9865, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9866(w_eco9866, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9867(w_eco9867, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9868(w_eco9868, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9869(w_eco9869, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9870(w_eco9870, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9871(w_eco9871, Tgdel[1], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_9872(w_eco9872, Tgdel[1], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_9873(w_eco9873, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9874(w_eco9874, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_9875(w_eco9875, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9876(w_eco9876, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_9877(w_eco9877, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9878(w_eco9878, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9879(w_eco9879, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], !prev_cnt[0], prev_cnt[1], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9880(w_eco9880, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9881(w_eco9881, Tsync[6], !Tgate[1], !Tgdel[1], !Tsync[1], prev_cnt[0], !prev_cnt[1], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9882(w_eco9882, !prev_cnt[0], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9883(w_eco9883, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9884(w_eco9884, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9885(w_eco9885, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9886(w_eco9886, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9887(w_eco9887, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9888(w_eco9888, Tgate[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9889(w_eco9889, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9890(w_eco9890, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9891(w_eco9891, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9892(w_eco9892, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9893(w_eco9893, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9894(w_eco9894, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9895(w_eco9895, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9896(w_eco9896, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9897(w_eco9897, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9898(w_eco9898, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9899(w_eco9899, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9900(w_eco9900, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9901(w_eco9901, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9902(w_eco9902, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9903(w_eco9903, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9904(w_eco9904, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9905(w_eco9905, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9906(w_eco9906, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9907(w_eco9907, !prev_cnt[0], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9908(w_eco9908, Tgdel[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_9909(w_eco9909, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9910(w_eco9910, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9911(w_eco9911, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9912(w_eco9912, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9913(w_eco9913, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9914(w_eco9914, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_9915(w_eco9915, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9916(w_eco9916, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_9917(w_eco9917, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_9918(w_eco9918, Tsync[6], !Tsync[1], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9919(w_eco9919, Tsync[6], !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_9920(w_eco9920, !prev_cnt[0], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9921(w_eco9921, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9922(w_eco9922, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9923(w_eco9923, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9924(w_eco9924, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9925(w_eco9925, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9926(w_eco9926, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9927(w_eco9927, Tgdel[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_9928(w_eco9928, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9929(w_eco9929, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9930(w_eco9930, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9931(w_eco9931, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9932(w_eco9932, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9933(w_eco9933, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9934(w_eco9934, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9935(w_eco9935, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9936(w_eco9936, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9937(w_eco9937, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9938(w_eco9938, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9939(w_eco9939, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9940(w_eco9940, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9941(w_eco9941, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9942(w_eco9942, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9943(w_eco9943, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9944(w_eco9944, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9945(w_eco9945, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9946(w_eco9946, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9947(w_eco9947, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9948(w_eco9948, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9949(w_eco9949, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9950(w_eco9950, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9951(w_eco9951, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9952(w_eco9952, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9953(w_eco9953, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9954(w_eco9954, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9955(w_eco9955, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9956(w_eco9956, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_9957(w_eco9957, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_9958(w_eco9958, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9959(w_eco9959, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9960(w_eco9960, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9961(w_eco9961, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9962(w_eco9962, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9963(w_eco9963, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9964(w_eco9964, prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_9965(w_eco9965, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_9966(w_eco9966, !prev_cnt[0], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_9967(w_eco9967, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9968(w_eco9968, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9969(w_eco9969, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9970(w_eco9970, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9971(w_eco9971, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9972(w_eco9972, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9973(w_eco9973, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9974(w_eco9974, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9975(w_eco9975, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9976(w_eco9976, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9977(w_eco9977, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9978(w_eco9978, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9979(w_eco9979, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_9980(w_eco9980, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9981(w_eco9981, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9982(w_eco9982, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9983(w_eco9983, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9984(w_eco9984, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9985(w_eco9985, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9986(w_eco9986, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9987(w_eco9987, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9988(w_eco9988, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9989(w_eco9989, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9990(w_eco9990, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9991(w_eco9991, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_9992(w_eco9992, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9993(w_eco9993, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_9994(w_eco9994, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9995(w_eco9995, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9996(w_eco9996, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_9997(w_eco9997, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_9998(w_eco9998, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_9999(w_eco9999, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10000(w_eco10000, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10001(w_eco10001, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10002(w_eco10002, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_10003(w_eco10003, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_10004(w_eco10004, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_10005(w_eco10005, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_10006(w_eco10006, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10007(w_eco10007, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10008(w_eco10008, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10009(w_eco10009, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10010(w_eco10010, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10011(w_eco10011, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10012(w_eco10012, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10013(w_eco10013, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10014(w_eco10014, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10015(w_eco10015, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10016(w_eco10016, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10017(w_eco10017, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10018(w_eco10018, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10019(w_eco10019, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10020(w_eco10020, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10021(w_eco10021, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10022(w_eco10022, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10023(w_eco10023, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10024(w_eco10024, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10025(w_eco10025, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10026(w_eco10026, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10027(w_eco10027, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10028(w_eco10028, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10029(w_eco10029, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10030(w_eco10030, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10031(w_eco10031, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10032(w_eco10032, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10033(w_eco10033, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10034(w_eco10034, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10035(w_eco10035, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10036(w_eco10036, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10037(w_eco10037, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10038(w_eco10038, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10039(w_eco10039, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10040(w_eco10040, !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10041(w_eco10041, prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10042(w_eco10042, !Tsync[6], Tsync[1], !prev_cnt[6], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10043(w_eco10043, !prev_cnt[14], prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_10044(w_eco10044, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_10045(w_eco10045, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10046(w_eco10046, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10047(w_eco10047, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10048(w_eco10048, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10049(w_eco10049, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10050(w_eco10050, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10051(w_eco10051, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10052(w_eco10052, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10053(w_eco10053, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10054(w_eco10054, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10055(w_eco10055, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10056(w_eco10056, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10057(w_eco10057, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10058(w_eco10058, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10059(w_eco10059, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10060(w_eco10060, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10061(w_eco10061, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10062(w_eco10062, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10063(w_eco10063, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10064(w_eco10064, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10065(w_eco10065, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10066(w_eco10066, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10067(w_eco10067, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10068(w_eco10068, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10069(w_eco10069, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10070(w_eco10070, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10071(w_eco10071, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10072(w_eco10072, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10073(w_eco10073, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10074(w_eco10074, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10075(w_eco10075, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10076(w_eco10076, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10077(w_eco10077, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10078(w_eco10078, !Tsync[6], Tsync[1], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10079(w_eco10079, !Tsync[6], Tsync[1], !prev_cnt[6], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10080(w_eco10080, !Tsync[6], Tsync[1], !prev_cnt[6], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10081(w_eco10081, !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_10082(w_eco10082, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10083(w_eco10083, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10084(w_eco10084, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10085(w_eco10085, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10086(w_eco10086, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10087(w_eco10087, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10088(w_eco10088, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10089(w_eco10089, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10090(w_eco10090, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10091(w_eco10091, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10092(w_eco10092, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10093(w_eco10093, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10094(w_eco10094, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10095(w_eco10095, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10096(w_eco10096, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10097(w_eco10097, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10098(w_eco10098, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10099(w_eco10099, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10100(w_eco10100, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10101(w_eco10101, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10102(w_eco10102, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10103(w_eco10103, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10104(w_eco10104, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10105(w_eco10105, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10106(w_eco10106, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10107(w_eco10107, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10108(w_eco10108, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10109(w_eco10109, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10110(w_eco10110, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10111(w_eco10111, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10112(w_eco10112, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10113(w_eco10113, !Tsync[6], Tsync[1], !prev_cnt[6], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10114(w_eco10114, Tsync[1], !prev_cnt[6], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10115(w_eco10115, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10116(w_eco10116, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10117(w_eco10117, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10118(w_eco10118, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10119(w_eco10119, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10120(w_eco10120, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10121(w_eco10121, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10122(w_eco10122, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10123(w_eco10123, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10124(w_eco10124, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10125(w_eco10125, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10126(w_eco10126, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10127(w_eco10127, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10128(w_eco10128, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10129(w_eco10129, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10130(w_eco10130, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10131(w_eco10131, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10132(w_eco10132, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10133(w_eco10133, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10134(w_eco10134, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10135(w_eco10135, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10136(w_eco10136, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10137(w_eco10137, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10138(w_eco10138, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10139(w_eco10139, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10140(w_eco10140, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10141(w_eco10141, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10142(w_eco10142, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10143(w_eco10143, !Tsync[6], Tsync[1], !prev_cnt[6], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10144(w_eco10144, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_10145(w_eco10145, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10146(w_eco10146, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10147(w_eco10147, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10148(w_eco10148, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10149(w_eco10149, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10150(w_eco10150, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10151(w_eco10151, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10152(w_eco10152, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10153(w_eco10153, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10154(w_eco10154, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10155(w_eco10155, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10156(w_eco10156, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10157(w_eco10157, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10158(w_eco10158, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10159(w_eco10159, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10160(w_eco10160, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10161(w_eco10161, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10162(w_eco10162, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10163(w_eco10163, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10164(w_eco10164, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10165(w_eco10165, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10166(w_eco10166, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10167(w_eco10167, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10168(w_eco10168, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10169(w_eco10169, prev_cnt[0], prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10170(w_eco10170, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10171(w_eco10171, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10172(w_eco10172, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10173(w_eco10173, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10174(w_eco10174, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10175(w_eco10175, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10176(w_eco10176, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10177(w_eco10177, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10178(w_eco10178, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10179(w_eco10179, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10180(w_eco10180, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10181(w_eco10181, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10182(w_eco10182, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10183(w_eco10183, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10184(w_eco10184, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10185(w_eco10185, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10186(w_eco10186, !prev_cnt[0], !prev_cnt[1], !prev_cnt[6], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10187(w_eco10187, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10188(w_eco10188, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10189(w_eco10189, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10190(w_eco10190, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10191(w_eco10191, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10192(w_eco10192, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10193(w_eco10193, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10194(w_eco10194, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10195(w_eco10195, Tsync[6], !prev_cnt[0], prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10196(w_eco10196, Tsync[6], prev_cnt[0], !prev_cnt[1], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10197(w_eco10197, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10198(w_eco10198, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10199(w_eco10199, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10200(w_eco10200, Tsync[6], !Tgate[1], !Tgdel[1], !prev_cnt[0], prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10201(w_eco10201, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10202(w_eco10202, Tsync[6], !Tgate[1], !Tgdel[1], prev_cnt[0], !prev_cnt[1], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10203(w_eco10203, Tsync[6], !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10204(w_eco10204, Tsync[6], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_10205(w_eco10205, w_eco9586, w_eco9587, w_eco9588, w_eco9589, w_eco9590, w_eco9591, w_eco9592, w_eco9593, w_eco9594, w_eco9595, w_eco9596, w_eco9597, w_eco9598, w_eco9599, w_eco9600, w_eco9601, w_eco9602, w_eco9603, w_eco9604, w_eco9605, w_eco9606, w_eco9607, w_eco9608, w_eco9609, w_eco9610, w_eco9611, w_eco9612, w_eco9613, w_eco9614, w_eco9615, w_eco9616, w_eco9617, w_eco9618, w_eco9619, w_eco9620, w_eco9621, w_eco9622, w_eco9623, w_eco9624, w_eco9625, w_eco9626, w_eco9627, w_eco9628, w_eco9629, w_eco9630, w_eco9631, w_eco9632, w_eco9633, w_eco9634, w_eco9635, w_eco9636, w_eco9637, w_eco9638, w_eco9639, w_eco9640, w_eco9641, w_eco9642, w_eco9643, w_eco9644, w_eco9645, w_eco9646, w_eco9647, w_eco9648, w_eco9649, w_eco9650, w_eco9651, w_eco9652, w_eco9653, w_eco9654, w_eco9655, w_eco9656, w_eco9657, w_eco9658, w_eco9659, w_eco9660, w_eco9661, w_eco9662, w_eco9663, w_eco9664, w_eco9665, w_eco9666, w_eco9667, w_eco9668, w_eco9669, w_eco9670, w_eco9671, w_eco9672, w_eco9673, w_eco9674, w_eco9675, w_eco9676, w_eco9677, w_eco9678, w_eco9679, w_eco9680, w_eco9681, w_eco9682, w_eco9683, w_eco9684, w_eco9685, w_eco9686, w_eco9687, w_eco9688, w_eco9689, w_eco9690, w_eco9691, w_eco9692, w_eco9693, w_eco9694, w_eco9695, w_eco9696, w_eco9697, w_eco9698, w_eco9699, w_eco9700, w_eco9701, w_eco9702, w_eco9703, w_eco9704, w_eco9705, w_eco9706, w_eco9707, w_eco9708, w_eco9709, w_eco9710, w_eco9711, w_eco9712, w_eco9713, w_eco9714, w_eco9715, w_eco9716, w_eco9717, w_eco9718, w_eco9719, w_eco9720, w_eco9721, w_eco9722, w_eco9723, w_eco9724, w_eco9725, w_eco9726, w_eco9727, w_eco9728, w_eco9729, w_eco9730, w_eco9731, w_eco9732, w_eco9733, w_eco9734, w_eco9735, w_eco9736, w_eco9737, w_eco9738, w_eco9739, w_eco9740, w_eco9741, w_eco9742, w_eco9743, w_eco9744, w_eco9745, w_eco9746, w_eco9747, w_eco9748, w_eco9749, w_eco9750, w_eco9751, w_eco9752, w_eco9753, w_eco9754, w_eco9755, w_eco9756, w_eco9757, w_eco9758, w_eco9759, w_eco9760, w_eco9761, w_eco9762, w_eco9763, w_eco9764, w_eco9765, w_eco9766, w_eco9767, w_eco9768, w_eco9769, w_eco9770, w_eco9771, w_eco9772, w_eco9773, w_eco9774, w_eco9775, w_eco9776, w_eco9777, w_eco9778, w_eco9779, w_eco9780, w_eco9781, w_eco9782, w_eco9783, w_eco9784, w_eco9785, w_eco9786, w_eco9787, w_eco9788, w_eco9789, w_eco9790, w_eco9791, w_eco9792, w_eco9793, w_eco9794, w_eco9795, w_eco9796, w_eco9797, w_eco9798, w_eco9799, w_eco9800, w_eco9801, w_eco9802, w_eco9803, w_eco9804, w_eco9805, w_eco9806, w_eco9807, w_eco9808, w_eco9809, w_eco9810, w_eco9811, w_eco9812, w_eco9813, w_eco9814, w_eco9815, w_eco9816, w_eco9817, w_eco9818, w_eco9819, w_eco9820, w_eco9821, w_eco9822, w_eco9823, w_eco9824, w_eco9825, w_eco9826, w_eco9827, w_eco9828, w_eco9829, w_eco9830, w_eco9831, w_eco9832, w_eco9833, w_eco9834, w_eco9835, w_eco9836, w_eco9837, w_eco9838, w_eco9839, w_eco9840, w_eco9841, w_eco9842, w_eco9843, w_eco9844, w_eco9845, w_eco9846, w_eco9847, w_eco9848, w_eco9849, w_eco9850, w_eco9851, w_eco9852, w_eco9853, w_eco9854, w_eco9855, w_eco9856, w_eco9857, w_eco9858, w_eco9859, w_eco9860, w_eco9861, w_eco9862, w_eco9863, w_eco9864, w_eco9865, w_eco9866, w_eco9867, w_eco9868, w_eco9869, w_eco9870, w_eco9871, w_eco9872, w_eco9873, w_eco9874, w_eco9875, w_eco9876, w_eco9877, w_eco9878, w_eco9879, w_eco9880, w_eco9881, w_eco9882, w_eco9883, w_eco9884, w_eco9885, w_eco9886, w_eco9887, w_eco9888, w_eco9889, w_eco9890, w_eco9891, w_eco9892, w_eco9893, w_eco9894, w_eco9895, w_eco9896, w_eco9897, w_eco9898, w_eco9899, w_eco9900, w_eco9901, w_eco9902, w_eco9903, w_eco9904, w_eco9905, w_eco9906, w_eco9907, w_eco9908, w_eco9909, w_eco9910, w_eco9911, w_eco9912, w_eco9913, w_eco9914, w_eco9915, w_eco9916, w_eco9917, w_eco9918, w_eco9919, w_eco9920, w_eco9921, w_eco9922, w_eco9923, w_eco9924, w_eco9925, w_eco9926, w_eco9927, w_eco9928, w_eco9929, w_eco9930, w_eco9931, w_eco9932, w_eco9933, w_eco9934, w_eco9935, w_eco9936, w_eco9937, w_eco9938, w_eco9939, w_eco9940, w_eco9941, w_eco9942, w_eco9943, w_eco9944, w_eco9945, w_eco9946, w_eco9947, w_eco9948, w_eco9949, w_eco9950, w_eco9951, w_eco9952, w_eco9953, w_eco9954, w_eco9955, w_eco9956, w_eco9957, w_eco9958, w_eco9959, w_eco9960, w_eco9961, w_eco9962, w_eco9963, w_eco9964, w_eco9965, w_eco9966, w_eco9967, w_eco9968, w_eco9969, w_eco9970, w_eco9971, w_eco9972, w_eco9973, w_eco9974, w_eco9975, w_eco9976, w_eco9977, w_eco9978, w_eco9979, w_eco9980, w_eco9981, w_eco9982, w_eco9983, w_eco9984, w_eco9985, w_eco9986, w_eco9987, w_eco9988, w_eco9989, w_eco9990, w_eco9991, w_eco9992, w_eco9993, w_eco9994, w_eco9995, w_eco9996, w_eco9997, w_eco9998, w_eco9999, w_eco10000, w_eco10001, w_eco10002, w_eco10003, w_eco10004, w_eco10005, w_eco10006, w_eco10007, w_eco10008, w_eco10009, w_eco10010, w_eco10011, w_eco10012, w_eco10013, w_eco10014, w_eco10015, w_eco10016, w_eco10017, w_eco10018, w_eco10019, w_eco10020, w_eco10021, w_eco10022, w_eco10023, w_eco10024, w_eco10025, w_eco10026, w_eco10027, w_eco10028, w_eco10029, w_eco10030, w_eco10031, w_eco10032, w_eco10033, w_eco10034, w_eco10035, w_eco10036, w_eco10037, w_eco10038, w_eco10039, w_eco10040, w_eco10041, w_eco10042, w_eco10043, w_eco10044, w_eco10045, w_eco10046, w_eco10047, w_eco10048, w_eco10049, w_eco10050, w_eco10051, w_eco10052, w_eco10053, w_eco10054, w_eco10055, w_eco10056, w_eco10057, w_eco10058, w_eco10059, w_eco10060, w_eco10061, w_eco10062, w_eco10063, w_eco10064, w_eco10065, w_eco10066, w_eco10067, w_eco10068, w_eco10069, w_eco10070, w_eco10071, w_eco10072, w_eco10073, w_eco10074, w_eco10075, w_eco10076, w_eco10077, w_eco10078, w_eco10079, w_eco10080, w_eco10081, w_eco10082, w_eco10083, w_eco10084, w_eco10085, w_eco10086, w_eco10087, w_eco10088, w_eco10089, w_eco10090, w_eco10091, w_eco10092, w_eco10093, w_eco10094, w_eco10095, w_eco10096, w_eco10097, w_eco10098, w_eco10099, w_eco10100, w_eco10101, w_eco10102, w_eco10103, w_eco10104, w_eco10105, w_eco10106, w_eco10107, w_eco10108, w_eco10109, w_eco10110, w_eco10111, w_eco10112, w_eco10113, w_eco10114, w_eco10115, w_eco10116, w_eco10117, w_eco10118, w_eco10119, w_eco10120, w_eco10121, w_eco10122, w_eco10123, w_eco10124, w_eco10125, w_eco10126, w_eco10127, w_eco10128, w_eco10129, w_eco10130, w_eco10131, w_eco10132, w_eco10133, w_eco10134, w_eco10135, w_eco10136, w_eco10137, w_eco10138, w_eco10139, w_eco10140, w_eco10141, w_eco10142, w_eco10143, w_eco10144, w_eco10145, w_eco10146, w_eco10147, w_eco10148, w_eco10149, w_eco10150, w_eco10151, w_eco10152, w_eco10153, w_eco10154, w_eco10155, w_eco10156, w_eco10157, w_eco10158, w_eco10159, w_eco10160, w_eco10161, w_eco10162, w_eco10163, w_eco10164, w_eco10165, w_eco10166, w_eco10167, w_eco10168, w_eco10169, w_eco10170, w_eco10171, w_eco10172, w_eco10173, w_eco10174, w_eco10175, w_eco10176, w_eco10177, w_eco10178, w_eco10179, w_eco10180, w_eco10181, w_eco10182, w_eco10183, w_eco10184, w_eco10185, w_eco10186, w_eco10187, w_eco10188, w_eco10189, w_eco10190, w_eco10191, w_eco10192, w_eco10193, w_eco10194, w_eco10195, w_eco10196, w_eco10197, w_eco10198, w_eco10199, w_eco10200, w_eco10201, w_eco10202, w_eco10203, w_eco10204);
	xor _ECO_out7(cnt[1], sub_wire7, w_eco10205);
	assign w_eco10206 = rst;
	and _ECO_10207(w_eco10207, Tsync[0], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10208(w_eco10208, Tsync[0], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10209(w_eco10209, Tsync[0], !prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_10210(w_eco10210, Tsync[0], !prev_cnt[7], ena, !prev_state[0]);
	and _ECO_10211(w_eco10211, !Tsync[0], prev_cnt[0], prev_cnt[11], !ena);
	and _ECO_10212(w_eco10212, Tgdel[0], !prev_cnt[0], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10213(w_eco10213, Tsync[0], !Tsync[7], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_10214(w_eco10214, Tgdel[0], !prev_cnt[0], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10215(w_eco10215, !prev_cnt[0], !prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_10216(w_eco10216, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_state[1]);
	and _ECO_10217(w_eco10217, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_10218(w_eco10218, !Tsync[0], prev_cnt[0], prev_cnt[15], !ena);
	and _ECO_10219(w_eco10219, Tgdel[0], !Tsync[7], !prev_cnt[0], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10220(w_eco10220, !Tsync[7], !prev_cnt[0], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10221(w_eco10221, !Tsync[7], !prev_cnt[0], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10222(w_eco10222, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_state[3], !prev_state[2]);
	and _ECO_10223(w_eco10223, !prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_10224(w_eco10224, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], prev_state[1]);
	and _ECO_10225(w_eco10225, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_state[4], !prev_state[2]);
	and _ECO_10226(w_eco10226, !prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10227(w_eco10227, !Tsync[7], !prev_cnt[0], !prev_cnt[7], ena, prev_state[0]);
	and _ECO_10228(w_eco10228, Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10229(w_eco10229, !prev_cnt[0], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10230(w_eco10230, !prev_cnt[0], !prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_10231(w_eco10231, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10232(w_eco10232, !prev_cnt[0], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10233(w_eco10233, !prev_cnt[0], !prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_10234(w_eco10234, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_10235(w_eco10235, !Tsync[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10236(w_eco10236, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], prev_state[1]);
	and _ECO_10237(w_eco10237, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10238(w_eco10238, !Tsync[0], prev_cnt[0], prev_cnt[9], !ena);
	and _ECO_10239(w_eco10239, Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10240(w_eco10240, !prev_cnt[0], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10241(w_eco10241, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10242(w_eco10242, !prev_cnt[0], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10243(w_eco10243, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_10244(w_eco10244, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_10245(w_eco10245, !Tsync[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10246(w_eco10246, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10247(w_eco10247, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_10248(w_eco10248, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10249(w_eco10249, !Tsync[0], prev_cnt[0], prev_cnt[6], !ena);
	and _ECO_10250(w_eco10250, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_10251(w_eco10251, !Tgdel[0], !Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10252(w_eco10252, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10253(w_eco10253, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], prev_state[1]);
	and _ECO_10254(w_eco10254, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_10255(w_eco10255, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10256(w_eco10256, !Tsync[0], prev_cnt[0], prev_cnt[8], !ena);
	and _ECO_10257(w_eco10257, Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10258(w_eco10258, Tgate[0], !prev_cnt[0], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10259(w_eco10259, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10260(w_eco10260, Tgate[0], !prev_cnt[0], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10261(w_eco10261, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_10262(w_eco10262, !Tsync[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10263(w_eco10263, !Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], prev_state[1]);
	and _ECO_10264(w_eco10264, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10265(w_eco10265, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10266(w_eco10266, !Tsync[0], prev_cnt[0], prev_cnt[10], !ena);
	and _ECO_10267(w_eco10267, Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10268(w_eco10268, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10269(w_eco10269, !prev_cnt[0], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10270(w_eco10270, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10271(w_eco10271, !prev_cnt[0], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10272(w_eco10272, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], prev_state[3], prev_state[0]);
	and _ECO_10273(w_eco10273, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_10274(w_eco10274, !Tsync[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10275(w_eco10275, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10276(w_eco10276, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], prev_state[1]);
	and _ECO_10277(w_eco10277, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_10278(w_eco10278, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10279(w_eco10279, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10280(w_eco10280, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10281(w_eco10281, !prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_10282(w_eco10282, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[12], !ena);
	and _ECO_10283(w_eco10283, !Tgate[0], !Tgdel[0], !Tsync[0], prev_cnt[0], !ena);
	and _ECO_10284(w_eco10284, Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10285(w_eco10285, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10286(w_eco10286, Tgdel[0], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10287(w_eco10287, !prev_cnt[0], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10288(w_eco10288, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10289(w_eco10289, Tgdel[0], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10290(w_eco10290, !prev_cnt[0], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10291(w_eco10291, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_10292(w_eco10292, !Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], !prev_state[4], !prev_state[2]);
	and _ECO_10293(w_eco10293, !Tsync[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10294(w_eco10294, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10295(w_eco10295, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10296(w_eco10296, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], prev_state[1]);
	and _ECO_10297(w_eco10297, Tgdel[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_10298(w_eco10298, !Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], !prev_state[3], prev_state[0]);
	and _ECO_10299(w_eco10299, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10300(w_eco10300, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10301(w_eco10301, !prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_10302(w_eco10302, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[13], !ena);
	and _ECO_10303(w_eco10303, Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10304(w_eco10304, Tgdel[0], !Tsync[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10305(w_eco10305, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10306(w_eco10306, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10307(w_eco10307, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10308(w_eco10308, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10309(w_eco10309, !prev_cnt[0], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10310(w_eco10310, Tgdel[0], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_10311(w_eco10311, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10312(w_eco10312, Tgdel[0], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_10313(w_eco10313, prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10314(w_eco10314, !prev_cnt[0], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10315(w_eco10315, Tgdel[0], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_10316(w_eco10316, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_10317(w_eco10317, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_10318(w_eco10318, Tgdel[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_10319(w_eco10319, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10320(w_eco10320, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10321(w_eco10321, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], prev_state[1]);
	and _ECO_10322(w_eco10322, !Tgate[0], !Tgdel[0], !Tsync[0], prev_cnt[0], prev_cnt[7], prev_state[1]);
	and _ECO_10323(w_eco10323, Tgate[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_10324(w_eco10324, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_10325(w_eco10325, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10326(w_eco10326, Tgdel[0], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10327(w_eco10327, prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10328(w_eco10328, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10329(w_eco10329, Tgdel[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10330(w_eco10330, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10331(w_eco10331, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10332(w_eco10332, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10333(w_eco10333, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10334(w_eco10334, !Tsync[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10335(w_eco10335, Tgdel[0], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_10336(w_eco10336, Tgdel[0], !Tsync[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_10337(w_eco10337, Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10338(w_eco10338, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10339(w_eco10339, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10340(w_eco10340, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10341(w_eco10341, !Tgate[0], !Tgdel[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10342(w_eco10342, Tgate[0], !Tsync[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10343(w_eco10343, Tgdel[0], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10344(w_eco10344, prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10345(w_eco10345, Tgate[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_10346(w_eco10346, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10347(w_eco10347, !Tgate[0], !Tgdel[0], !Tsync[0], Tsync[7], prev_cnt[0], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10348(w_eco10348, Tgate[0], !Tsync[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10349(w_eco10349, prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10350(w_eco10350, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_10351(w_eco10351, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_10352(w_eco10352, !Tgate[0], !Tgdel[0], !Tsync[0], Tsync[7], prev_cnt[0], prev_state[3], prev_state[0]);
	and _ECO_10353(w_eco10353, !Tsync[0], !prev_cnt[14], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10354(w_eco10354, prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10355(w_eco10355, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10356(w_eco10356, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10357(w_eco10357, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10358(w_eco10358, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10359(w_eco10359, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10360(w_eco10360, Tgate[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10361(w_eco10361, !prev_cnt[0], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10362(w_eco10362, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], prev_state[1]);
	and _ECO_10363(w_eco10363, Tgdel[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_10364(w_eco10364, !Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_10365(w_eco10365, Tgdel[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10366(w_eco10366, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10367(w_eco10367, !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10368(w_eco10368, prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10369(w_eco10369, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10370(w_eco10370, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10371(w_eco10371, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10372(w_eco10372, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10373(w_eco10373, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10374(w_eco10374, Tgate[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10375(w_eco10375, Tgdel[0], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_10376(w_eco10376, Tgate[0], !Tsync[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_10377(w_eco10377, !Tgate[0], Tgdel[0], !Tsync[0], prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[0]);
	and _ECO_10378(w_eco10378, Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10379(w_eco10379, Tgdel[0], !Tsync[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10380(w_eco10380, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10381(w_eco10381, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10382(w_eco10382, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10383(w_eco10383, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10384(w_eco10384, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10385(w_eco10385, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10386(w_eco10386, !prev_cnt[14], !prev_cnt[0], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10387(w_eco10387, Tgdel[0], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_10388(w_eco10388, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10389(w_eco10389, Tgdel[0], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_10390(w_eco10390, !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10391(w_eco10391, prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10392(w_eco10392, Tgate[0], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10393(w_eco10393, !prev_cnt[0], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10394(w_eco10394, !prev_cnt[14], !prev_cnt[0], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10395(w_eco10395, Tgdel[0], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_10396(w_eco10396, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_10397(w_eco10397, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_10398(w_eco10398, !Tgate[0], !Tgdel[0], !Tsync[0], prev_cnt[0], prev_cnt[7], !prev_state[4], !prev_state[2]);
	and _ECO_10399(w_eco10399, prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10400(w_eco10400, Tgdel[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_10401(w_eco10401, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10402(w_eco10402, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10403(w_eco10403, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10404(w_eco10404, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10405(w_eco10405, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10406(w_eco10406, Tgate[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_10407(w_eco10407, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_10408(w_eco10408, !Tgate[0], !Tgdel[0], !Tsync[0], prev_cnt[0], prev_cnt[7], !prev_state[3], prev_state[0]);
	and _ECO_10409(w_eco10409, Tgdel[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10410(w_eco10410, !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10411(w_eco10411, prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10412(w_eco10412, !Tgate[0], !Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_10413(w_eco10413, !prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_10414(w_eco10414, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10415(w_eco10415, Tgdel[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10416(w_eco10416, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10417(w_eco10417, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10418(w_eco10418, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10419(w_eco10419, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10420(w_eco10420, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10421(w_eco10421, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10422(w_eco10422, !Tsync[0], !prev_cnt[14], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10423(w_eco10423, !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10424(w_eco10424, prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10425(w_eco10425, Tgdel[0], !Tsync[7], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_10426(w_eco10426, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10427(w_eco10427, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10428(w_eco10428, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10429(w_eco10429, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10430(w_eco10430, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10431(w_eco10431, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10432(w_eco10432, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10433(w_eco10433, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10434(w_eco10434, Tgate[0], !Tsync[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10435(w_eco10435, Tgate[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_10436(w_eco10436, Tgate[0], !Tsync[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10437(w_eco10437, !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10438(w_eco10438, prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10439(w_eco10439, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_10440(w_eco10440, !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10441(w_eco10441, prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10442(w_eco10442, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10443(w_eco10443, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10444(w_eco10444, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10445(w_eco10445, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10446(w_eco10446, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10447(w_eco10447, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10448(w_eco10448, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10449(w_eco10449, Tgate[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10450(w_eco10450, !prev_cnt[14], !prev_cnt[0], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10451(w_eco10451, !Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_10452(w_eco10452, !prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_10453(w_eco10453, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10454(w_eco10454, !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10455(w_eco10455, prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10456(w_eco10456, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10457(w_eco10457, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10458(w_eco10458, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10459(w_eco10459, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10460(w_eco10460, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10461(w_eco10461, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10462(w_eco10462, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10463(w_eco10463, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10464(w_eco10464, Tgate[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10465(w_eco10465, Tgdel[0], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_10466(w_eco10466, Tgate[0], !Tsync[7], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_10467(w_eco10467, !Tgate[0], Tgdel[0], !Tsync[0], prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[0]);
	and _ECO_10468(w_eco10468, !prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_10469(w_eco10469, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10470(w_eco10470, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10471(w_eco10471, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10472(w_eco10472, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10473(w_eco10473, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10474(w_eco10474, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10475(w_eco10475, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10476(w_eco10476, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10477(w_eco10477, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10478(w_eco10478, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10479(w_eco10479, !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10480(w_eco10480, prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10481(w_eco10481, Tgate[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10482(w_eco10482, !prev_cnt[14], !prev_cnt[0], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10483(w_eco10483, !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10484(w_eco10484, prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10485(w_eco10485, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10486(w_eco10486, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10487(w_eco10487, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10488(w_eco10488, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10489(w_eco10489, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10490(w_eco10490, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10491(w_eco10491, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10492(w_eco10492, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10493(w_eco10493, Tgdel[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10494(w_eco10494, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10495(w_eco10495, !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10496(w_eco10496, prev_cnt[14], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10497(w_eco10497, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10498(w_eco10498, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10499(w_eco10499, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10500(w_eco10500, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10501(w_eco10501, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10502(w_eco10502, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10503(w_eco10503, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10504(w_eco10504, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10505(w_eco10505, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10506(w_eco10506, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10507(w_eco10507, Tgdel[0], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_10508(w_eco10508, !prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_10509(w_eco10509, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10510(w_eco10510, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10511(w_eco10511, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10512(w_eco10512, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10513(w_eco10513, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10514(w_eco10514, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10515(w_eco10515, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10516(w_eco10516, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10517(w_eco10517, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10518(w_eco10518, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10519(w_eco10519, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10520(w_eco10520, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10521(w_eco10521, !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10522(w_eco10522, prev_cnt[14], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10523(w_eco10523, !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10524(w_eco10524, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10525(w_eco10525, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10526(w_eco10526, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10527(w_eco10527, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10528(w_eco10528, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10529(w_eco10529, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10530(w_eco10530, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10531(w_eco10531, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10532(w_eco10532, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10533(w_eco10533, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10534(w_eco10534, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10535(w_eco10535, !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10536(w_eco10536, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10537(w_eco10537, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10538(w_eco10538, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10539(w_eco10539, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10540(w_eco10540, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10541(w_eco10541, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10542(w_eco10542, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10543(w_eco10543, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10544(w_eco10544, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10545(w_eco10545, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10546(w_eco10546, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10547(w_eco10547, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10548(w_eco10548, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10549(w_eco10549, !prev_cnt[14], !prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_10550(w_eco10550, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10551(w_eco10551, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10552(w_eco10552, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10553(w_eco10553, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10554(w_eco10554, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10555(w_eco10555, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10556(w_eco10556, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10557(w_eco10557, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10558(w_eco10558, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10559(w_eco10559, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10560(w_eco10560, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10561(w_eco10561, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10562(w_eco10562, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10563(w_eco10563, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10564(w_eco10564, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_10565(w_eco10565, !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10566(w_eco10566, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_10567(w_eco10567, !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10568(w_eco10568, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10569(w_eco10569, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10570(w_eco10570, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10571(w_eco10571, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10572(w_eco10572, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10573(w_eco10573, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10574(w_eco10574, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10575(w_eco10575, Tsync[0], !Tsync[7], !prev_cnt[7], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10576(w_eco10576, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10577(w_eco10577, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10578(w_eco10578, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10579(w_eco10579, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10580(w_eco10580, !Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10581(w_eco10581, !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10582(w_eco10582, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10583(w_eco10583, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10584(w_eco10584, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10585(w_eco10585, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10586(w_eco10586, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10587(w_eco10587, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10588(w_eco10588, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10589(w_eco10589, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10590(w_eco10590, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10591(w_eco10591, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10592(w_eco10592, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10593(w_eco10593, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10594(w_eco10594, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10595(w_eco10595, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10596(w_eco10596, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10597(w_eco10597, !prev_cnt[14], !prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_10598(w_eco10598, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10599(w_eco10599, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10600(w_eco10600, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10601(w_eco10601, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10602(w_eco10602, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10603(w_eco10603, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10604(w_eco10604, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10605(w_eco10605, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10606(w_eco10606, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10607(w_eco10607, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10608(w_eco10608, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10609(w_eco10609, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10610(w_eco10610, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10611(w_eco10611, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10612(w_eco10612, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10613(w_eco10613, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10614(w_eco10614, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10615(w_eco10615, !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10616(w_eco10616, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10617(w_eco10617, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10618(w_eco10618, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10619(w_eco10619, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10620(w_eco10620, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10621(w_eco10621, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10622(w_eco10622, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10623(w_eco10623, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10624(w_eco10624, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10625(w_eco10625, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10626(w_eco10626, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10627(w_eco10627, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10628(w_eco10628, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10629(w_eco10629, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10630(w_eco10630, Tsync[0], !Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10631(w_eco10631, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10632(w_eco10632, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10633(w_eco10633, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10634(w_eco10634, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10635(w_eco10635, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10636(w_eco10636, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10637(w_eco10637, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10638(w_eco10638, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10639(w_eco10639, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10640(w_eco10640, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10641(w_eco10641, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10642(w_eco10642, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10643(w_eco10643, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10644(w_eco10644, Tsync[0], !Tsync[7], !prev_cnt[7], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10645(w_eco10645, Tsync[0], !Tsync[7], !prev_cnt[7], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10646(w_eco10646, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10647(w_eco10647, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10648(w_eco10648, !Tgate[0], !Tgdel[0], !Tsync[0], Tsync[7], prev_cnt[0], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10649(w_eco10649, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10650(w_eco10650, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10651(w_eco10651, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10652(w_eco10652, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10653(w_eco10653, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10654(w_eco10654, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10655(w_eco10655, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10656(w_eco10656, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10657(w_eco10657, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10658(w_eco10658, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10659(w_eco10659, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10660(w_eco10660, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10661(w_eco10661, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10662(w_eco10662, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10663(w_eco10663, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10664(w_eco10664, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10665(w_eco10665, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10666(w_eco10666, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10667(w_eco10667, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10668(w_eco10668, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10669(w_eco10669, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10670(w_eco10670, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10671(w_eco10671, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10672(w_eco10672, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10673(w_eco10673, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10674(w_eco10674, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10675(w_eco10675, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10676(w_eco10676, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10677(w_eco10677, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10678(w_eco10678, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10679(w_eco10679, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10680(w_eco10680, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10681(w_eco10681, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10682(w_eco10682, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10683(w_eco10683, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10684(w_eco10684, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10685(w_eco10685, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10686(w_eco10686, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10687(w_eco10687, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10688(w_eco10688, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10689(w_eco10689, Tsync[0], !Tsync[7], !prev_cnt[7], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10690(w_eco10690, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10691(w_eco10691, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10692(w_eco10692, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_10693(w_eco10693, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10694(w_eco10694, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10695(w_eco10695, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10696(w_eco10696, !Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10697(w_eco10697, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10698(w_eco10698, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10699(w_eco10699, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10700(w_eco10700, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10701(w_eco10701, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10702(w_eco10702, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10703(w_eco10703, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10704(w_eco10704, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10705(w_eco10705, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10706(w_eco10706, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10707(w_eco10707, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10708(w_eco10708, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10709(w_eco10709, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10710(w_eco10710, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10711(w_eco10711, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10712(w_eco10712, Tsync[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10713(w_eco10713, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10714(w_eco10714, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10715(w_eco10715, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10716(w_eco10716, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10717(w_eco10717, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10718(w_eco10718, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10719(w_eco10719, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10720(w_eco10720, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10721(w_eco10721, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10722(w_eco10722, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10723(w_eco10723, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10724(w_eco10724, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10725(w_eco10725, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10726(w_eco10726, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10727(w_eco10727, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10728(w_eco10728, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10729(w_eco10729, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10730(w_eco10730, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10731(w_eco10731, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10732(w_eco10732, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10733(w_eco10733, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10734(w_eco10734, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10735(w_eco10735, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10736(w_eco10736, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10737(w_eco10737, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10738(w_eco10738, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10739(w_eco10739, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10740(w_eco10740, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10741(w_eco10741, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10742(w_eco10742, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10743(w_eco10743, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10744(w_eco10744, Tsync[0], !Tsync[7], !prev_cnt[7], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10745(w_eco10745, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10746(w_eco10746, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10747(w_eco10747, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10748(w_eco10748, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10749(w_eco10749, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10750(w_eco10750, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10751(w_eco10751, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10752(w_eco10752, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10753(w_eco10753, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10754(w_eco10754, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10755(w_eco10755, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10756(w_eco10756, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10757(w_eco10757, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10758(w_eco10758, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10759(w_eco10759, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10760(w_eco10760, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10761(w_eco10761, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10762(w_eco10762, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10763(w_eco10763, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10764(w_eco10764, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10765(w_eco10765, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10766(w_eco10766, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10767(w_eco10767, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10768(w_eco10768, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10769(w_eco10769, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10770(w_eco10770, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10771(w_eco10771, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10772(w_eco10772, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10773(w_eco10773, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[6], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10774(w_eco10774, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10775(w_eco10775, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10776(w_eco10776, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10777(w_eco10777, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10778(w_eco10778, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10779(w_eco10779, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10780(w_eco10780, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10781(w_eco10781, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_10782(w_eco10782, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10783(w_eco10783, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10784(w_eco10784, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10785(w_eco10785, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10786(w_eco10786, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10787(w_eco10787, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10788(w_eco10788, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10789(w_eco10789, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10790(w_eco10790, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_10791(w_eco10791, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10792(w_eco10792, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10793(w_eco10793, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10794(w_eco10794, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10795(w_eco10795, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10796(w_eco10796, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10797(w_eco10797, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10798(w_eco10798, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10799(w_eco10799, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10800(w_eco10800, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10801(w_eco10801, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10802(w_eco10802, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10803(w_eco10803, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10804(w_eco10804, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10805(w_eco10805, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10806(w_eco10806, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10807(w_eco10807, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10808(w_eco10808, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10809(w_eco10809, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10810(w_eco10810, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10811(w_eco10811, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10812(w_eco10812, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10813(w_eco10813, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10814(w_eco10814, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10815(w_eco10815, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10816(w_eco10816, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10817(w_eco10817, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10818(w_eco10818, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10819(w_eco10819, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10820(w_eco10820, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10821(w_eco10821, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10822(w_eco10822, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10823(w_eco10823, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10824(w_eco10824, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10825(w_eco10825, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10826(w_eco10826, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10827(w_eco10827, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10828(w_eco10828, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10829(w_eco10829, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10830(w_eco10830, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10831(w_eco10831, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10832(w_eco10832, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10833(w_eco10833, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10834(w_eco10834, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10835(w_eco10835, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10836(w_eco10836, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10837(w_eco10837, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10838(w_eco10838, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10839(w_eco10839, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10840(w_eco10840, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10841(w_eco10841, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10842(w_eco10842, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10843(w_eco10843, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10844(w_eco10844, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10845(w_eco10845, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10846(w_eco10846, prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10847(w_eco10847, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10848(w_eco10848, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10849(w_eco10849, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10850(w_eco10850, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10851(w_eco10851, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10852(w_eco10852, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10853(w_eco10853, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10854(w_eco10854, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10855(w_eco10855, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10856(w_eco10856, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10857(w_eco10857, Tsync[0], Tsync[7], prev_cnt[0], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10858(w_eco10858, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10859(w_eco10859, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10860(w_eco10860, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10861(w_eco10861, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10862(w_eco10862, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10863(w_eco10863, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10864(w_eco10864, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10865(w_eco10865, Tsync[0], prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10866(w_eco10866, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10867(w_eco10867, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10868(w_eco10868, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10869(w_eco10869, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10870(w_eco10870, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10871(w_eco10871, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10872(w_eco10872, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10873(w_eco10873, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10874(w_eco10874, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10875(w_eco10875, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10876(w_eco10876, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10877(w_eco10877, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10878(w_eco10878, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10879(w_eco10879, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10880(w_eco10880, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10881(w_eco10881, !prev_cnt[0], !prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10882(w_eco10882, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10883(w_eco10883, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10884(w_eco10884, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10885(w_eco10885, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10886(w_eco10886, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10887(w_eco10887, !Tgate[0], !Tgdel[0], Tsync[0], Tsync[7], prev_cnt[0], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10888(w_eco10888, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10889(w_eco10889, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10890(w_eco10890, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10891(w_eco10891, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10892(w_eco10892, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10893(w_eco10893, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10894(w_eco10894, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10895(w_eco10895, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10896(w_eco10896, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10897(w_eco10897, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10898(w_eco10898, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10899(w_eco10899, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10900(w_eco10900, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10901(w_eco10901, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10902(w_eco10902, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10903(w_eco10903, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10904(w_eco10904, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10905(w_eco10905, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10906(w_eco10906, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10907(w_eco10907, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10908(w_eco10908, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_10909(w_eco10909, Tsync[0], prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10910(w_eco10910, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10911(w_eco10911, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10912(w_eco10912, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_10913(w_eco10913, !Tgate[0], !Tsync[0], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10914(w_eco10914, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10915(w_eco10915, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10916(w_eco10916, !Tgate[0], !Tgdel[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10917(w_eco10917, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10918(w_eco10918, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10919(w_eco10919, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10920(w_eco10920, !Tgate[0], !Tgdel[0], Tsync[0], prev_cnt[0], prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10921(w_eco10921, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_10922(w_eco10922, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10923(w_eco10923, Tsync[0], !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_10924(w_eco10924, !Tgate[0], !Tsync[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_10925(w_eco10925, w_eco10206, w_eco10207, w_eco10208, w_eco10209, w_eco10210, w_eco10211, w_eco10212, w_eco10213, w_eco10214, w_eco10215, w_eco10216, w_eco10217, w_eco10218, w_eco10219, w_eco10220, w_eco10221, w_eco10222, w_eco10223, w_eco10224, w_eco10225, w_eco10226, w_eco10227, w_eco10228, w_eco10229, w_eco10230, w_eco10231, w_eco10232, w_eco10233, w_eco10234, w_eco10235, w_eco10236, w_eco10237, w_eco10238, w_eco10239, w_eco10240, w_eco10241, w_eco10242, w_eco10243, w_eco10244, w_eco10245, w_eco10246, w_eco10247, w_eco10248, w_eco10249, w_eco10250, w_eco10251, w_eco10252, w_eco10253, w_eco10254, w_eco10255, w_eco10256, w_eco10257, w_eco10258, w_eco10259, w_eco10260, w_eco10261, w_eco10262, w_eco10263, w_eco10264, w_eco10265, w_eco10266, w_eco10267, w_eco10268, w_eco10269, w_eco10270, w_eco10271, w_eco10272, w_eco10273, w_eco10274, w_eco10275, w_eco10276, w_eco10277, w_eco10278, w_eco10279, w_eco10280, w_eco10281, w_eco10282, w_eco10283, w_eco10284, w_eco10285, w_eco10286, w_eco10287, w_eco10288, w_eco10289, w_eco10290, w_eco10291, w_eco10292, w_eco10293, w_eco10294, w_eco10295, w_eco10296, w_eco10297, w_eco10298, w_eco10299, w_eco10300, w_eco10301, w_eco10302, w_eco10303, w_eco10304, w_eco10305, w_eco10306, w_eco10307, w_eco10308, w_eco10309, w_eco10310, w_eco10311, w_eco10312, w_eco10313, w_eco10314, w_eco10315, w_eco10316, w_eco10317, w_eco10318, w_eco10319, w_eco10320, w_eco10321, w_eco10322, w_eco10323, w_eco10324, w_eco10325, w_eco10326, w_eco10327, w_eco10328, w_eco10329, w_eco10330, w_eco10331, w_eco10332, w_eco10333, w_eco10334, w_eco10335, w_eco10336, w_eco10337, w_eco10338, w_eco10339, w_eco10340, w_eco10341, w_eco10342, w_eco10343, w_eco10344, w_eco10345, w_eco10346, w_eco10347, w_eco10348, w_eco10349, w_eco10350, w_eco10351, w_eco10352, w_eco10353, w_eco10354, w_eco10355, w_eco10356, w_eco10357, w_eco10358, w_eco10359, w_eco10360, w_eco10361, w_eco10362, w_eco10363, w_eco10364, w_eco10365, w_eco10366, w_eco10367, w_eco10368, w_eco10369, w_eco10370, w_eco10371, w_eco10372, w_eco10373, w_eco10374, w_eco10375, w_eco10376, w_eco10377, w_eco10378, w_eco10379, w_eco10380, w_eco10381, w_eco10382, w_eco10383, w_eco10384, w_eco10385, w_eco10386, w_eco10387, w_eco10388, w_eco10389, w_eco10390, w_eco10391, w_eco10392, w_eco10393, w_eco10394, w_eco10395, w_eco10396, w_eco10397, w_eco10398, w_eco10399, w_eco10400, w_eco10401, w_eco10402, w_eco10403, w_eco10404, w_eco10405, w_eco10406, w_eco10407, w_eco10408, w_eco10409, w_eco10410, w_eco10411, w_eco10412, w_eco10413, w_eco10414, w_eco10415, w_eco10416, w_eco10417, w_eco10418, w_eco10419, w_eco10420, w_eco10421, w_eco10422, w_eco10423, w_eco10424, w_eco10425, w_eco10426, w_eco10427, w_eco10428, w_eco10429, w_eco10430, w_eco10431, w_eco10432, w_eco10433, w_eco10434, w_eco10435, w_eco10436, w_eco10437, w_eco10438, w_eco10439, w_eco10440, w_eco10441, w_eco10442, w_eco10443, w_eco10444, w_eco10445, w_eco10446, w_eco10447, w_eco10448, w_eco10449, w_eco10450, w_eco10451, w_eco10452, w_eco10453, w_eco10454, w_eco10455, w_eco10456, w_eco10457, w_eco10458, w_eco10459, w_eco10460, w_eco10461, w_eco10462, w_eco10463, w_eco10464, w_eco10465, w_eco10466, w_eco10467, w_eco10468, w_eco10469, w_eco10470, w_eco10471, w_eco10472, w_eco10473, w_eco10474, w_eco10475, w_eco10476, w_eco10477, w_eco10478, w_eco10479, w_eco10480, w_eco10481, w_eco10482, w_eco10483, w_eco10484, w_eco10485, w_eco10486, w_eco10487, w_eco10488, w_eco10489, w_eco10490, w_eco10491, w_eco10492, w_eco10493, w_eco10494, w_eco10495, w_eco10496, w_eco10497, w_eco10498, w_eco10499, w_eco10500, w_eco10501, w_eco10502, w_eco10503, w_eco10504, w_eco10505, w_eco10506, w_eco10507, w_eco10508, w_eco10509, w_eco10510, w_eco10511, w_eco10512, w_eco10513, w_eco10514, w_eco10515, w_eco10516, w_eco10517, w_eco10518, w_eco10519, w_eco10520, w_eco10521, w_eco10522, w_eco10523, w_eco10524, w_eco10525, w_eco10526, w_eco10527, w_eco10528, w_eco10529, w_eco10530, w_eco10531, w_eco10532, w_eco10533, w_eco10534, w_eco10535, w_eco10536, w_eco10537, w_eco10538, w_eco10539, w_eco10540, w_eco10541, w_eco10542, w_eco10543, w_eco10544, w_eco10545, w_eco10546, w_eco10547, w_eco10548, w_eco10549, w_eco10550, w_eco10551, w_eco10552, w_eco10553, w_eco10554, w_eco10555, w_eco10556, w_eco10557, w_eco10558, w_eco10559, w_eco10560, w_eco10561, w_eco10562, w_eco10563, w_eco10564, w_eco10565, w_eco10566, w_eco10567, w_eco10568, w_eco10569, w_eco10570, w_eco10571, w_eco10572, w_eco10573, w_eco10574, w_eco10575, w_eco10576, w_eco10577, w_eco10578, w_eco10579, w_eco10580, w_eco10581, w_eco10582, w_eco10583, w_eco10584, w_eco10585, w_eco10586, w_eco10587, w_eco10588, w_eco10589, w_eco10590, w_eco10591, w_eco10592, w_eco10593, w_eco10594, w_eco10595, w_eco10596, w_eco10597, w_eco10598, w_eco10599, w_eco10600, w_eco10601, w_eco10602, w_eco10603, w_eco10604, w_eco10605, w_eco10606, w_eco10607, w_eco10608, w_eco10609, w_eco10610, w_eco10611, w_eco10612, w_eco10613, w_eco10614, w_eco10615, w_eco10616, w_eco10617, w_eco10618, w_eco10619, w_eco10620, w_eco10621, w_eco10622, w_eco10623, w_eco10624, w_eco10625, w_eco10626, w_eco10627, w_eco10628, w_eco10629, w_eco10630, w_eco10631, w_eco10632, w_eco10633, w_eco10634, w_eco10635, w_eco10636, w_eco10637, w_eco10638, w_eco10639, w_eco10640, w_eco10641, w_eco10642, w_eco10643, w_eco10644, w_eco10645, w_eco10646, w_eco10647, w_eco10648, w_eco10649, w_eco10650, w_eco10651, w_eco10652, w_eco10653, w_eco10654, w_eco10655, w_eco10656, w_eco10657, w_eco10658, w_eco10659, w_eco10660, w_eco10661, w_eco10662, w_eco10663, w_eco10664, w_eco10665, w_eco10666, w_eco10667, w_eco10668, w_eco10669, w_eco10670, w_eco10671, w_eco10672, w_eco10673, w_eco10674, w_eco10675, w_eco10676, w_eco10677, w_eco10678, w_eco10679, w_eco10680, w_eco10681, w_eco10682, w_eco10683, w_eco10684, w_eco10685, w_eco10686, w_eco10687, w_eco10688, w_eco10689, w_eco10690, w_eco10691, w_eco10692, w_eco10693, w_eco10694, w_eco10695, w_eco10696, w_eco10697, w_eco10698, w_eco10699, w_eco10700, w_eco10701, w_eco10702, w_eco10703, w_eco10704, w_eco10705, w_eco10706, w_eco10707, w_eco10708, w_eco10709, w_eco10710, w_eco10711, w_eco10712, w_eco10713, w_eco10714, w_eco10715, w_eco10716, w_eco10717, w_eco10718, w_eco10719, w_eco10720, w_eco10721, w_eco10722, w_eco10723, w_eco10724, w_eco10725, w_eco10726, w_eco10727, w_eco10728, w_eco10729, w_eco10730, w_eco10731, w_eco10732, w_eco10733, w_eco10734, w_eco10735, w_eco10736, w_eco10737, w_eco10738, w_eco10739, w_eco10740, w_eco10741, w_eco10742, w_eco10743, w_eco10744, w_eco10745, w_eco10746, w_eco10747, w_eco10748, w_eco10749, w_eco10750, w_eco10751, w_eco10752, w_eco10753, w_eco10754, w_eco10755, w_eco10756, w_eco10757, w_eco10758, w_eco10759, w_eco10760, w_eco10761, w_eco10762, w_eco10763, w_eco10764, w_eco10765, w_eco10766, w_eco10767, w_eco10768, w_eco10769, w_eco10770, w_eco10771, w_eco10772, w_eco10773, w_eco10774, w_eco10775, w_eco10776, w_eco10777, w_eco10778, w_eco10779, w_eco10780, w_eco10781, w_eco10782, w_eco10783, w_eco10784, w_eco10785, w_eco10786, w_eco10787, w_eco10788, w_eco10789, w_eco10790, w_eco10791, w_eco10792, w_eco10793, w_eco10794, w_eco10795, w_eco10796, w_eco10797, w_eco10798, w_eco10799, w_eco10800, w_eco10801, w_eco10802, w_eco10803, w_eco10804, w_eco10805, w_eco10806, w_eco10807, w_eco10808, w_eco10809, w_eco10810, w_eco10811, w_eco10812, w_eco10813, w_eco10814, w_eco10815, w_eco10816, w_eco10817, w_eco10818, w_eco10819, w_eco10820, w_eco10821, w_eco10822, w_eco10823, w_eco10824, w_eco10825, w_eco10826, w_eco10827, w_eco10828, w_eco10829, w_eco10830, w_eco10831, w_eco10832, w_eco10833, w_eco10834, w_eco10835, w_eco10836, w_eco10837, w_eco10838, w_eco10839, w_eco10840, w_eco10841, w_eco10842, w_eco10843, w_eco10844, w_eco10845, w_eco10846, w_eco10847, w_eco10848, w_eco10849, w_eco10850, w_eco10851, w_eco10852, w_eco10853, w_eco10854, w_eco10855, w_eco10856, w_eco10857, w_eco10858, w_eco10859, w_eco10860, w_eco10861, w_eco10862, w_eco10863, w_eco10864, w_eco10865, w_eco10866, w_eco10867, w_eco10868, w_eco10869, w_eco10870, w_eco10871, w_eco10872, w_eco10873, w_eco10874, w_eco10875, w_eco10876, w_eco10877, w_eco10878, w_eco10879, w_eco10880, w_eco10881, w_eco10882, w_eco10883, w_eco10884, w_eco10885, w_eco10886, w_eco10887, w_eco10888, w_eco10889, w_eco10890, w_eco10891, w_eco10892, w_eco10893, w_eco10894, w_eco10895, w_eco10896, w_eco10897, w_eco10898, w_eco10899, w_eco10900, w_eco10901, w_eco10902, w_eco10903, w_eco10904, w_eco10905, w_eco10906, w_eco10907, w_eco10908, w_eco10909, w_eco10910, w_eco10911, w_eco10912, w_eco10913, w_eco10914, w_eco10915, w_eco10916, w_eco10917, w_eco10918, w_eco10919, w_eco10920, w_eco10921, w_eco10922, w_eco10923, w_eco10924);
	xor _ECO_out8(cnt[0], sub_wire8, w_eco10925);
	assign w_eco10926 = rst;
	and _ECO_10927(w_eco10927, Tsync[7], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10928(w_eco10928, Tsync[7], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_10929(w_eco10929, Tsync[7], !prev_cnt[0], ena, !prev_state[3], prev_state[1]);
	and _ECO_10930(w_eco10930, Tsync[7], !prev_cnt[0], ena, !prev_state[0]);
	and _ECO_10931(w_eco10931, !Tsync[0], Tsync[7], ena, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1]);
	and _ECO_10932(w_eco10932, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_state[1]);
	and _ECO_10933(w_eco10933, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_state[3], !prev_state[2]);
	and _ECO_10934(w_eco10934, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_state[4], !prev_state[2]);
	and _ECO_10935(w_eco10935, !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_10936(w_eco10936, Tgate[7], prev_cnt[1], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10937(w_eco10937, Tgate[7], prev_cnt[1], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10938(w_eco10938, Tgate[7], !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_10939(w_eco10939, !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_10940(w_eco10940, !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_10941(w_eco10941, !Tsync[0], Tgate[7], prev_cnt[1], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10942(w_eco10942, Tgate[7], prev_cnt[2], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10943(w_eco10943, Tgdel[7], prev_cnt[1], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10944(w_eco10944, Tgate[7], !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_10945(w_eco10945, !Tsync[0], prev_cnt[1], prev_cnt[7], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10946(w_eco10946, Tgate[7], prev_cnt[2], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10947(w_eco10947, Tgdel[7], prev_cnt[1], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10948(w_eco10948, !Tsync[7], prev_cnt[0], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10949(w_eco10949, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], prev_state[1]);
	and _ECO_10950(w_eco10950, Tgate[7], !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_10951(w_eco10951, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_10952(w_eco10952, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10953(w_eco10953, !Tsync[0], !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[0]);
	and _ECO_10954(w_eco10954, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_10955(w_eco10955, !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_10956(w_eco10956, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[1], !prev_cnt[7], !ena);
	and _ECO_10957(w_eco10957, Tsync[0], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10958(w_eco10958, !Tsync[0], Tgate[7], prev_cnt[2], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10959(w_eco10959, Tgate[7], prev_cnt[3], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10960(w_eco10960, Tgdel[7], prev_cnt[2], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10961(w_eco10961, prev_cnt[1], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10962(w_eco10962, !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_10963(w_eco10963, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10964(w_eco10964, !Tsync[0], prev_cnt[2], prev_cnt[7], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10965(w_eco10965, Tgate[7], prev_cnt[3], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10966(w_eco10966, Tgdel[7], prev_cnt[2], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10967(w_eco10967, prev_cnt[1], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10968(w_eco10968, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_10969(w_eco10969, !Tsync[7], prev_cnt[0], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10970(w_eco10970, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], prev_state[1]);
	and _ECO_10971(w_eco10971, Tgate[7], !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_10972(w_eco10972, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_10973(w_eco10973, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10974(w_eco10974, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_10975(w_eco10975, !Tsync[0], !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[0]);
	and _ECO_10976(w_eco10976, Tgate[7], !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_10977(w_eco10977, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_10978(w_eco10978, !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_10979(w_eco10979, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[2], !prev_cnt[7], !ena);
	and _ECO_10980(w_eco10980, Tsync[0], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10981(w_eco10981, Tsync[0], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_10982(w_eco10982, !Tsync[0], Tgate[7], prev_cnt[3], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10983(w_eco10983, Tgate[7], prev_cnt[0], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10984(w_eco10984, Tgdel[7], prev_cnt[3], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10985(w_eco10985, prev_cnt[1], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10986(w_eco10986, prev_cnt[2], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_10987(w_eco10987, !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_10988(w_eco10988, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_10989(w_eco10989, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_10990(w_eco10990, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10991(w_eco10991, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_10992(w_eco10992, !Tsync[0], prev_cnt[3], prev_cnt[7], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_10993(w_eco10993, !Tsync[0], Tgdel[7], prev_cnt[0], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_10994(w_eco10994, !Tsync[0], prev_cnt[0], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_10995(w_eco10995, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_10996(w_eco10996, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_10997(w_eco10997, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_10998(w_eco10998, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], !prev_state[4], !prev_state[2]);
	and _ECO_10999(w_eco10999, !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11000(w_eco11000, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11001(w_eco11001, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11002(w_eco11002, Tgate[7], !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_11003(w_eco11003, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_11004(w_eco11004, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_state[1]);
	and _ECO_11005(w_eco11005, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], !prev_state[3], prev_state[0]);
	and _ECO_11006(w_eco11006, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11007(w_eco11007, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11008(w_eco11008, !Tsync[0], !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[0]);
	and _ECO_11009(w_eco11009, Tgate[7], !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_11010(w_eco11010, !Tsync[7], prev_cnt[6], !prev_cnt[7], !ena);
	and _ECO_11011(w_eco11011, Tsync[0], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11012(w_eco11012, Tsync[0], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11013(w_eco11013, Tsync[0], !Tgate[7], !Tgdel[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11014(w_eco11014, Tgate[7], !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11015(w_eco11015, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11016(w_eco11016, Tgate[7], !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_11017(w_eco11017, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11018(w_eco11018, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11019(w_eco11019, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11020(w_eco11020, !Tsync[0], prev_cnt[0], prev_cnt[7], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_11021(w_eco11021, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11022(w_eco11022, Tgate[7], prev_cnt[0], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11023(w_eco11023, Tgate[7], !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11024(w_eco11024, Tgdel[7], prev_cnt[3], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11025(w_eco11025, prev_cnt[1], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11026(w_eco11026, prev_cnt[2], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11027(w_eco11027, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11028(w_eco11028, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11029(w_eco11029, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_11030(w_eco11030, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_11031(w_eco11031, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11032(w_eco11032, !Tsync[7], prev_cnt[0], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11033(w_eco11033, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11034(w_eco11034, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11035(w_eco11035, Tgdel[7], prev_cnt[0], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11036(w_eco11036, prev_cnt[2], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11037(w_eco11037, prev_cnt[3], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11038(w_eco11038, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], prev_state[1]);
	and _ECO_11039(w_eco11039, Tgate[7], !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_11040(w_eco11040, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_11041(w_eco11041, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_11042(w_eco11042, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11043(w_eco11043, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11044(w_eco11044, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11045(w_eco11045, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_11046(w_eco11046, !Tsync[0], !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[0]);
	and _ECO_11047(w_eco11047, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_11048(w_eco11048, !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11049(w_eco11049, !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_11050(w_eco11050, Tsync[0], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11051(w_eco11051, Tsync[0], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11052(w_eco11052, Tsync[0], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11053(w_eco11053, Tsync[0], !Tgate[7], !Tgdel[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11054(w_eco11054, Tgate[7], !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11055(w_eco11055, Tgdel[7], prev_cnt[4], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11056(w_eco11056, prev_cnt[1], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11057(w_eco11057, prev_cnt[3], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11058(w_eco11058, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11059(w_eco11059, !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11060(w_eco11060, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_11061(w_eco11061, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[3], !prev_cnt[7], !ena);
	and _ECO_11062(w_eco11062, Tgate[7], !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_11063(w_eco11063, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11064(w_eco11064, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11065(w_eco11065, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11066(w_eco11066, Tsync[0], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], prev_state[0]);
	and _ECO_11067(w_eco11067, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11068(w_eco11068, Tgate[7], !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11069(w_eco11069, Tgdel[7], prev_cnt[0], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11070(w_eco11070, prev_cnt[2], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11071(w_eco11071, prev_cnt[3], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11072(w_eco11072, Tgdel[7], prev_cnt[4], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11073(w_eco11073, prev_cnt[1], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11074(w_eco11074, prev_cnt[3], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11075(w_eco11075, prev_cnt[0], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11076(w_eco11076, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11077(w_eco11077, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11078(w_eco11078, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11079(w_eco11079, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], !prev_state[4], !prev_state[2]);
	and _ECO_11080(w_eco11080, !Tsync[7], prev_cnt[0], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11081(w_eco11081, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11082(w_eco11082, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11083(w_eco11083, !Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], prev_state[1]);
	and _ECO_11084(w_eco11084, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_11085(w_eco11085, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_11086(w_eco11086, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], !prev_state[3], prev_state[0]);
	and _ECO_11087(w_eco11087, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11088(w_eco11088, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11089(w_eco11089, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11090(w_eco11090, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11091(w_eco11091, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_11092(w_eco11092, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_11093(w_eco11093, !Tsync[0], !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[0]);
	and _ECO_11094(w_eco11094, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_11095(w_eco11095, !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11096(w_eco11096, !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11097(w_eco11097, !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_11098(w_eco11098, !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_11099(w_eco11099, !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], !ena);
	and _ECO_11100(w_eco11100, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11101(w_eco11101, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11102(w_eco11102, Tgdel[7], prev_cnt[5], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11103(w_eco11103, prev_cnt[6], prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11104(w_eco11104, !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11105(w_eco11105, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], !ena);
	and _ECO_11106(w_eco11106, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_11107(w_eco11107, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[4], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11108(w_eco11108, Tsync[0], !Tsync[7], prev_cnt[6], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11109(w_eco11109, Tgdel[7], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11110(w_eco11110, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11111(w_eco11111, Tgdel[7], prev_cnt[5], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11112(w_eco11112, prev_cnt[6], prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11113(w_eco11113, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[3], !prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11114(w_eco11114, Tsync[0], !Tsync[7], prev_cnt[6], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11115(w_eco11115, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], !prev_state[4], !prev_state[2]);
	and _ECO_11116(w_eco11116, !Tsync[7], prev_cnt[0], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11117(w_eco11117, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11118(w_eco11118, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], prev_state[1]);
	and _ECO_11119(w_eco11119, !prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[3], prev_state[1]);
	and _ECO_11120(w_eco11120, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], !prev_state[3], prev_state[0]);
	and _ECO_11121(w_eco11121, Tsync[0], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11122(w_eco11122, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11123(w_eco11123, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11124(w_eco11124, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11125(w_eco11125, Tgdel[7], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11126(w_eco11126, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11127(w_eco11127, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11128(w_eco11128, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11129(w_eco11129, !Tsync[0], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], ena, prev_state[0]);
	and _ECO_11130(w_eco11130, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_11131(w_eco11131, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11132(w_eco11132, !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11133(w_eco11133, !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11134(w_eco11134, !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_11135(w_eco11135, !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], !ena);
	and _ECO_11136(w_eco11136, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[4], !prev_cnt[7], !ena);
	and _ECO_11137(w_eco11137, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11138(w_eco11138, prev_cnt[1], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11139(w_eco11139, prev_cnt[2], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11140(w_eco11140, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11141(w_eco11141, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11142(w_eco11142, !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11143(w_eco11143, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11144(w_eco11144, !prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, prev_state[1], !prev_state[0]);
	and _ECO_11145(w_eco11145, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], prev_state[1], !prev_state[0]);
	and _ECO_11146(w_eco11146, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11147(w_eco11147, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11148(w_eco11148, Tsync[0], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], prev_state[0]);
	and _ECO_11149(w_eco11149, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11150(w_eco11150, Tgdel[7], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11151(w_eco11151, prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11152(w_eco11152, prev_cnt[1], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11153(w_eco11153, prev_cnt[2], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11154(w_eco11154, prev_cnt[0], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11155(w_eco11155, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11156(w_eco11156, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11157(w_eco11157, !Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], !prev_state[4], !prev_state[2]);
	and _ECO_11158(w_eco11158, !Tsync[7], prev_cnt[0], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11159(w_eco11159, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11160(w_eco11160, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11161(w_eco11161, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11162(w_eco11162, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], prev_state[1]);
	and _ECO_11163(w_eco11163, Tgate[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_11164(w_eco11164, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11165(w_eco11165, !Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], !prev_state[3], prev_state[0]);
	and _ECO_11166(w_eco11166, Tsync[0], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11167(w_eco11167, Tsync[0], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11168(w_eco11168, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11169(w_eco11169, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11170(w_eco11170, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11171(w_eco11171, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11172(w_eco11172, Tgdel[7], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11173(w_eco11173, prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11174(w_eco11174, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11175(w_eco11175, !prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11176(w_eco11176, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11177(w_eco11177, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11178(w_eco11178, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11179(w_eco11179, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11180(w_eco11180, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_11181(w_eco11181, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_11182(w_eco11182, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], prev_state[3], prev_state[0]);
	and _ECO_11183(w_eco11183, !Tsync[0], !prev_cnt[0], prev_cnt[6], prev_cnt[7], ena, prev_state[0]);
	and _ECO_11184(w_eco11184, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11185(w_eco11185, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11186(w_eco11186, !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11187(w_eco11187, !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11188(w_eco11188, !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11189(w_eco11189, !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[5], !prev_cnt[7], !ena);
	and _ECO_11190(w_eco11190, !Tgate[7], !Tgdel[7], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], !ena);
	and _ECO_11191(w_eco11191, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11192(w_eco11192, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11193(w_eco11193, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11194(w_eco11194, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11195(w_eco11195, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11196(w_eco11196, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11197(w_eco11197, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11198(w_eco11198, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11199(w_eco11199, Tgate[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11200(w_eco11200, prev_cnt[1], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11201(w_eco11201, prev_cnt[2], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11202(w_eco11202, prev_cnt[3], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11203(w_eco11203, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11204(w_eco11204, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11205(w_eco11205, !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11206(w_eco11206, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11207(w_eco11207, Tgate[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11208(w_eco11208, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11209(w_eco11209, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11210(w_eco11210, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11211(w_eco11211, !Tsync[0], Tgate[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_11212(w_eco11212, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_state[0]);
	and _ECO_11213(w_eco11213, Tgdel[7], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11214(w_eco11214, Tgdel[7], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11215(w_eco11215, prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11216(w_eco11216, Tgate[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11217(w_eco11217, prev_cnt[1], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11218(w_eco11218, prev_cnt[2], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11219(w_eco11219, prev_cnt[3], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11220(w_eco11220, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11221(w_eco11221, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11222(w_eco11222, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11223(w_eco11223, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11224(w_eco11224, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], !prev_state[4], !prev_state[2]);
	and _ECO_11225(w_eco11225, !Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11226(w_eco11226, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11227(w_eco11227, prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11228(w_eco11228, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11229(w_eco11229, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11230(w_eco11230, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11231(w_eco11231, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11232(w_eco11232, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], prev_state[1]);
	and _ECO_11233(w_eco11233, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_11234(w_eco11234, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11235(w_eco11235, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11236(w_eco11236, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11237(w_eco11237, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], !prev_state[3], prev_state[0]);
	and _ECO_11238(w_eco11238, !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_11239(w_eco11239, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11240(w_eco11240, Tsync[0], !Tsync[7], prev_cnt[6], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11241(w_eco11241, Tgdel[7], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11242(w_eco11242, Tgdel[7], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11243(w_eco11243, prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11244(w_eco11244, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11245(w_eco11245, Tgate[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11246(w_eco11246, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11247(w_eco11247, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11248(w_eco11248, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11249(w_eco11249, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11250(w_eco11250, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11251(w_eco11251, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11252(w_eco11252, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11253(w_eco11253, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_11254(w_eco11254, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_11255(w_eco11255, !Tsync[0], Tgate[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_11256(w_eco11256, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11257(w_eco11257, !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11258(w_eco11258, !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11259(w_eco11259, !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11260(w_eco11260, !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], !ena);
	and _ECO_11261(w_eco11261, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11262(w_eco11262, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11263(w_eco11263, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11264(w_eco11264, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11265(w_eco11265, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11266(w_eco11266, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11267(w_eco11267, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11268(w_eco11268, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11269(w_eco11269, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11270(w_eco11270, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11271(w_eco11271, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11272(w_eco11272, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11273(w_eco11273, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11274(w_eco11274, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11275(w_eco11275, !prev_cnt[14], prev_cnt[1], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11276(w_eco11276, prev_cnt[2], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11277(w_eco11277, prev_cnt[3], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11278(w_eco11278, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11279(w_eco11279, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11280(w_eco11280, !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11281(w_eco11281, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11282(w_eco11282, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11283(w_eco11283, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11284(w_eco11284, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11285(w_eco11285, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11286(w_eco11286, Tsync[0], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], prev_state[0]);
	and _ECO_11287(w_eco11287, !Tsync[0], Tgdel[7], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_11288(w_eco11288, Tgdel[7], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11289(w_eco11289, Tgdel[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11290(w_eco11290, prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11291(w_eco11291, prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11292(w_eco11292, !prev_cnt[14], prev_cnt[1], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11293(w_eco11293, prev_cnt[2], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11294(w_eco11294, prev_cnt[3], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11295(w_eco11295, prev_cnt[0], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11296(w_eco11296, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11297(w_eco11297, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11298(w_eco11298, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11299(w_eco11299, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11300(w_eco11300, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], !prev_state[4], !prev_state[2]);
	and _ECO_11301(w_eco11301, !Tsync[7], !prev_cnt[14], prev_cnt[0], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11302(w_eco11302, Tgdel[7], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11303(w_eco11303, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11304(w_eco11304, prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11305(w_eco11305, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11306(w_eco11306, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11307(w_eco11307, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11308(w_eco11308, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11309(w_eco11309, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11310(w_eco11310, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11311(w_eco11311, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11312(w_eco11312, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11313(w_eco11313, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], prev_state[1]);
	and _ECO_11314(w_eco11314, Tgate[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_11315(w_eco11315, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11316(w_eco11316, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11317(w_eco11317, !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], !prev_state[3], prev_state[0]);
	and _ECO_11318(w_eco11318, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11319(w_eco11319, !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11320(w_eco11320, !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_11321(w_eco11321, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11322(w_eco11322, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11323(w_eco11323, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11324(w_eco11324, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11325(w_eco11325, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11326(w_eco11326, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11327(w_eco11327, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11328(w_eco11328, Tgdel[7], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11329(w_eco11329, Tgdel[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11330(w_eco11330, prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11331(w_eco11331, prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11332(w_eco11332, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0]);
	and _ECO_11333(w_eco11333, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11334(w_eco11334, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11335(w_eco11335, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11336(w_eco11336, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11337(w_eco11337, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11338(w_eco11338, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11339(w_eco11339, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11340(w_eco11340, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11341(w_eco11341, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11342(w_eco11342, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11343(w_eco11343, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_state[3], prev_state[0]);
	and _ECO_11344(w_eco11344, !Tsync[0], Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_11345(w_eco11345, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11346(w_eco11346, !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11347(w_eco11347, !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11348(w_eco11348, !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], !ena);
	and _ECO_11349(w_eco11349, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11350(w_eco11350, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11351(w_eco11351, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11352(w_eco11352, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11353(w_eco11353, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11354(w_eco11354, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11355(w_eco11355, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11356(w_eco11356, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11357(w_eco11357, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11358(w_eco11358, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11359(w_eco11359, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11360(w_eco11360, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11361(w_eco11361, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11362(w_eco11362, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11363(w_eco11363, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11364(w_eco11364, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11365(w_eco11365, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11366(w_eco11366, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11367(w_eco11367, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11368(w_eco11368, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11369(w_eco11369, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11370(w_eco11370, Tgate[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11371(w_eco11371, !prev_cnt[14], prev_cnt[1], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11372(w_eco11372, !prev_cnt[14], prev_cnt[2], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11373(w_eco11373, prev_cnt[3], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11374(w_eco11374, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11375(w_eco11375, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11376(w_eco11376, !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11377(w_eco11377, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11378(w_eco11378, Tgate[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11379(w_eco11379, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11380(w_eco11380, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11381(w_eco11381, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11382(w_eco11382, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11383(w_eco11383, Tsync[0], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], prev_state[0]);
	and _ECO_11384(w_eco11384, !Tsync[0], Tgate[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_11385(w_eco11385, Tgdel[7], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11386(w_eco11386, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11387(w_eco11387, prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11388(w_eco11388, prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11389(w_eco11389, !Tsync[0], Tgate[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_11390(w_eco11390, Tgate[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11391(w_eco11391, !prev_cnt[14], prev_cnt[1], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11392(w_eco11392, !prev_cnt[14], prev_cnt[2], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11393(w_eco11393, prev_cnt[3], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11394(w_eco11394, prev_cnt[0], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11395(w_eco11395, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11396(w_eco11396, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11397(w_eco11397, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11398(w_eco11398, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11399(w_eco11399, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_11400(w_eco11400, Tgdel[7], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11401(w_eco11401, !prev_cnt[0], prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11402(w_eco11402, prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11403(w_eco11403, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11404(w_eco11404, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11405(w_eco11405, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11406(w_eco11406, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11407(w_eco11407, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11408(w_eco11408, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11409(w_eco11409, Tgdel[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_11410(w_eco11410, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11411(w_eco11411, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_11412(w_eco11412, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11413(w_eco11413, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11414(w_eco11414, !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11415(w_eco11415, !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_11416(w_eco11416, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11417(w_eco11417, Tsync[0], !Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11418(w_eco11418, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11419(w_eco11419, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11420(w_eco11420, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11421(w_eco11421, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11422(w_eco11422, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11423(w_eco11423, Tgdel[7], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11424(w_eco11424, prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11425(w_eco11425, prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11426(w_eco11426, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[0]);
	and _ECO_11427(w_eco11427, Tgate[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11428(w_eco11428, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11429(w_eco11429, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11430(w_eco11430, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11431(w_eco11431, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11432(w_eco11432, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11433(w_eco11433, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11434(w_eco11434, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11435(w_eco11435, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11436(w_eco11436, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11437(w_eco11437, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11438(w_eco11438, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11439(w_eco11439, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11440(w_eco11440, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_11441(w_eco11441, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11442(w_eco11442, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11443(w_eco11443, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11444(w_eco11444, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], prev_state[3], prev_state[0]);
	and _ECO_11445(w_eco11445, !Tsync[0], Tgate[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_11446(w_eco11446, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11447(w_eco11447, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11448(w_eco11448, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11449(w_eco11449, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11450(w_eco11450, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11451(w_eco11451, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11452(w_eco11452, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_11453(w_eco11453, !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11454(w_eco11454, !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11455(w_eco11455, !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], !ena);
	and _ECO_11456(w_eco11456, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11457(w_eco11457, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11458(w_eco11458, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11459(w_eco11459, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11460(w_eco11460, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11461(w_eco11461, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11462(w_eco11462, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11463(w_eco11463, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11464(w_eco11464, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11465(w_eco11465, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11466(w_eco11466, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11467(w_eco11467, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11468(w_eco11468, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11469(w_eco11469, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11470(w_eco11470, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11471(w_eco11471, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11472(w_eco11472, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11473(w_eco11473, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11474(w_eco11474, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11475(w_eco11475, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11476(w_eco11476, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11477(w_eco11477, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11478(w_eco11478, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11479(w_eco11479, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11480(w_eco11480, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11481(w_eco11481, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11482(w_eco11482, !prev_cnt[14], prev_cnt[2], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11483(w_eco11483, !prev_cnt[14], prev_cnt[3], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11484(w_eco11484, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11485(w_eco11485, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11486(w_eco11486, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11487(w_eco11487, !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11488(w_eco11488, Tgdel[7], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11489(w_eco11489, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11490(w_eco11490, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11491(w_eco11491, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11492(w_eco11492, Tsync[0], !Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], prev_state[0]);
	and _ECO_11493(w_eco11493, !Tsync[0], Tgdel[7], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_11494(w_eco11494, !Tsync[0], Tgdel[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_11495(w_eco11495, Tgdel[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[1], !prev_state[0]);
	and _ECO_11496(w_eco11496, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11497(w_eco11497, prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11498(w_eco11498, prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11499(w_eco11499, !Tsync[0], Tgate[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_11500(w_eco11500, !Tsync[0], Tgdel[7], prev_cnt[14], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_11501(w_eco11501, Tgdel[7], !prev_cnt[0], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11502(w_eco11502, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11503(w_eco11503, Tgdel[7], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11504(w_eco11504, !prev_cnt[0], prev_cnt[2], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11505(w_eco11505, Tgdel[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_11506(w_eco11506, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11507(w_eco11507, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11508(w_eco11508, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11509(w_eco11509, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11510(w_eco11510, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11511(w_eco11511, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11512(w_eco11512, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11513(w_eco11513, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11514(w_eco11514, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11515(w_eco11515, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11516(w_eco11516, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11517(w_eco11517, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11518(w_eco11518, !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_11519(w_eco11519, !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11520(w_eco11520, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_11521(w_eco11521, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11522(w_eco11522, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11523(w_eco11523, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11524(w_eco11524, Tsync[0], !Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11525(w_eco11525, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11526(w_eco11526, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11527(w_eco11527, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11528(w_eco11528, Tsync[0], !Tgate[7], !Tgdel[7], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11529(w_eco11529, Tgdel[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11530(w_eco11530, prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11531(w_eco11531, prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_11532(w_eco11532, Tgdel[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_11533(w_eco11533, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11534(w_eco11534, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11535(w_eco11535, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11536(w_eco11536, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11537(w_eco11537, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11538(w_eco11538, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11539(w_eco11539, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11540(w_eco11540, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11541(w_eco11541, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11542(w_eco11542, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11543(w_eco11543, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11544(w_eco11544, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11545(w_eco11545, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11546(w_eco11546, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11547(w_eco11547, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], prev_state[3], prev_state[0]);
	and _ECO_11548(w_eco11548, !Tsync[0], Tgdel[7], !prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_11549(w_eco11549, !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11550(w_eco11550, !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11551(w_eco11551, !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], !ena);
	and _ECO_11552(w_eco11552, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11553(w_eco11553, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11554(w_eco11554, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11555(w_eco11555, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11556(w_eco11556, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11557(w_eco11557, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11558(w_eco11558, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11559(w_eco11559, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11560(w_eco11560, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11561(w_eco11561, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11562(w_eco11562, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11563(w_eco11563, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11564(w_eco11564, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11565(w_eco11565, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11566(w_eco11566, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11567(w_eco11567, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11568(w_eco11568, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11569(w_eco11569, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11570(w_eco11570, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11571(w_eco11571, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11572(w_eco11572, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11573(w_eco11573, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11574(w_eco11574, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11575(w_eco11575, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11576(w_eco11576, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11577(w_eco11577, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11578(w_eco11578, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11579(w_eco11579, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11580(w_eco11580, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11581(w_eco11581, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11582(w_eco11582, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11583(w_eco11583, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11584(w_eco11584, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11585(w_eco11585, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11586(w_eco11586, Tgdel[7], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11587(w_eco11587, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11588(w_eco11588, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11589(w_eco11589, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], prev_state[0]);
	and _ECO_11590(w_eco11590, !Tsync[0], Tgdel[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1]);
	and _ECO_11591(w_eco11591, Tgdel[7], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11592(w_eco11592, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11593(w_eco11593, !prev_cnt[14], prev_cnt[2], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11594(w_eco11594, !prev_cnt[14], prev_cnt[3], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11595(w_eco11595, prev_cnt[0], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11596(w_eco11596, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11597(w_eco11597, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11598(w_eco11598, !prev_cnt[14], prev_cnt[3], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11599(w_eco11599, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11600(w_eco11600, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11601(w_eco11601, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11602(w_eco11602, prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11603(w_eco11603, prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11604(w_eco11604, !Tsync[0], Tgdel[7], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_11605(w_eco11605, Tgdel[7], !prev_cnt[0], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11606(w_eco11606, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11607(w_eco11607, !prev_cnt[0], prev_cnt[3], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11608(w_eco11608, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11609(w_eco11609, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11610(w_eco11610, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11611(w_eco11611, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11612(w_eco11612, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11613(w_eco11613, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11614(w_eco11614, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11615(w_eco11615, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11616(w_eco11616, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11617(w_eco11617, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11618(w_eco11618, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11619(w_eco11619, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11620(w_eco11620, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11621(w_eco11621, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11622(w_eco11622, !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_11623(w_eco11623, !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_11624(w_eco11624, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11625(w_eco11625, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_11626(w_eco11626, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11627(w_eco11627, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11628(w_eco11628, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11629(w_eco11629, Tsync[0], !Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11630(w_eco11630, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11631(w_eco11631, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11632(w_eco11632, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11633(w_eco11633, prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11634(w_eco11634, prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_11635(w_eco11635, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11636(w_eco11636, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11637(w_eco11637, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11638(w_eco11638, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11639(w_eco11639, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11640(w_eco11640, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11641(w_eco11641, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11642(w_eco11642, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11643(w_eco11643, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11644(w_eco11644, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11645(w_eco11645, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11646(w_eco11646, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11647(w_eco11647, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11648(w_eco11648, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11649(w_eco11649, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11650(w_eco11650, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11651(w_eco11651, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11652(w_eco11652, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], prev_state[3], prev_state[0]);
	and _ECO_11653(w_eco11653, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11654(w_eco11654, !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11655(w_eco11655, !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], !ena);
	and _ECO_11656(w_eco11656, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11657(w_eco11657, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11658(w_eco11658, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11659(w_eco11659, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11660(w_eco11660, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11661(w_eco11661, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11662(w_eco11662, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11663(w_eco11663, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11664(w_eco11664, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11665(w_eco11665, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11666(w_eco11666, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11667(w_eco11667, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11668(w_eco11668, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11669(w_eco11669, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11670(w_eco11670, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11671(w_eco11671, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11672(w_eco11672, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11673(w_eco11673, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11674(w_eco11674, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11675(w_eco11675, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11676(w_eco11676, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11677(w_eco11677, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11678(w_eco11678, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11679(w_eco11679, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11680(w_eco11680, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11681(w_eco11681, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11682(w_eco11682, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11683(w_eco11683, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11684(w_eco11684, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11685(w_eco11685, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11686(w_eco11686, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11687(w_eco11687, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11688(w_eco11688, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11689(w_eco11689, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11690(w_eco11690, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11691(w_eco11691, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11692(w_eco11692, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11693(w_eco11693, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11694(w_eco11694, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11695(w_eco11695, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11696(w_eco11696, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11697(w_eco11697, Tgdel[7], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11698(w_eco11698, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11699(w_eco11699, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_11700(w_eco11700, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], prev_state[0]);
	and _ECO_11701(w_eco11701, Tgdel[7], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11702(w_eco11702, !prev_cnt[0], prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11703(w_eco11703, !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_11704(w_eco11704, !prev_cnt[14], prev_cnt[3], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11705(w_eco11705, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11706(w_eco11706, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11707(w_eco11707, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11708(w_eco11708, Tgdel[7], !prev_cnt[0], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11709(w_eco11709, Tgdel[7], prev_cnt[14], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11710(w_eco11710, Tgdel[7], prev_cnt[14], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11711(w_eco11711, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11712(w_eco11712, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11713(w_eco11713, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], prev_state[3], prev_state[0]);
	and _ECO_11714(w_eco11714, !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_11715(w_eco11715, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11716(w_eco11716, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11717(w_eco11717, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11718(w_eco11718, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11719(w_eco11719, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11720(w_eco11720, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11721(w_eco11721, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11722(w_eco11722, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11723(w_eco11723, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11724(w_eco11724, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11725(w_eco11725, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11726(w_eco11726, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11727(w_eco11727, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11728(w_eco11728, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11729(w_eco11729, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11730(w_eco11730, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11731(w_eco11731, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11732(w_eco11732, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11733(w_eco11733, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11734(w_eco11734, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11735(w_eco11735, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11736(w_eco11736, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11737(w_eco11737, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11738(w_eco11738, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11739(w_eco11739, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11740(w_eco11740, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11741(w_eco11741, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11742(w_eco11742, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11743(w_eco11743, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11744(w_eco11744, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11745(w_eco11745, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11746(w_eco11746, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11747(w_eco11747, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11748(w_eco11748, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11749(w_eco11749, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11750(w_eco11750, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11751(w_eco11751, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11752(w_eco11752, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11753(w_eco11753, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11754(w_eco11754, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11755(w_eco11755, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11756(w_eco11756, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11757(w_eco11757, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11758(w_eco11758, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11759(w_eco11759, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11760(w_eco11760, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11761(w_eco11761, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11762(w_eco11762, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11763(w_eco11763, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11764(w_eco11764, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11765(w_eco11765, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11766(w_eco11766, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11767(w_eco11767, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11768(w_eco11768, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11769(w_eco11769, Tgdel[7], !prev_cnt[0], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11770(w_eco11770, Tgdel[7], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[1], !prev_state[0]);
	and _ECO_11771(w_eco11771, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11772(w_eco11772, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11773(w_eco11773, !prev_cnt[0], prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11774(w_eco11774, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11775(w_eco11775, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11776(w_eco11776, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11777(w_eco11777, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11778(w_eco11778, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11779(w_eco11779, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11780(w_eco11780, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11781(w_eco11781, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11782(w_eco11782, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11783(w_eco11783, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11784(w_eco11784, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11785(w_eco11785, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11786(w_eco11786, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11787(w_eco11787, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11788(w_eco11788, !prev_cnt[14], prev_cnt[0], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_11789(w_eco11789, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11790(w_eco11790, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11791(w_eco11791, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11792(w_eco11792, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11793(w_eco11793, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11794(w_eco11794, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11795(w_eco11795, !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_11796(w_eco11796, !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_11797(w_eco11797, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_11798(w_eco11798, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11799(w_eco11799, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11800(w_eco11800, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11801(w_eco11801, Tsync[0], !Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11802(w_eco11802, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11803(w_eco11803, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11804(w_eco11804, !prev_cnt[0], prev_cnt[4], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_11805(w_eco11805, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11806(w_eco11806, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11807(w_eco11807, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11808(w_eco11808, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11809(w_eco11809, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11810(w_eco11810, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11811(w_eco11811, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11812(w_eco11812, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11813(w_eco11813, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11814(w_eco11814, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11815(w_eco11815, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11816(w_eco11816, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11817(w_eco11817, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11818(w_eco11818, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11819(w_eco11819, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11820(w_eco11820, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11821(w_eco11821, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11822(w_eco11822, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], prev_state[3], prev_state[0]);
	and _ECO_11823(w_eco11823, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11824(w_eco11824, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11825(w_eco11825, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11826(w_eco11826, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11827(w_eco11827, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11828(w_eco11828, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11829(w_eco11829, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11830(w_eco11830, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11831(w_eco11831, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11832(w_eco11832, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11833(w_eco11833, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11834(w_eco11834, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11835(w_eco11835, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11836(w_eco11836, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11837(w_eco11837, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11838(w_eco11838, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11839(w_eco11839, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11840(w_eco11840, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11841(w_eco11841, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11842(w_eco11842, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11843(w_eco11843, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11844(w_eco11844, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11845(w_eco11845, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11846(w_eco11846, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11847(w_eco11847, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11848(w_eco11848, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11849(w_eco11849, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11850(w_eco11850, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11851(w_eco11851, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11852(w_eco11852, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11853(w_eco11853, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11854(w_eco11854, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11855(w_eco11855, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11856(w_eco11856, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11857(w_eco11857, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11858(w_eco11858, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11859(w_eco11859, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11860(w_eco11860, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11861(w_eco11861, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11862(w_eco11862, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11863(w_eco11863, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11864(w_eco11864, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11865(w_eco11865, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11866(w_eco11866, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11867(w_eco11867, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11868(w_eco11868, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11869(w_eco11869, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11870(w_eco11870, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11871(w_eco11871, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11872(w_eco11872, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11873(w_eco11873, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11874(w_eco11874, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11875(w_eco11875, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11876(w_eco11876, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11877(w_eco11877, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11878(w_eco11878, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11879(w_eco11879, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11880(w_eco11880, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11881(w_eco11881, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11882(w_eco11882, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11883(w_eco11883, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11884(w_eco11884, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11885(w_eco11885, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11886(w_eco11886, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11887(w_eco11887, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_11888(w_eco11888, Tgdel[7], !prev_cnt[0], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11889(w_eco11889, Tgdel[7], !prev_cnt[0], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_11890(w_eco11890, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11891(w_eco11891, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11892(w_eco11892, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11893(w_eco11893, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11894(w_eco11894, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11895(w_eco11895, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11896(w_eco11896, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11897(w_eco11897, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11898(w_eco11898, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11899(w_eco11899, !Tsync[0], Tsync[7], !prev_cnt[0], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11900(w_eco11900, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11901(w_eco11901, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11902(w_eco11902, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11903(w_eco11903, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11904(w_eco11904, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11905(w_eco11905, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11906(w_eco11906, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_11907(w_eco11907, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11908(w_eco11908, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11909(w_eco11909, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_11910(w_eco11910, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11911(w_eco11911, !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_11912(w_eco11912, !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_11913(w_eco11913, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_11914(w_eco11914, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11915(w_eco11915, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11916(w_eco11916, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11917(w_eco11917, Tsync[0], !Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11918(w_eco11918, Tsync[0], !Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_11919(w_eco11919, !prev_cnt[0], prev_cnt[5], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_11920(w_eco11920, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11921(w_eco11921, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11922(w_eco11922, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11923(w_eco11923, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11924(w_eco11924, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11925(w_eco11925, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11926(w_eco11926, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11927(w_eco11927, prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11928(w_eco11928, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11929(w_eco11929, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11930(w_eco11930, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11931(w_eco11931, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11932(w_eco11932, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11933(w_eco11933, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11934(w_eco11934, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_11935(w_eco11935, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11936(w_eco11936, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_11937(w_eco11937, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11938(w_eco11938, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11939(w_eco11939, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[0]);
	and _ECO_11940(w_eco11940, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11941(w_eco11941, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11942(w_eco11942, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11943(w_eco11943, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11944(w_eco11944, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11945(w_eco11945, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11946(w_eco11946, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11947(w_eco11947, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11948(w_eco11948, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11949(w_eco11949, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11950(w_eco11950, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11951(w_eco11951, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11952(w_eco11952, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11953(w_eco11953, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11954(w_eco11954, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11955(w_eco11955, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11956(w_eco11956, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11957(w_eco11957, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11958(w_eco11958, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11959(w_eco11959, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11960(w_eco11960, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11961(w_eco11961, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11962(w_eco11962, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11963(w_eco11963, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_11964(w_eco11964, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11965(w_eco11965, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11966(w_eco11966, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11967(w_eco11967, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11968(w_eco11968, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11969(w_eco11969, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11970(w_eco11970, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11971(w_eco11971, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11972(w_eco11972, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11973(w_eco11973, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11974(w_eco11974, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11975(w_eco11975, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11976(w_eco11976, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11977(w_eco11977, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11978(w_eco11978, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11979(w_eco11979, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11980(w_eco11980, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11981(w_eco11981, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11982(w_eco11982, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11983(w_eco11983, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11984(w_eco11984, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11985(w_eco11985, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11986(w_eco11986, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11987(w_eco11987, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11988(w_eco11988, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11989(w_eco11989, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11990(w_eco11990, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_11991(w_eco11991, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11992(w_eco11992, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11993(w_eco11993, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_11994(w_eco11994, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11995(w_eco11995, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11996(w_eco11996, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11997(w_eco11997, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11998(w_eco11998, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_11999(w_eco11999, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12000(w_eco12000, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12001(w_eco12001, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12002(w_eco12002, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12003(w_eco12003, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12004(w_eco12004, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12005(w_eco12005, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12006(w_eco12006, !Tsync[0], Tsync[7], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12007(w_eco12007, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12008(w_eco12008, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12009(w_eco12009, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12010(w_eco12010, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12011(w_eco12011, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12012(w_eco12012, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12013(w_eco12013, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12014(w_eco12014, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12015(w_eco12015, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12016(w_eco12016, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12017(w_eco12017, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12018(w_eco12018, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12019(w_eco12019, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12020(w_eco12020, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12021(w_eco12021, !Tsync[0], Tsync[7], !prev_cnt[0], ena, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12022(w_eco12022, !Tsync[0], Tsync[7], !prev_cnt[0], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12023(w_eco12023, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_12024(w_eco12024, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12025(w_eco12025, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12026(w_eco12026, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12027(w_eco12027, !prev_cnt[14], !prev_cnt[0], prev_cnt[1], prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_12028(w_eco12028, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12029(w_eco12029, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12030(w_eco12030, !prev_cnt[14], !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_12031(w_eco12031, !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_12032(w_eco12032, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_12033(w_eco12033, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[9], ena, prev_state[1], !prev_state[0]);
	and _ECO_12034(w_eco12034, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12035(w_eco12035, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12036(w_eco12036, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12037(w_eco12037, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12038(w_eco12038, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12039(w_eco12039, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12040(w_eco12040, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12041(w_eco12041, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12042(w_eco12042, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12043(w_eco12043, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12044(w_eco12044, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12045(w_eco12045, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12046(w_eco12046, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12047(w_eco12047, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12048(w_eco12048, prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12049(w_eco12049, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12050(w_eco12050, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12051(w_eco12051, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12052(w_eco12052, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12053(w_eco12053, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12054(w_eco12054, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12055(w_eco12055, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12056(w_eco12056, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12057(w_eco12057, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12058(w_eco12058, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12059(w_eco12059, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12060(w_eco12060, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12061(w_eco12061, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12062(w_eco12062, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12063(w_eco12063, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12064(w_eco12064, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12065(w_eco12065, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12066(w_eco12066, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12067(w_eco12067, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12068(w_eco12068, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12069(w_eco12069, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12070(w_eco12070, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12071(w_eco12071, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12072(w_eco12072, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12073(w_eco12073, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12074(w_eco12074, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12075(w_eco12075, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12076(w_eco12076, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12077(w_eco12077, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12078(w_eco12078, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12079(w_eco12079, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12080(w_eco12080, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12081(w_eco12081, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12082(w_eco12082, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12083(w_eco12083, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12084(w_eco12084, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12085(w_eco12085, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12086(w_eco12086, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12087(w_eco12087, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12088(w_eco12088, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12089(w_eco12089, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12090(w_eco12090, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12091(w_eco12091, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12092(w_eco12092, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12093(w_eco12093, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12094(w_eco12094, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12095(w_eco12095, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12096(w_eco12096, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12097(w_eco12097, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12098(w_eco12098, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[1], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12099(w_eco12099, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12100(w_eco12100, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12101(w_eco12101, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12102(w_eco12102, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12103(w_eco12103, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12104(w_eco12104, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12105(w_eco12105, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12106(w_eco12106, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12107(w_eco12107, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12108(w_eco12108, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12109(w_eco12109, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12110(w_eco12110, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12111(w_eco12111, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12112(w_eco12112, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12113(w_eco12113, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12114(w_eco12114, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12115(w_eco12115, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12116(w_eco12116, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12117(w_eco12117, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12118(w_eco12118, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12119(w_eco12119, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12120(w_eco12120, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12121(w_eco12121, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12122(w_eco12122, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12123(w_eco12123, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12124(w_eco12124, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12125(w_eco12125, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12126(w_eco12126, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12127(w_eco12127, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12128(w_eco12128, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12129(w_eco12129, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12130(w_eco12130, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12131(w_eco12131, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12132(w_eco12132, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12133(w_eco12133, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12134(w_eco12134, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12135(w_eco12135, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12136(w_eco12136, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12137(w_eco12137, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12138(w_eco12138, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12139(w_eco12139, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12140(w_eco12140, !Tsync[0], Tsync[7], !prev_cnt[0], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12141(w_eco12141, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12142(w_eco12142, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12143(w_eco12143, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12144(w_eco12144, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12145(w_eco12145, !prev_cnt[14], !prev_cnt[0], prev_cnt[2], prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_12146(w_eco12146, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12147(w_eco12147, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12148(w_eco12148, !prev_cnt[14], !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_12149(w_eco12149, !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_12150(w_eco12150, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[8], ena, prev_state[1], !prev_state[0]);
	and _ECO_12151(w_eco12151, Tsync[0], !Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12152(w_eco12152, Tsync[0], !Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12153(w_eco12153, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12154(w_eco12154, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12155(w_eco12155, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12156(w_eco12156, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12157(w_eco12157, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12158(w_eco12158, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12159(w_eco12159, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12160(w_eco12160, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12161(w_eco12161, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12162(w_eco12162, !Tgate[7], !Tgdel[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12163(w_eco12163, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12164(w_eco12164, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12165(w_eco12165, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12166(w_eco12166, Tsync[7], !prev_cnt[0], ena, !prev_state[4], !prev_state[3], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12167(w_eco12167, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12168(w_eco12168, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12169(w_eco12169, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12170(w_eco12170, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12171(w_eco12171, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12172(w_eco12172, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12173(w_eco12173, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12174(w_eco12174, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12175(w_eco12175, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12176(w_eco12176, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12177(w_eco12177, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12178(w_eco12178, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12179(w_eco12179, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12180(w_eco12180, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12181(w_eco12181, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12182(w_eco12182, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12183(w_eco12183, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12184(w_eco12184, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12185(w_eco12185, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12186(w_eco12186, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12187(w_eco12187, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12188(w_eco12188, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12189(w_eco12189, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12190(w_eco12190, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12191(w_eco12191, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12192(w_eco12192, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12193(w_eco12193, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12194(w_eco12194, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12195(w_eco12195, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12196(w_eco12196, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12197(w_eco12197, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12198(w_eco12198, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12199(w_eco12199, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12200(w_eco12200, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12201(w_eco12201, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12202(w_eco12202, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12203(w_eco12203, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12204(w_eco12204, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12205(w_eco12205, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12206(w_eco12206, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12207(w_eco12207, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12208(w_eco12208, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12209(w_eco12209, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12210(w_eco12210, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12211(w_eco12211, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12212(w_eco12212, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12213(w_eco12213, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12214(w_eco12214, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12215(w_eco12215, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12216(w_eco12216, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12217(w_eco12217, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12218(w_eco12218, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12219(w_eco12219, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12220(w_eco12220, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12221(w_eco12221, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[2], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12222(w_eco12222, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12223(w_eco12223, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12224(w_eco12224, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12225(w_eco12225, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12226(w_eco12226, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12227(w_eco12227, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12228(w_eco12228, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12229(w_eco12229, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12230(w_eco12230, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12231(w_eco12231, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12232(w_eco12232, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12233(w_eco12233, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12234(w_eco12234, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12235(w_eco12235, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12236(w_eco12236, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12237(w_eco12237, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12238(w_eco12238, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12239(w_eco12239, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12240(w_eco12240, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12241(w_eco12241, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12242(w_eco12242, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12243(w_eco12243, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12244(w_eco12244, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12245(w_eco12245, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12246(w_eco12246, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12247(w_eco12247, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12248(w_eco12248, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12249(w_eco12249, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12250(w_eco12250, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12251(w_eco12251, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12252(w_eco12252, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12253(w_eco12253, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12254(w_eco12254, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12255(w_eco12255, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12256(w_eco12256, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12257(w_eco12257, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12258(w_eco12258, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12259(w_eco12259, !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12260(w_eco12260, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12261(w_eco12261, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12262(w_eco12262, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12263(w_eco12263, !Tsync[0], Tsync[7], !prev_cnt[0], ena, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12264(w_eco12264, !prev_cnt[14], !prev_cnt[0], prev_cnt[3], prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_12265(w_eco12265, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12266(w_eco12266, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12267(w_eco12267, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12268(w_eco12268, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12269(w_eco12269, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12270(w_eco12270, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12271(w_eco12271, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_12272(w_eco12272, !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[10], ena, prev_state[1], !prev_state[0]);
	and _ECO_12273(w_eco12273, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12274(w_eco12274, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12275(w_eco12275, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12276(w_eco12276, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12277(w_eco12277, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12278(w_eco12278, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12279(w_eco12279, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12280(w_eco12280, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12281(w_eco12281, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12282(w_eco12282, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12283(w_eco12283, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12284(w_eco12284, prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12285(w_eco12285, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12286(w_eco12286, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12287(w_eco12287, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12288(w_eco12288, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12289(w_eco12289, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12290(w_eco12290, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12291(w_eco12291, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12292(w_eco12292, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12293(w_eco12293, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12294(w_eco12294, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12295(w_eco12295, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12296(w_eco12296, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12297(w_eco12297, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12298(w_eco12298, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12299(w_eco12299, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12300(w_eco12300, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12301(w_eco12301, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12302(w_eco12302, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12303(w_eco12303, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12304(w_eco12304, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12305(w_eco12305, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12306(w_eco12306, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12307(w_eco12307, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12308(w_eco12308, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12309(w_eco12309, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12310(w_eco12310, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12311(w_eco12311, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12312(w_eco12312, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12313(w_eco12313, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12314(w_eco12314, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12315(w_eco12315, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12316(w_eco12316, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12317(w_eco12317, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12318(w_eco12318, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12319(w_eco12319, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12320(w_eco12320, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12321(w_eco12321, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12322(w_eco12322, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12323(w_eco12323, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12324(w_eco12324, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12325(w_eco12325, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12326(w_eco12326, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12327(w_eco12327, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12328(w_eco12328, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12329(w_eco12329, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12330(w_eco12330, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12331(w_eco12331, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12332(w_eco12332, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12333(w_eco12333, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12334(w_eco12334, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12335(w_eco12335, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12336(w_eco12336, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12337(w_eco12337, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12338(w_eco12338, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12339(w_eco12339, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12340(w_eco12340, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12341(w_eco12341, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12342(w_eco12342, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12343(w_eco12343, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12344(w_eco12344, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12345(w_eco12345, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12346(w_eco12346, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12347(w_eco12347, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12348(w_eco12348, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12349(w_eco12349, Tsync[0], Tsync[7], prev_cnt[6], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12350(w_eco12350, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12351(w_eco12351, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12352(w_eco12352, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12353(w_eco12353, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12354(w_eco12354, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12355(w_eco12355, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12356(w_eco12356, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12357(w_eco12357, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12358(w_eco12358, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12359(w_eco12359, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12360(w_eco12360, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12361(w_eco12361, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12362(w_eco12362, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12363(w_eco12363, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12364(w_eco12364, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12365(w_eco12365, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12366(w_eco12366, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12367(w_eco12367, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12368(w_eco12368, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12369(w_eco12369, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12370(w_eco12370, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12371(w_eco12371, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12372(w_eco12372, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12373(w_eco12373, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12374(w_eco12374, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12375(w_eco12375, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12376(w_eco12376, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12377(w_eco12377, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12378(w_eco12378, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12379(w_eco12379, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12380(w_eco12380, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12381(w_eco12381, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12382(w_eco12382, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12383(w_eco12383, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12384(w_eco12384, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12385(w_eco12385, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12386(w_eco12386, !prev_cnt[14], !prev_cnt[0], prev_cnt[4], prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_12387(w_eco12387, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[12], ena, prev_state[1], !prev_state[0]);
	and _ECO_12388(w_eco12388, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12389(w_eco12389, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12390(w_eco12390, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12391(w_eco12391, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12392(w_eco12392, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12393(w_eco12393, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12394(w_eco12394, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12395(w_eco12395, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12396(w_eco12396, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12397(w_eco12397, prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12398(w_eco12398, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12399(w_eco12399, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12400(w_eco12400, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12401(w_eco12401, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12402(w_eco12402, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12403(w_eco12403, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12404(w_eco12404, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12405(w_eco12405, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12406(w_eco12406, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12407(w_eco12407, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12408(w_eco12408, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12409(w_eco12409, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12410(w_eco12410, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12411(w_eco12411, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12412(w_eco12412, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12413(w_eco12413, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12414(w_eco12414, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12415(w_eco12415, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12416(w_eco12416, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12417(w_eco12417, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12418(w_eco12418, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12419(w_eco12419, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12420(w_eco12420, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12421(w_eco12421, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12422(w_eco12422, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12423(w_eco12423, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12424(w_eco12424, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12425(w_eco12425, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12426(w_eco12426, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12427(w_eco12427, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12428(w_eco12428, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12429(w_eco12429, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12430(w_eco12430, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12431(w_eco12431, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12432(w_eco12432, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12433(w_eco12433, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12434(w_eco12434, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12435(w_eco12435, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12436(w_eco12436, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12437(w_eco12437, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12438(w_eco12438, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12439(w_eco12439, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12440(w_eco12440, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12441(w_eco12441, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12442(w_eco12442, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12443(w_eco12443, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12444(w_eco12444, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12445(w_eco12445, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12446(w_eco12446, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12447(w_eco12447, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12448(w_eco12448, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12449(w_eco12449, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12450(w_eco12450, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12451(w_eco12451, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12452(w_eco12452, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12453(w_eco12453, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12454(w_eco12454, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12455(w_eco12455, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12456(w_eco12456, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12457(w_eco12457, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12458(w_eco12458, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12459(w_eco12459, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12460(w_eco12460, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12461(w_eco12461, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12462(w_eco12462, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12463(w_eco12463, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12464(w_eco12464, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12465(w_eco12465, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12466(w_eco12466, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[3], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12467(w_eco12467, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12468(w_eco12468, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12469(w_eco12469, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12470(w_eco12470, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12471(w_eco12471, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12472(w_eco12472, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12473(w_eco12473, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12474(w_eco12474, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12475(w_eco12475, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12476(w_eco12476, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_12477(w_eco12477, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12478(w_eco12478, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12479(w_eco12479, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12480(w_eco12480, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12481(w_eco12481, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12482(w_eco12482, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12483(w_eco12483, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12484(w_eco12484, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12485(w_eco12485, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12486(w_eco12486, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12487(w_eco12487, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12488(w_eco12488, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12489(w_eco12489, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12490(w_eco12490, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12491(w_eco12491, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12492(w_eco12492, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12493(w_eco12493, Tsync[7], prev_cnt[0], prev_cnt[6], !prev_cnt[7], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12494(w_eco12494, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12495(w_eco12495, !prev_cnt[14], !prev_cnt[0], prev_cnt[5], prev_cnt[7], prev_cnt[13], ena, prev_state[1], !prev_state[0]);
	and _ECO_12496(w_eco12496, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12497(w_eco12497, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12498(w_eco12498, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12499(w_eco12499, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12500(w_eco12500, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12501(w_eco12501, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12502(w_eco12502, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12503(w_eco12503, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12504(w_eco12504, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12505(w_eco12505, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12506(w_eco12506, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12507(w_eco12507, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12508(w_eco12508, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12509(w_eco12509, prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12510(w_eco12510, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12511(w_eco12511, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12512(w_eco12512, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12513(w_eco12513, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12514(w_eco12514, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12515(w_eco12515, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12516(w_eco12516, !prev_cnt[0], prev_cnt[1], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12517(w_eco12517, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12518(w_eco12518, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12519(w_eco12519, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12520(w_eco12520, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12521(w_eco12521, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12522(w_eco12522, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12523(w_eco12523, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12524(w_eco12524, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12525(w_eco12525, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12526(w_eco12526, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12527(w_eco12527, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12528(w_eco12528, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12529(w_eco12529, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12530(w_eco12530, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12531(w_eco12531, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12532(w_eco12532, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12533(w_eco12533, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12534(w_eco12534, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12535(w_eco12535, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12536(w_eco12536, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12537(w_eco12537, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12538(w_eco12538, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12539(w_eco12539, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12540(w_eco12540, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12541(w_eco12541, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12542(w_eco12542, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12543(w_eco12543, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12544(w_eco12544, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12545(w_eco12545, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12546(w_eco12546, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12547(w_eco12547, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12548(w_eco12548, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12549(w_eco12549, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12550(w_eco12550, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12551(w_eco12551, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12552(w_eco12552, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12553(w_eco12553, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12554(w_eco12554, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12555(w_eco12555, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12556(w_eco12556, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12557(w_eco12557, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12558(w_eco12558, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12559(w_eco12559, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12560(w_eco12560, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12561(w_eco12561, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12562(w_eco12562, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12563(w_eco12563, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12564(w_eco12564, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12565(w_eco12565, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12566(w_eco12566, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12567(w_eco12567, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12568(w_eco12568, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12569(w_eco12569, Tsync[0], Tsync[7], prev_cnt[1], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12570(w_eco12570, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12571(w_eco12571, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12572(w_eco12572, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12573(w_eco12573, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12574(w_eco12574, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[11], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12575(w_eco12575, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12576(w_eco12576, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12577(w_eco12577, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[0], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12578(w_eco12578, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12579(w_eco12579, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12580(w_eco12580, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12581(w_eco12581, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12582(w_eco12582, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12583(w_eco12583, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12584(w_eco12584, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12585(w_eco12585, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12586(w_eco12586, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12587(w_eco12587, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12588(w_eco12588, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12589(w_eco12589, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12590(w_eco12590, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12591(w_eco12591, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12592(w_eco12592, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12593(w_eco12593, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12594(w_eco12594, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12595(w_eco12595, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12596(w_eco12596, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12597(w_eco12597, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12598(w_eco12598, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12599(w_eco12599, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12600(w_eco12600, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12601(w_eco12601, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12602(w_eco12602, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12603(w_eco12603, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12604(w_eco12604, prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12605(w_eco12605, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12606(w_eco12606, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12607(w_eco12607, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12608(w_eco12608, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12609(w_eco12609, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12610(w_eco12610, !prev_cnt[0], prev_cnt[2], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12611(w_eco12611, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12612(w_eco12612, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12613(w_eco12613, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12614(w_eco12614, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12615(w_eco12615, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12616(w_eco12616, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12617(w_eco12617, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12618(w_eco12618, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12619(w_eco12619, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12620(w_eco12620, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12621(w_eco12621, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12622(w_eco12622, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12623(w_eco12623, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12624(w_eco12624, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12625(w_eco12625, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12626(w_eco12626, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12627(w_eco12627, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12628(w_eco12628, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12629(w_eco12629, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12630(w_eco12630, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12631(w_eco12631, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_12632(w_eco12632, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12633(w_eco12633, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12634(w_eco12634, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12635(w_eco12635, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12636(w_eco12636, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12637(w_eco12637, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12638(w_eco12638, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12639(w_eco12639, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12640(w_eco12640, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12641(w_eco12641, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12642(w_eco12642, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12643(w_eco12643, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12644(w_eco12644, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12645(w_eco12645, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12646(w_eco12646, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12647(w_eco12647, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12648(w_eco12648, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12649(w_eco12649, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12650(w_eco12650, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12651(w_eco12651, Tsync[0], Tsync[7], prev_cnt[2], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12652(w_eco12652, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12653(w_eco12653, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12654(w_eco12654, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12655(w_eco12655, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[15], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12656(w_eco12656, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[4], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12657(w_eco12657, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12658(w_eco12658, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12659(w_eco12659, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12660(w_eco12660, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12661(w_eco12661, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12662(w_eco12662, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12663(w_eco12663, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12664(w_eco12664, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12665(w_eco12665, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12666(w_eco12666, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12667(w_eco12667, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12668(w_eco12668, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12669(w_eco12669, Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12670(w_eco12670, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12671(w_eco12671, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_12672(w_eco12672, !Tgate[7], !Tsync[7], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12673(w_eco12673, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12674(w_eco12674, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12675(w_eco12675, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12676(w_eco12676, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12677(w_eco12677, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12678(w_eco12678, !prev_cnt[0], prev_cnt[3], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12679(w_eco12679, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12680(w_eco12680, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12681(w_eco12681, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12682(w_eco12682, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12683(w_eco12683, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12684(w_eco12684, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12685(w_eco12685, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12686(w_eco12686, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12687(w_eco12687, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12688(w_eco12688, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12689(w_eco12689, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12690(w_eco12690, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12691(w_eco12691, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12692(w_eco12692, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12693(w_eco12693, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12694(w_eco12694, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12695(w_eco12695, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12696(w_eco12696, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12697(w_eco12697, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12698(w_eco12698, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12699(w_eco12699, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12700(w_eco12700, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12701(w_eco12701, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12702(w_eco12702, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12703(w_eco12703, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12704(w_eco12704, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12705(w_eco12705, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12706(w_eco12706, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12707(w_eco12707, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12708(w_eco12708, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12709(w_eco12709, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[1], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12710(w_eco12710, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12711(w_eco12711, Tsync[0], Tsync[7], prev_cnt[3], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12712(w_eco12712, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12713(w_eco12713, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12714(w_eco12714, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], prev_cnt[5], !prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12715(w_eco12715, Tsync[0], !Tgate[7], !Tgdel[7], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12716(w_eco12716, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12717(w_eco12717, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12718(w_eco12718, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12719(w_eco12719, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12720(w_eco12720, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12721(w_eco12721, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12722(w_eco12722, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12723(w_eco12723, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12724(w_eco12724, !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[3], !prev_state[1], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12725(w_eco12725, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12726(w_eco12726, !prev_cnt[0], prev_cnt[4], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12727(w_eco12727, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12728(w_eco12728, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12729(w_eco12729, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12730(w_eco12730, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12731(w_eco12731, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12732(w_eco12732, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12733(w_eco12733, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12734(w_eco12734, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12735(w_eco12735, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12736(w_eco12736, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12737(w_eco12737, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12738(w_eco12738, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12739(w_eco12739, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12740(w_eco12740, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12741(w_eco12741, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12742(w_eco12742, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12743(w_eco12743, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12744(w_eco12744, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12745(w_eco12745, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12746(w_eco12746, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12747(w_eco12747, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12748(w_eco12748, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[2], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12749(w_eco12749, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12750(w_eco12750, Tsync[0], Tsync[7], prev_cnt[0], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12751(w_eco12751, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12752(w_eco12752, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12753(w_eco12753, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[9], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12754(w_eco12754, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12755(w_eco12755, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12756(w_eco12756, Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, !prev_state[3], prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12757(w_eco12757, !Tgate[7], !Tsync[7], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_12758(w_eco12758, !prev_cnt[0], prev_cnt[5], prev_cnt[7], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12759(w_eco12759, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12760(w_eco12760, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12761(w_eco12761, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12762(w_eco12762, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12763(w_eco12763, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12764(w_eco12764, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12765(w_eco12765, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12766(w_eco12766, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12767(w_eco12767, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12768(w_eco12768, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12769(w_eco12769, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12770(w_eco12770, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12771(w_eco12771, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12772(w_eco12772, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12773(w_eco12773, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[3], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12774(w_eco12774, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12775(w_eco12775, Tsync[0], Tsync[7], prev_cnt[4], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12776(w_eco12776, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12777(w_eco12777, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[8], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12778(w_eco12778, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12779(w_eco12779, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12780(w_eco12780, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12781(w_eco12781, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12782(w_eco12782, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12783(w_eco12783, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12784(w_eco12784, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_12785(w_eco12785, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[0], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12786(w_eco12786, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12787(w_eco12787, Tsync[0], Tsync[7], prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12788(w_eco12788, Tsync[0], Tsync[7], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[10], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12789(w_eco12789, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12790(w_eco12790, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12791(w_eco12791, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[4], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12792(w_eco12792, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12793(w_eco12793, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[12], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12794(w_eco12794, Tsync[0], Tsync[7], !prev_cnt[14], prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_12795(w_eco12795, Tsync[0], Tsync[7], !prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], prev_cnt[7], prev_cnt[13], ena, prev_state[2], !prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_12796(w_eco12796, w_eco10926, w_eco10927, w_eco10928, w_eco10929, w_eco10930, w_eco10931, w_eco10932, w_eco10933, w_eco10934, w_eco10935, w_eco10936, w_eco10937, w_eco10938, w_eco10939, w_eco10940, w_eco10941, w_eco10942, w_eco10943, w_eco10944, w_eco10945, w_eco10946, w_eco10947, w_eco10948, w_eco10949, w_eco10950, w_eco10951, w_eco10952, w_eco10953, w_eco10954, w_eco10955, w_eco10956, w_eco10957, w_eco10958, w_eco10959, w_eco10960, w_eco10961, w_eco10962, w_eco10963, w_eco10964, w_eco10965, w_eco10966, w_eco10967, w_eco10968, w_eco10969, w_eco10970, w_eco10971, w_eco10972, w_eco10973, w_eco10974, w_eco10975, w_eco10976, w_eco10977, w_eco10978, w_eco10979, w_eco10980, w_eco10981, w_eco10982, w_eco10983, w_eco10984, w_eco10985, w_eco10986, w_eco10987, w_eco10988, w_eco10989, w_eco10990, w_eco10991, w_eco10992, w_eco10993, w_eco10994, w_eco10995, w_eco10996, w_eco10997, w_eco10998, w_eco10999, w_eco11000, w_eco11001, w_eco11002, w_eco11003, w_eco11004, w_eco11005, w_eco11006, w_eco11007, w_eco11008, w_eco11009, w_eco11010, w_eco11011, w_eco11012, w_eco11013, w_eco11014, w_eco11015, w_eco11016, w_eco11017, w_eco11018, w_eco11019, w_eco11020, w_eco11021, w_eco11022, w_eco11023, w_eco11024, w_eco11025, w_eco11026, w_eco11027, w_eco11028, w_eco11029, w_eco11030, w_eco11031, w_eco11032, w_eco11033, w_eco11034, w_eco11035, w_eco11036, w_eco11037, w_eco11038, w_eco11039, w_eco11040, w_eco11041, w_eco11042, w_eco11043, w_eco11044, w_eco11045, w_eco11046, w_eco11047, w_eco11048, w_eco11049, w_eco11050, w_eco11051, w_eco11052, w_eco11053, w_eco11054, w_eco11055, w_eco11056, w_eco11057, w_eco11058, w_eco11059, w_eco11060, w_eco11061, w_eco11062, w_eco11063, w_eco11064, w_eco11065, w_eco11066, w_eco11067, w_eco11068, w_eco11069, w_eco11070, w_eco11071, w_eco11072, w_eco11073, w_eco11074, w_eco11075, w_eco11076, w_eco11077, w_eco11078, w_eco11079, w_eco11080, w_eco11081, w_eco11082, w_eco11083, w_eco11084, w_eco11085, w_eco11086, w_eco11087, w_eco11088, w_eco11089, w_eco11090, w_eco11091, w_eco11092, w_eco11093, w_eco11094, w_eco11095, w_eco11096, w_eco11097, w_eco11098, w_eco11099, w_eco11100, w_eco11101, w_eco11102, w_eco11103, w_eco11104, w_eco11105, w_eco11106, w_eco11107, w_eco11108, w_eco11109, w_eco11110, w_eco11111, w_eco11112, w_eco11113, w_eco11114, w_eco11115, w_eco11116, w_eco11117, w_eco11118, w_eco11119, w_eco11120, w_eco11121, w_eco11122, w_eco11123, w_eco11124, w_eco11125, w_eco11126, w_eco11127, w_eco11128, w_eco11129, w_eco11130, w_eco11131, w_eco11132, w_eco11133, w_eco11134, w_eco11135, w_eco11136, w_eco11137, w_eco11138, w_eco11139, w_eco11140, w_eco11141, w_eco11142, w_eco11143, w_eco11144, w_eco11145, w_eco11146, w_eco11147, w_eco11148, w_eco11149, w_eco11150, w_eco11151, w_eco11152, w_eco11153, w_eco11154, w_eco11155, w_eco11156, w_eco11157, w_eco11158, w_eco11159, w_eco11160, w_eco11161, w_eco11162, w_eco11163, w_eco11164, w_eco11165, w_eco11166, w_eco11167, w_eco11168, w_eco11169, w_eco11170, w_eco11171, w_eco11172, w_eco11173, w_eco11174, w_eco11175, w_eco11176, w_eco11177, w_eco11178, w_eco11179, w_eco11180, w_eco11181, w_eco11182, w_eco11183, w_eco11184, w_eco11185, w_eco11186, w_eco11187, w_eco11188, w_eco11189, w_eco11190, w_eco11191, w_eco11192, w_eco11193, w_eco11194, w_eco11195, w_eco11196, w_eco11197, w_eco11198, w_eco11199, w_eco11200, w_eco11201, w_eco11202, w_eco11203, w_eco11204, w_eco11205, w_eco11206, w_eco11207, w_eco11208, w_eco11209, w_eco11210, w_eco11211, w_eco11212, w_eco11213, w_eco11214, w_eco11215, w_eco11216, w_eco11217, w_eco11218, w_eco11219, w_eco11220, w_eco11221, w_eco11222, w_eco11223, w_eco11224, w_eco11225, w_eco11226, w_eco11227, w_eco11228, w_eco11229, w_eco11230, w_eco11231, w_eco11232, w_eco11233, w_eco11234, w_eco11235, w_eco11236, w_eco11237, w_eco11238, w_eco11239, w_eco11240, w_eco11241, w_eco11242, w_eco11243, w_eco11244, w_eco11245, w_eco11246, w_eco11247, w_eco11248, w_eco11249, w_eco11250, w_eco11251, w_eco11252, w_eco11253, w_eco11254, w_eco11255, w_eco11256, w_eco11257, w_eco11258, w_eco11259, w_eco11260, w_eco11261, w_eco11262, w_eco11263, w_eco11264, w_eco11265, w_eco11266, w_eco11267, w_eco11268, w_eco11269, w_eco11270, w_eco11271, w_eco11272, w_eco11273, w_eco11274, w_eco11275, w_eco11276, w_eco11277, w_eco11278, w_eco11279, w_eco11280, w_eco11281, w_eco11282, w_eco11283, w_eco11284, w_eco11285, w_eco11286, w_eco11287, w_eco11288, w_eco11289, w_eco11290, w_eco11291, w_eco11292, w_eco11293, w_eco11294, w_eco11295, w_eco11296, w_eco11297, w_eco11298, w_eco11299, w_eco11300, w_eco11301, w_eco11302, w_eco11303, w_eco11304, w_eco11305, w_eco11306, w_eco11307, w_eco11308, w_eco11309, w_eco11310, w_eco11311, w_eco11312, w_eco11313, w_eco11314, w_eco11315, w_eco11316, w_eco11317, w_eco11318, w_eco11319, w_eco11320, w_eco11321, w_eco11322, w_eco11323, w_eco11324, w_eco11325, w_eco11326, w_eco11327, w_eco11328, w_eco11329, w_eco11330, w_eco11331, w_eco11332, w_eco11333, w_eco11334, w_eco11335, w_eco11336, w_eco11337, w_eco11338, w_eco11339, w_eco11340, w_eco11341, w_eco11342, w_eco11343, w_eco11344, w_eco11345, w_eco11346, w_eco11347, w_eco11348, w_eco11349, w_eco11350, w_eco11351, w_eco11352, w_eco11353, w_eco11354, w_eco11355, w_eco11356, w_eco11357, w_eco11358, w_eco11359, w_eco11360, w_eco11361, w_eco11362, w_eco11363, w_eco11364, w_eco11365, w_eco11366, w_eco11367, w_eco11368, w_eco11369, w_eco11370, w_eco11371, w_eco11372, w_eco11373, w_eco11374, w_eco11375, w_eco11376, w_eco11377, w_eco11378, w_eco11379, w_eco11380, w_eco11381, w_eco11382, w_eco11383, w_eco11384, w_eco11385, w_eco11386, w_eco11387, w_eco11388, w_eco11389, w_eco11390, w_eco11391, w_eco11392, w_eco11393, w_eco11394, w_eco11395, w_eco11396, w_eco11397, w_eco11398, w_eco11399, w_eco11400, w_eco11401, w_eco11402, w_eco11403, w_eco11404, w_eco11405, w_eco11406, w_eco11407, w_eco11408, w_eco11409, w_eco11410, w_eco11411, w_eco11412, w_eco11413, w_eco11414, w_eco11415, w_eco11416, w_eco11417, w_eco11418, w_eco11419, w_eco11420, w_eco11421, w_eco11422, w_eco11423, w_eco11424, w_eco11425, w_eco11426, w_eco11427, w_eco11428, w_eco11429, w_eco11430, w_eco11431, w_eco11432, w_eco11433, w_eco11434, w_eco11435, w_eco11436, w_eco11437, w_eco11438, w_eco11439, w_eco11440, w_eco11441, w_eco11442, w_eco11443, w_eco11444, w_eco11445, w_eco11446, w_eco11447, w_eco11448, w_eco11449, w_eco11450, w_eco11451, w_eco11452, w_eco11453, w_eco11454, w_eco11455, w_eco11456, w_eco11457, w_eco11458, w_eco11459, w_eco11460, w_eco11461, w_eco11462, w_eco11463, w_eco11464, w_eco11465, w_eco11466, w_eco11467, w_eco11468, w_eco11469, w_eco11470, w_eco11471, w_eco11472, w_eco11473, w_eco11474, w_eco11475, w_eco11476, w_eco11477, w_eco11478, w_eco11479, w_eco11480, w_eco11481, w_eco11482, w_eco11483, w_eco11484, w_eco11485, w_eco11486, w_eco11487, w_eco11488, w_eco11489, w_eco11490, w_eco11491, w_eco11492, w_eco11493, w_eco11494, w_eco11495, w_eco11496, w_eco11497, w_eco11498, w_eco11499, w_eco11500, w_eco11501, w_eco11502, w_eco11503, w_eco11504, w_eco11505, w_eco11506, w_eco11507, w_eco11508, w_eco11509, w_eco11510, w_eco11511, w_eco11512, w_eco11513, w_eco11514, w_eco11515, w_eco11516, w_eco11517, w_eco11518, w_eco11519, w_eco11520, w_eco11521, w_eco11522, w_eco11523, w_eco11524, w_eco11525, w_eco11526, w_eco11527, w_eco11528, w_eco11529, w_eco11530, w_eco11531, w_eco11532, w_eco11533, w_eco11534, w_eco11535, w_eco11536, w_eco11537, w_eco11538, w_eco11539, w_eco11540, w_eco11541, w_eco11542, w_eco11543, w_eco11544, w_eco11545, w_eco11546, w_eco11547, w_eco11548, w_eco11549, w_eco11550, w_eco11551, w_eco11552, w_eco11553, w_eco11554, w_eco11555, w_eco11556, w_eco11557, w_eco11558, w_eco11559, w_eco11560, w_eco11561, w_eco11562, w_eco11563, w_eco11564, w_eco11565, w_eco11566, w_eco11567, w_eco11568, w_eco11569, w_eco11570, w_eco11571, w_eco11572, w_eco11573, w_eco11574, w_eco11575, w_eco11576, w_eco11577, w_eco11578, w_eco11579, w_eco11580, w_eco11581, w_eco11582, w_eco11583, w_eco11584, w_eco11585, w_eco11586, w_eco11587, w_eco11588, w_eco11589, w_eco11590, w_eco11591, w_eco11592, w_eco11593, w_eco11594, w_eco11595, w_eco11596, w_eco11597, w_eco11598, w_eco11599, w_eco11600, w_eco11601, w_eco11602, w_eco11603, w_eco11604, w_eco11605, w_eco11606, w_eco11607, w_eco11608, w_eco11609, w_eco11610, w_eco11611, w_eco11612, w_eco11613, w_eco11614, w_eco11615, w_eco11616, w_eco11617, w_eco11618, w_eco11619, w_eco11620, w_eco11621, w_eco11622, w_eco11623, w_eco11624, w_eco11625, w_eco11626, w_eco11627, w_eco11628, w_eco11629, w_eco11630, w_eco11631, w_eco11632, w_eco11633, w_eco11634, w_eco11635, w_eco11636, w_eco11637, w_eco11638, w_eco11639, w_eco11640, w_eco11641, w_eco11642, w_eco11643, w_eco11644, w_eco11645, w_eco11646, w_eco11647, w_eco11648, w_eco11649, w_eco11650, w_eco11651, w_eco11652, w_eco11653, w_eco11654, w_eco11655, w_eco11656, w_eco11657, w_eco11658, w_eco11659, w_eco11660, w_eco11661, w_eco11662, w_eco11663, w_eco11664, w_eco11665, w_eco11666, w_eco11667, w_eco11668, w_eco11669, w_eco11670, w_eco11671, w_eco11672, w_eco11673, w_eco11674, w_eco11675, w_eco11676, w_eco11677, w_eco11678, w_eco11679, w_eco11680, w_eco11681, w_eco11682, w_eco11683, w_eco11684, w_eco11685, w_eco11686, w_eco11687, w_eco11688, w_eco11689, w_eco11690, w_eco11691, w_eco11692, w_eco11693, w_eco11694, w_eco11695, w_eco11696, w_eco11697, w_eco11698, w_eco11699, w_eco11700, w_eco11701, w_eco11702, w_eco11703, w_eco11704, w_eco11705, w_eco11706, w_eco11707, w_eco11708, w_eco11709, w_eco11710, w_eco11711, w_eco11712, w_eco11713, w_eco11714, w_eco11715, w_eco11716, w_eco11717, w_eco11718, w_eco11719, w_eco11720, w_eco11721, w_eco11722, w_eco11723, w_eco11724, w_eco11725, w_eco11726, w_eco11727, w_eco11728, w_eco11729, w_eco11730, w_eco11731, w_eco11732, w_eco11733, w_eco11734, w_eco11735, w_eco11736, w_eco11737, w_eco11738, w_eco11739, w_eco11740, w_eco11741, w_eco11742, w_eco11743, w_eco11744, w_eco11745, w_eco11746, w_eco11747, w_eco11748, w_eco11749, w_eco11750, w_eco11751, w_eco11752, w_eco11753, w_eco11754, w_eco11755, w_eco11756, w_eco11757, w_eco11758, w_eco11759, w_eco11760, w_eco11761, w_eco11762, w_eco11763, w_eco11764, w_eco11765, w_eco11766, w_eco11767, w_eco11768, w_eco11769, w_eco11770, w_eco11771, w_eco11772, w_eco11773, w_eco11774, w_eco11775, w_eco11776, w_eco11777, w_eco11778, w_eco11779, w_eco11780, w_eco11781, w_eco11782, w_eco11783, w_eco11784, w_eco11785, w_eco11786, w_eco11787, w_eco11788, w_eco11789, w_eco11790, w_eco11791, w_eco11792, w_eco11793, w_eco11794, w_eco11795, w_eco11796, w_eco11797, w_eco11798, w_eco11799, w_eco11800, w_eco11801, w_eco11802, w_eco11803, w_eco11804, w_eco11805, w_eco11806, w_eco11807, w_eco11808, w_eco11809, w_eco11810, w_eco11811, w_eco11812, w_eco11813, w_eco11814, w_eco11815, w_eco11816, w_eco11817, w_eco11818, w_eco11819, w_eco11820, w_eco11821, w_eco11822, w_eco11823, w_eco11824, w_eco11825, w_eco11826, w_eco11827, w_eco11828, w_eco11829, w_eco11830, w_eco11831, w_eco11832, w_eco11833, w_eco11834, w_eco11835, w_eco11836, w_eco11837, w_eco11838, w_eco11839, w_eco11840, w_eco11841, w_eco11842, w_eco11843, w_eco11844, w_eco11845, w_eco11846, w_eco11847, w_eco11848, w_eco11849, w_eco11850, w_eco11851, w_eco11852, w_eco11853, w_eco11854, w_eco11855, w_eco11856, w_eco11857, w_eco11858, w_eco11859, w_eco11860, w_eco11861, w_eco11862, w_eco11863, w_eco11864, w_eco11865, w_eco11866, w_eco11867, w_eco11868, w_eco11869, w_eco11870, w_eco11871, w_eco11872, w_eco11873, w_eco11874, w_eco11875, w_eco11876, w_eco11877, w_eco11878, w_eco11879, w_eco11880, w_eco11881, w_eco11882, w_eco11883, w_eco11884, w_eco11885, w_eco11886, w_eco11887, w_eco11888, w_eco11889, w_eco11890, w_eco11891, w_eco11892, w_eco11893, w_eco11894, w_eco11895, w_eco11896, w_eco11897, w_eco11898, w_eco11899, w_eco11900, w_eco11901, w_eco11902, w_eco11903, w_eco11904, w_eco11905, w_eco11906, w_eco11907, w_eco11908, w_eco11909, w_eco11910, w_eco11911, w_eco11912, w_eco11913, w_eco11914, w_eco11915, w_eco11916, w_eco11917, w_eco11918, w_eco11919, w_eco11920, w_eco11921, w_eco11922, w_eco11923, w_eco11924, w_eco11925, w_eco11926, w_eco11927, w_eco11928, w_eco11929, w_eco11930, w_eco11931, w_eco11932, w_eco11933, w_eco11934, w_eco11935, w_eco11936, w_eco11937, w_eco11938, w_eco11939, w_eco11940, w_eco11941, w_eco11942, w_eco11943, w_eco11944, w_eco11945, w_eco11946, w_eco11947, w_eco11948, w_eco11949, w_eco11950, w_eco11951, w_eco11952, w_eco11953, w_eco11954, w_eco11955, w_eco11956, w_eco11957, w_eco11958, w_eco11959, w_eco11960, w_eco11961, w_eco11962, w_eco11963, w_eco11964, w_eco11965, w_eco11966, w_eco11967, w_eco11968, w_eco11969, w_eco11970, w_eco11971, w_eco11972, w_eco11973, w_eco11974, w_eco11975, w_eco11976, w_eco11977, w_eco11978, w_eco11979, w_eco11980, w_eco11981, w_eco11982, w_eco11983, w_eco11984, w_eco11985, w_eco11986, w_eco11987, w_eco11988, w_eco11989, w_eco11990, w_eco11991, w_eco11992, w_eco11993, w_eco11994, w_eco11995, w_eco11996, w_eco11997, w_eco11998, w_eco11999, w_eco12000, w_eco12001, w_eco12002, w_eco12003, w_eco12004, w_eco12005, w_eco12006, w_eco12007, w_eco12008, w_eco12009, w_eco12010, w_eco12011, w_eco12012, w_eco12013, w_eco12014, w_eco12015, w_eco12016, w_eco12017, w_eco12018, w_eco12019, w_eco12020, w_eco12021, w_eco12022, w_eco12023, w_eco12024, w_eco12025, w_eco12026, w_eco12027, w_eco12028, w_eco12029, w_eco12030, w_eco12031, w_eco12032, w_eco12033, w_eco12034, w_eco12035, w_eco12036, w_eco12037, w_eco12038, w_eco12039, w_eco12040, w_eco12041, w_eco12042, w_eco12043, w_eco12044, w_eco12045, w_eco12046, w_eco12047, w_eco12048, w_eco12049, w_eco12050, w_eco12051, w_eco12052, w_eco12053, w_eco12054, w_eco12055, w_eco12056, w_eco12057, w_eco12058, w_eco12059, w_eco12060, w_eco12061, w_eco12062, w_eco12063, w_eco12064, w_eco12065, w_eco12066, w_eco12067, w_eco12068, w_eco12069, w_eco12070, w_eco12071, w_eco12072, w_eco12073, w_eco12074, w_eco12075, w_eco12076, w_eco12077, w_eco12078, w_eco12079, w_eco12080, w_eco12081, w_eco12082, w_eco12083, w_eco12084, w_eco12085, w_eco12086, w_eco12087, w_eco12088, w_eco12089, w_eco12090, w_eco12091, w_eco12092, w_eco12093, w_eco12094, w_eco12095, w_eco12096, w_eco12097, w_eco12098, w_eco12099, w_eco12100, w_eco12101, w_eco12102, w_eco12103, w_eco12104, w_eco12105, w_eco12106, w_eco12107, w_eco12108, w_eco12109, w_eco12110, w_eco12111, w_eco12112, w_eco12113, w_eco12114, w_eco12115, w_eco12116, w_eco12117, w_eco12118, w_eco12119, w_eco12120, w_eco12121, w_eco12122, w_eco12123, w_eco12124, w_eco12125, w_eco12126, w_eco12127, w_eco12128, w_eco12129, w_eco12130, w_eco12131, w_eco12132, w_eco12133, w_eco12134, w_eco12135, w_eco12136, w_eco12137, w_eco12138, w_eco12139, w_eco12140, w_eco12141, w_eco12142, w_eco12143, w_eco12144, w_eco12145, w_eco12146, w_eco12147, w_eco12148, w_eco12149, w_eco12150, w_eco12151, w_eco12152, w_eco12153, w_eco12154, w_eco12155, w_eco12156, w_eco12157, w_eco12158, w_eco12159, w_eco12160, w_eco12161, w_eco12162, w_eco12163, w_eco12164, w_eco12165, w_eco12166, w_eco12167, w_eco12168, w_eco12169, w_eco12170, w_eco12171, w_eco12172, w_eco12173, w_eco12174, w_eco12175, w_eco12176, w_eco12177, w_eco12178, w_eco12179, w_eco12180, w_eco12181, w_eco12182, w_eco12183, w_eco12184, w_eco12185, w_eco12186, w_eco12187, w_eco12188, w_eco12189, w_eco12190, w_eco12191, w_eco12192, w_eco12193, w_eco12194, w_eco12195, w_eco12196, w_eco12197, w_eco12198, w_eco12199, w_eco12200, w_eco12201, w_eco12202, w_eco12203, w_eco12204, w_eco12205, w_eco12206, w_eco12207, w_eco12208, w_eco12209, w_eco12210, w_eco12211, w_eco12212, w_eco12213, w_eco12214, w_eco12215, w_eco12216, w_eco12217, w_eco12218, w_eco12219, w_eco12220, w_eco12221, w_eco12222, w_eco12223, w_eco12224, w_eco12225, w_eco12226, w_eco12227, w_eco12228, w_eco12229, w_eco12230, w_eco12231, w_eco12232, w_eco12233, w_eco12234, w_eco12235, w_eco12236, w_eco12237, w_eco12238, w_eco12239, w_eco12240, w_eco12241, w_eco12242, w_eco12243, w_eco12244, w_eco12245, w_eco12246, w_eco12247, w_eco12248, w_eco12249, w_eco12250, w_eco12251, w_eco12252, w_eco12253, w_eco12254, w_eco12255, w_eco12256, w_eco12257, w_eco12258, w_eco12259, w_eco12260, w_eco12261, w_eco12262, w_eco12263, w_eco12264, w_eco12265, w_eco12266, w_eco12267, w_eco12268, w_eco12269, w_eco12270, w_eco12271, w_eco12272, w_eco12273, w_eco12274, w_eco12275, w_eco12276, w_eco12277, w_eco12278, w_eco12279, w_eco12280, w_eco12281, w_eco12282, w_eco12283, w_eco12284, w_eco12285, w_eco12286, w_eco12287, w_eco12288, w_eco12289, w_eco12290, w_eco12291, w_eco12292, w_eco12293, w_eco12294, w_eco12295, w_eco12296, w_eco12297, w_eco12298, w_eco12299, w_eco12300, w_eco12301, w_eco12302, w_eco12303, w_eco12304, w_eco12305, w_eco12306, w_eco12307, w_eco12308, w_eco12309, w_eco12310, w_eco12311, w_eco12312, w_eco12313, w_eco12314, w_eco12315, w_eco12316, w_eco12317, w_eco12318, w_eco12319, w_eco12320, w_eco12321, w_eco12322, w_eco12323, w_eco12324, w_eco12325, w_eco12326, w_eco12327, w_eco12328, w_eco12329, w_eco12330, w_eco12331, w_eco12332, w_eco12333, w_eco12334, w_eco12335, w_eco12336, w_eco12337, w_eco12338, w_eco12339, w_eco12340, w_eco12341, w_eco12342, w_eco12343, w_eco12344, w_eco12345, w_eco12346, w_eco12347, w_eco12348, w_eco12349, w_eco12350, w_eco12351, w_eco12352, w_eco12353, w_eco12354, w_eco12355, w_eco12356, w_eco12357, w_eco12358, w_eco12359, w_eco12360, w_eco12361, w_eco12362, w_eco12363, w_eco12364, w_eco12365, w_eco12366, w_eco12367, w_eco12368, w_eco12369, w_eco12370, w_eco12371, w_eco12372, w_eco12373, w_eco12374, w_eco12375, w_eco12376, w_eco12377, w_eco12378, w_eco12379, w_eco12380, w_eco12381, w_eco12382, w_eco12383, w_eco12384, w_eco12385, w_eco12386, w_eco12387, w_eco12388, w_eco12389, w_eco12390, w_eco12391, w_eco12392, w_eco12393, w_eco12394, w_eco12395, w_eco12396, w_eco12397, w_eco12398, w_eco12399, w_eco12400, w_eco12401, w_eco12402, w_eco12403, w_eco12404, w_eco12405, w_eco12406, w_eco12407, w_eco12408, w_eco12409, w_eco12410, w_eco12411, w_eco12412, w_eco12413, w_eco12414, w_eco12415, w_eco12416, w_eco12417, w_eco12418, w_eco12419, w_eco12420, w_eco12421, w_eco12422, w_eco12423, w_eco12424, w_eco12425, w_eco12426, w_eco12427, w_eco12428, w_eco12429, w_eco12430, w_eco12431, w_eco12432, w_eco12433, w_eco12434, w_eco12435, w_eco12436, w_eco12437, w_eco12438, w_eco12439, w_eco12440, w_eco12441, w_eco12442, w_eco12443, w_eco12444, w_eco12445, w_eco12446, w_eco12447, w_eco12448, w_eco12449, w_eco12450, w_eco12451, w_eco12452, w_eco12453, w_eco12454, w_eco12455, w_eco12456, w_eco12457, w_eco12458, w_eco12459, w_eco12460, w_eco12461, w_eco12462, w_eco12463, w_eco12464, w_eco12465, w_eco12466, w_eco12467, w_eco12468, w_eco12469, w_eco12470, w_eco12471, w_eco12472, w_eco12473, w_eco12474, w_eco12475, w_eco12476, w_eco12477, w_eco12478, w_eco12479, w_eco12480, w_eco12481, w_eco12482, w_eco12483, w_eco12484, w_eco12485, w_eco12486, w_eco12487, w_eco12488, w_eco12489, w_eco12490, w_eco12491, w_eco12492, w_eco12493, w_eco12494, w_eco12495, w_eco12496, w_eco12497, w_eco12498, w_eco12499, w_eco12500, w_eco12501, w_eco12502, w_eco12503, w_eco12504, w_eco12505, w_eco12506, w_eco12507, w_eco12508, w_eco12509, w_eco12510, w_eco12511, w_eco12512, w_eco12513, w_eco12514, w_eco12515, w_eco12516, w_eco12517, w_eco12518, w_eco12519, w_eco12520, w_eco12521, w_eco12522, w_eco12523, w_eco12524, w_eco12525, w_eco12526, w_eco12527, w_eco12528, w_eco12529, w_eco12530, w_eco12531, w_eco12532, w_eco12533, w_eco12534, w_eco12535, w_eco12536, w_eco12537, w_eco12538, w_eco12539, w_eco12540, w_eco12541, w_eco12542, w_eco12543, w_eco12544, w_eco12545, w_eco12546, w_eco12547, w_eco12548, w_eco12549, w_eco12550, w_eco12551, w_eco12552, w_eco12553, w_eco12554, w_eco12555, w_eco12556, w_eco12557, w_eco12558, w_eco12559, w_eco12560, w_eco12561, w_eco12562, w_eco12563, w_eco12564, w_eco12565, w_eco12566, w_eco12567, w_eco12568, w_eco12569, w_eco12570, w_eco12571, w_eco12572, w_eco12573, w_eco12574, w_eco12575, w_eco12576, w_eco12577, w_eco12578, w_eco12579, w_eco12580, w_eco12581, w_eco12582, w_eco12583, w_eco12584, w_eco12585, w_eco12586, w_eco12587, w_eco12588, w_eco12589, w_eco12590, w_eco12591, w_eco12592, w_eco12593, w_eco12594, w_eco12595, w_eco12596, w_eco12597, w_eco12598, w_eco12599, w_eco12600, w_eco12601, w_eco12602, w_eco12603, w_eco12604, w_eco12605, w_eco12606, w_eco12607, w_eco12608, w_eco12609, w_eco12610, w_eco12611, w_eco12612, w_eco12613, w_eco12614, w_eco12615, w_eco12616, w_eco12617, w_eco12618, w_eco12619, w_eco12620, w_eco12621, w_eco12622, w_eco12623, w_eco12624, w_eco12625, w_eco12626, w_eco12627, w_eco12628, w_eco12629, w_eco12630, w_eco12631, w_eco12632, w_eco12633, w_eco12634, w_eco12635, w_eco12636, w_eco12637, w_eco12638, w_eco12639, w_eco12640, w_eco12641, w_eco12642, w_eco12643, w_eco12644, w_eco12645, w_eco12646, w_eco12647, w_eco12648, w_eco12649, w_eco12650, w_eco12651, w_eco12652, w_eco12653, w_eco12654, w_eco12655, w_eco12656, w_eco12657, w_eco12658, w_eco12659, w_eco12660, w_eco12661, w_eco12662, w_eco12663, w_eco12664, w_eco12665, w_eco12666, w_eco12667, w_eco12668, w_eco12669, w_eco12670, w_eco12671, w_eco12672, w_eco12673, w_eco12674, w_eco12675, w_eco12676, w_eco12677, w_eco12678, w_eco12679, w_eco12680, w_eco12681, w_eco12682, w_eco12683, w_eco12684, w_eco12685, w_eco12686, w_eco12687, w_eco12688, w_eco12689, w_eco12690, w_eco12691, w_eco12692, w_eco12693, w_eco12694, w_eco12695, w_eco12696, w_eco12697, w_eco12698, w_eco12699, w_eco12700, w_eco12701, w_eco12702, w_eco12703, w_eco12704, w_eco12705, w_eco12706, w_eco12707, w_eco12708, w_eco12709, w_eco12710, w_eco12711, w_eco12712, w_eco12713, w_eco12714, w_eco12715, w_eco12716, w_eco12717, w_eco12718, w_eco12719, w_eco12720, w_eco12721, w_eco12722, w_eco12723, w_eco12724, w_eco12725, w_eco12726, w_eco12727, w_eco12728, w_eco12729, w_eco12730, w_eco12731, w_eco12732, w_eco12733, w_eco12734, w_eco12735, w_eco12736, w_eco12737, w_eco12738, w_eco12739, w_eco12740, w_eco12741, w_eco12742, w_eco12743, w_eco12744, w_eco12745, w_eco12746, w_eco12747, w_eco12748, w_eco12749, w_eco12750, w_eco12751, w_eco12752, w_eco12753, w_eco12754, w_eco12755, w_eco12756, w_eco12757, w_eco12758, w_eco12759, w_eco12760, w_eco12761, w_eco12762, w_eco12763, w_eco12764, w_eco12765, w_eco12766, w_eco12767, w_eco12768, w_eco12769, w_eco12770, w_eco12771, w_eco12772, w_eco12773, w_eco12774, w_eco12775, w_eco12776, w_eco12777, w_eco12778, w_eco12779, w_eco12780, w_eco12781, w_eco12782, w_eco12783, w_eco12784, w_eco12785, w_eco12786, w_eco12787, w_eco12788, w_eco12789, w_eco12790, w_eco12791, w_eco12792, w_eco12793, w_eco12794, w_eco12795);
	xor _ECO_out9(cnt[7], sub_wire9, w_eco12796);
	assign w_eco12797 = rst;
	and _ECO_12798(w_eco12798, prev_cnt[1], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12799(w_eco12799, prev_cnt[11], !prev_cnt[15], !ena);
	and _ECO_12800(w_eco12800, prev_cnt[1], prev_cnt[11], !prev_cnt[15], prev_state[1]);
	and _ECO_12801(w_eco12801, prev_cnt[1], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12802(w_eco12802, !Tgate[15], prev_cnt[14], !prev_cnt[15], !ena);
	and _ECO_12803(w_eco12803, !Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[15], prev_state[1]);
	and _ECO_12804(w_eco12804, !prev_cnt[1], prev_cnt[11], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12805(w_eco12805, prev_cnt[1], prev_cnt[11], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12806(w_eco12806, prev_cnt[14], prev_cnt[1], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12807(w_eco12807, prev_cnt[9], !prev_cnt[15], !ena);
	and _ECO_12808(w_eco12808, Tsync[1], prev_cnt[1], prev_cnt[11], !prev_cnt[15], prev_state[0]);
	and _ECO_12809(w_eco12809, prev_cnt[11], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12810(w_eco12810, !Tsync[1], prev_cnt[11], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12811(w_eco12811, !Tsync[1], !prev_cnt[1], prev_cnt[11], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12812(w_eco12812, !Tsync[1], prev_cnt[11], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12813(w_eco12813, prev_cnt[11], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12814(w_eco12814, prev_cnt[1], prev_cnt[11], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12815(w_eco12815, prev_cnt[1], prev_cnt[9], !prev_cnt[15], prev_state[1]);
	and _ECO_12816(w_eco12816, prev_cnt[14], !prev_cnt[1], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12817(w_eco12817, !Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12818(w_eco12818, !prev_cnt[1], prev_cnt[11], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12819(w_eco12819, !prev_cnt[14], prev_cnt[1], prev_cnt[12], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12820(w_eco12820, Tsync[1], prev_cnt[11], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12821(w_eco12821, prev_cnt[6], !prev_cnt[15], !ena);
	and _ECO_12822(w_eco12822, Tsync[1], !Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[15], prev_state[0]);
	and _ECO_12823(w_eco12823, prev_cnt[14], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12824(w_eco12824, !Tsync[1], prev_cnt[14], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12825(w_eco12825, !prev_cnt[1], prev_cnt[11], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12826(w_eco12826, !Tsync[1], prev_cnt[14], !prev_cnt[1], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12827(w_eco12827, !Tsync[1], prev_cnt[14], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12828(w_eco12828, prev_cnt[14], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12829(w_eco12829, !Tsync[1], !prev_cnt[1], prev_cnt[11], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12830(w_eco12830, Tsync[1], prev_cnt[11], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12831(w_eco12831, !Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12832(w_eco12832, prev_cnt[1], prev_cnt[6], !prev_cnt[15], prev_state[1]);
	and _ECO_12833(w_eco12833, !prev_cnt[1], prev_cnt[12], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12834(w_eco12834, Tsync[1], prev_cnt[11], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12835(w_eco12835, prev_cnt[1], prev_cnt[9], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12836(w_eco12836, prev_cnt[14], !prev_cnt[1], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12837(w_eco12837, Tsync[1], !Tgate[15], prev_cnt[14], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12838(w_eco12838, prev_cnt[8], !prev_cnt[15], !ena);
	and _ECO_12839(w_eco12839, Tsync[1], prev_cnt[1], prev_cnt[9], !prev_cnt[15], prev_state[0]);
	and _ECO_12840(w_eco12840, prev_cnt[12], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12841(w_eco12841, !Tsync[1], prev_cnt[12], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12842(w_eco12842, prev_cnt[14], !prev_cnt[1], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12843(w_eco12843, !Tsync[1], !prev_cnt[1], prev_cnt[12], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12844(w_eco12844, !Tsync[1], prev_cnt[12], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12845(w_eco12845, prev_cnt[12], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12846(w_eco12846, !Tsync[1], prev_cnt[14], !prev_cnt[1], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12847(w_eco12847, Tsync[1], !Tgate[15], prev_cnt[14], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12848(w_eco12848, prev_cnt[1], prev_cnt[9], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12849(w_eco12849, prev_cnt[1], prev_cnt[8], !prev_cnt[15], prev_state[1]);
	and _ECO_12850(w_eco12850, !prev_cnt[1], prev_cnt[13], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12851(w_eco12851, Tsync[1], !Tgate[15], prev_cnt[14], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12852(w_eco12852, prev_cnt[1], prev_cnt[6], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12853(w_eco12853, !prev_cnt[1], prev_cnt[12], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12854(w_eco12854, Tsync[1], prev_cnt[9], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12855(w_eco12855, prev_cnt[10], !prev_cnt[15], !ena);
	and _ECO_12856(w_eco12856, !prev_cnt[14], prev_cnt[12], !prev_cnt[15], !ena);
	and _ECO_12857(w_eco12857, Tsync[1], prev_cnt[1], prev_cnt[6], !prev_cnt[15], prev_state[0]);
	and _ECO_12858(w_eco12858, prev_cnt[13], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12859(w_eco12859, !Tsync[1], prev_cnt[13], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12860(w_eco12860, !prev_cnt[1], prev_cnt[12], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12861(w_eco12861, !Tsync[1], !prev_cnt[1], prev_cnt[13], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12862(w_eco12862, !Tsync[1], prev_cnt[13], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12863(w_eco12863, prev_cnt[13], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12864(w_eco12864, !Tsync[1], !prev_cnt[1], prev_cnt[12], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12865(w_eco12865, Tsync[1], prev_cnt[9], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12866(w_eco12866, prev_cnt[1], prev_cnt[6], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12867(w_eco12867, prev_cnt[1], prev_cnt[10], !prev_cnt[15], prev_state[1]);
	and _ECO_12868(w_eco12868, !prev_cnt[14], prev_cnt[1], prev_cnt[12], !prev_cnt[15], prev_state[1]);
	and _ECO_12869(w_eco12869, !prev_cnt[1], prev_cnt[9], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12870(w_eco12870, Tsync[1], prev_cnt[9], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12871(w_eco12871, prev_cnt[1], prev_cnt[8], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12872(w_eco12872, !prev_cnt[1], prev_cnt[13], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12873(w_eco12873, Tsync[1], prev_cnt[6], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12874(w_eco12874, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12875(w_eco12875, !prev_cnt[14], prev_cnt[13], !prev_cnt[15], !ena);
	and _ECO_12876(w_eco12876, Tsync[1], prev_cnt[1], prev_cnt[8], !prev_cnt[15], prev_state[0]);
	and _ECO_12877(w_eco12877, prev_cnt[9], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12878(w_eco12878, !Tsync[1], prev_cnt[9], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12879(w_eco12879, !prev_cnt[1], prev_cnt[13], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12880(w_eco12880, !Tsync[1], !prev_cnt[1], prev_cnt[9], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12881(w_eco12881, !Tsync[1], prev_cnt[9], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12882(w_eco12882, prev_cnt[9], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12883(w_eco12883, !Tsync[1], !prev_cnt[1], prev_cnt[13], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12884(w_eco12884, Tsync[1], prev_cnt[6], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12885(w_eco12885, prev_cnt[1], prev_cnt[8], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12886(w_eco12886, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[1]);
	and _ECO_12887(w_eco12887, !prev_cnt[14], prev_cnt[1], prev_cnt[13], !prev_cnt[15], prev_state[1]);
	and _ECO_12888(w_eco12888, !prev_cnt[1], prev_cnt[6], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12889(w_eco12889, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_12890(w_eco12890, !prev_cnt[1], prev_cnt[8], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12891(w_eco12891, Tsync[1], prev_cnt[6], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12892(w_eco12892, prev_cnt[1], prev_cnt[10], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12893(w_eco12893, !prev_cnt[1], prev_cnt[9], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12894(w_eco12894, Tsync[1], prev_cnt[8], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12895(w_eco12895, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12896(w_eco12896, Tsync[1], prev_cnt[1], prev_cnt[10], !prev_cnt[15], prev_state[0]);
	and _ECO_12897(w_eco12897, Tsync[1], !prev_cnt[14], prev_cnt[1], prev_cnt[12], !prev_cnt[15], prev_state[0]);
	and _ECO_12898(w_eco12898, prev_cnt[6], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12899(w_eco12899, Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12900(w_eco12900, !Tsync[1], prev_cnt[6], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12901(w_eco12901, !Tsync[1], Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12902(w_eco12902, !Tsync[1], prev_cnt[8], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12903(w_eco12903, !prev_cnt[1], prev_cnt[9], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12904(w_eco12904, !Tsync[1], !prev_cnt[1], prev_cnt[6], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12905(w_eco12905, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_12906(w_eco12906, !Tsync[1], !prev_cnt[1], prev_cnt[8], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12907(w_eco12907, !Tsync[1], prev_cnt[6], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12908(w_eco12908, !Tsync[1], Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12909(w_eco12909, !Tsync[1], prev_cnt[8], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12910(w_eco12910, prev_cnt[6], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12911(w_eco12911, Tgate[15], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12912(w_eco12912, !Tsync[1], !prev_cnt[1], prev_cnt[9], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12913(w_eco12913, Tsync[1], prev_cnt[8], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12914(w_eco12914, prev_cnt[1], prev_cnt[10], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12915(w_eco12915, !prev_cnt[14], prev_cnt[1], prev_cnt[12], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12916(w_eco12916, !prev_cnt[1], prev_cnt[10], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_12917(w_eco12917, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_12918(w_eco12918, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_12919(w_eco12919, Tsync[1], prev_cnt[8], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12920(w_eco12920, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12921(w_eco12921, !prev_cnt[14], prev_cnt[1], prev_cnt[13], !prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_12922(w_eco12922, !prev_cnt[1], prev_cnt[6], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12923(w_eco12923, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12924(w_eco12924, !prev_cnt[1], prev_cnt[8], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12925(w_eco12925, Tsync[1], prev_cnt[10], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12926(w_eco12926, Tsync[1], !prev_cnt[14], prev_cnt[12], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12927(w_eco12927, Tsync[1], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[0]);
	and _ECO_12928(w_eco12928, Tsync[1], !prev_cnt[14], prev_cnt[1], prev_cnt[13], !prev_cnt[15], prev_state[0]);
	and _ECO_12929(w_eco12929, prev_cnt[8], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12930(w_eco12930, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_12931(w_eco12931, !prev_cnt[1], prev_cnt[6], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12932(w_eco12932, !Tsync[1], prev_cnt[10], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_12933(w_eco12933, !Tsync[1], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12934(w_eco12934, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_12935(w_eco12935, !Tsync[1], !prev_cnt[1], prev_cnt[6], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12936(w_eco12936, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_12937(w_eco12937, !prev_cnt[1], prev_cnt[8], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12938(w_eco12938, !Tsync[1], !prev_cnt[1], prev_cnt[10], prev_cnt[15], ena, prev_state[1]);
	and _ECO_12939(w_eco12939, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2]);
	and _ECO_12940(w_eco12940, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_12941(w_eco12941, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12942(w_eco12942, !Tsync[1], prev_cnt[10], prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12943(w_eco12943, !Tsync[1], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_12944(w_eco12944, prev_cnt[8], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12945(w_eco12945, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_12946(w_eco12946, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_12947(w_eco12947, !Tsync[1], !prev_cnt[1], prev_cnt[8], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12948(w_eco12948, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_12949(w_eco12949, Tsync[1], prev_cnt[10], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12950(w_eco12950, Tsync[1], !prev_cnt[14], prev_cnt[12], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12951(w_eco12951, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12952(w_eco12952, !prev_cnt[14], prev_cnt[1], prev_cnt[13], !prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_12953(w_eco12953, Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_12954(w_eco12954, Tsync[1], prev_cnt[10], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12955(w_eco12955, Tsync[1], !prev_cnt[14], prev_cnt[12], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12956(w_eco12956, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12957(w_eco12957, !prev_cnt[1], prev_cnt[10], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12958(w_eco12958, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12959(w_eco12959, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_12960(w_eco12960, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12961(w_eco12961, Tsync[1], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12962(w_eco12962, Tsync[1], !prev_cnt[14], prev_cnt[13], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12963(w_eco12963, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_12964(w_eco12964, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12965(w_eco12965, prev_cnt[10], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12966(w_eco12966, Tgate[15], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12967(w_eco12967, prev_cnt[10], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12968(w_eco12968, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_12969(w_eco12969, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_12970(w_eco12970, !prev_cnt[1], prev_cnt[10], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_12971(w_eco12971, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_12972(w_eco12972, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_12973(w_eco12973, !Tsync[1], Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_12974(w_eco12974, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_12975(w_eco12975, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_12976(w_eco12976, !Tsync[1], !prev_cnt[1], prev_cnt[10], prev_cnt[15], ena, prev_state[0]);
	and _ECO_12977(w_eco12977, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_12978(w_eco12978, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12979(w_eco12979, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_12980(w_eco12980, Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_12981(w_eco12981, !Tsync[1], Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_12982(w_eco12982, Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_12983(w_eco12983, !Tsync[1], Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena);
	and _ECO_12984(w_eco12984, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_12985(w_eco12985, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_12986(w_eco12986, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_12987(w_eco12987, Tsync[1], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12988(w_eco12988, Tsync[1], !prev_cnt[14], prev_cnt[13], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_12989(w_eco12989, Tsync[1], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12990(w_eco12990, Tsync[1], !prev_cnt[14], prev_cnt[13], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_12991(w_eco12991, Tsync[1], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_12992(w_eco12992, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_12993(w_eco12993, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12994(w_eco12994, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !prev_cnt[15], !ena);
	and _ECO_12995(w_eco12995, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_12996(w_eco12996, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_12997(w_eco12997, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_12998(w_eco12998, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_12999(w_eco12999, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_13000(w_eco13000, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_13001(w_eco13001, !Tsync[1], Tgate[15], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena);
	and _ECO_13002(w_eco13002, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_13003(w_eco13003, !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_13004(w_eco13004, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13005(w_eco13005, Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_13006(w_eco13006, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13007(w_eco13007, Tgate[15], prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13008(w_eco13008, Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_13009(w_eco13009, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_13010(w_eco13010, !Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_13011(w_eco13011, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena);
	and _ECO_13012(w_eco13012, Tgate[15], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_13013(w_eco13013, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_13014(w_eco13014, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_13015(w_eco13015, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_13016(w_eco13016, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_13017(w_eco13017, !Tsync[1], Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena);
	and _ECO_13018(w_eco13018, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1]);
	and _ECO_13019(w_eco13019, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_13020(w_eco13020, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_13021(w_eco13021, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13022(w_eco13022, Tgate[15], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_13023(w_eco13023, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_13024(w_eco13024, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_13025(w_eco13025, Tsync[1], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13026(w_eco13026, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_13027(w_eco13027, Tsync[1], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13028(w_eco13028, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13029(w_eco13029, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2]);
	and _ECO_13030(w_eco13030, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13031(w_eco13031, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13032(w_eco13032, Tsync[1], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_13033(w_eco13033, Tsync[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_13034(w_eco13034, Tsync[1], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_13035(w_eco13035, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_13036(w_eco13036, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_13037(w_eco13037, !Tsync[1], !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_13038(w_eco13038, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_13039(w_eco13039, Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_13040(w_eco13040, !Tsync[1], Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[0]);
	and _ECO_13041(w_eco13041, Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[1], !prev_state[0]);
	and _ECO_13042(w_eco13042, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_13043(w_eco13043, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_13044(w_eco13044, !Tsync[1], !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2]);
	and _ECO_13045(w_eco13045, !Tsync[1], !prev_cnt[14], !prev_cnt[0], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], ena, prev_state[1]);
	and _ECO_13046(w_eco13046, Tgate[15], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_13047(w_eco13047, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_13048(w_eco13048, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_13049(w_eco13049, Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13050(w_eco13050, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_13051(w_eco13051, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_13052(w_eco13052, Tsync[1], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13053(w_eco13053, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13054(w_eco13054, Tgate[15], !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2]);
	and _ECO_13055(w_eco13055, Tgate[15], prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13056(w_eco13056, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13057(w_eco13057, Tsync[1], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[3], prev_state[0]);
	and _ECO_13058(w_eco13058, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_13059(w_eco13059, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_13060(w_eco13060, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13061(w_eco13061, !Tsync[1], !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[0]);
	and _ECO_13062(w_eco13062, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_13063(w_eco13063, !Tsync[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[0]);
	and _ECO_13064(w_eco13064, Tgate[15], !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[0]);
	and _ECO_13065(w_eco13065, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[0]);
	and _ECO_13066(w_eco13066, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13067(w_eco13067, Tgate[15], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_13068(w_eco13068, Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[3], prev_state[1]);
	and _ECO_13069(w_eco13069, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_13070(w_eco13070, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_13071(w_eco13071, Tsync[1], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13072(w_eco13072, Tsync[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13073(w_eco13073, Tsync[1], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13074(w_eco13074, Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_13075(w_eco13075, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_13076(w_eco13076, Tsync[1], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13077(w_eco13077, Tsync[1], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], !prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13078(w_eco13078, Tsync[1], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13079(w_eco13079, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13080(w_eco13080, Tgate[15], !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2]);
	and _ECO_13081(w_eco13081, Tgate[15], prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13082(w_eco13082, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13083(w_eco13083, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13084(w_eco13084, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[0]);
	and _ECO_13085(w_eco13085, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13086(w_eco13086, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13087(w_eco13087, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13088(w_eco13088, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13089(w_eco13089, !prev_cnt[14], !prev_cnt[0], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], ena, prev_state[1], !prev_state[0]);
	and _ECO_13090(w_eco13090, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13091(w_eco13091, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[3], prev_state[1], prev_state[0]);
	and _ECO_13092(w_eco13092, !prev_cnt[14], !prev_cnt[0], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], ena, !prev_state[3], prev_state[1]);
	and _ECO_13093(w_eco13093, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_13094(w_eco13094, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13095(w_eco13095, Tsync[1], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13096(w_eco13096, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[0]);
	and _ECO_13097(w_eco13097, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13098(w_eco13098, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_13099(w_eco13099, Tsync[1], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], prev_state[4], !prev_state[1], prev_state[0]);
	and _ECO_13100(w_eco13100, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[1], !prev_state[0]);
	and _ECO_13101(w_eco13101, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13102(w_eco13102, !prev_cnt[14], !prev_cnt[0], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[6], !prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], ena, !prev_state[4], !prev_state[3], !prev_state[2], prev_state[0]);
	and _ECO_13103(w_eco13103, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13104(w_eco13104, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13105(w_eco13105, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13106(w_eco13106, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13107(w_eco13107, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13108(w_eco13108, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[3], !prev_state[2], !prev_state[0]);
	and _ECO_13109(w_eco13109, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[0]);
	and _ECO_13110(w_eco13110, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13111(w_eco13111, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13112(w_eco13112, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13113(w_eco13113, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13114(w_eco13114, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13115(w_eco13115, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13116(w_eco13116, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13117(w_eco13117, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13118(w_eco13118, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13119(w_eco13119, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13120(w_eco13120, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13121(w_eco13121, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13122(w_eco13122, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13123(w_eco13123, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13124(w_eco13124, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13125(w_eco13125, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13126(w_eco13126, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13127(w_eco13127, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13128(w_eco13128, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13129(w_eco13129, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13130(w_eco13130, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13131(w_eco13131, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13132(w_eco13132, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13133(w_eco13133, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13134(w_eco13134, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13135(w_eco13135, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13136(w_eco13136, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13137(w_eco13137, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13138(w_eco13138, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13139(w_eco13139, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13140(w_eco13140, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13141(w_eco13141, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13142(w_eco13142, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13143(w_eco13143, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13144(w_eco13144, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13145(w_eco13145, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13146(w_eco13146, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13147(w_eco13147, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13148(w_eco13148, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13149(w_eco13149, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13150(w_eco13150, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13151(w_eco13151, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13152(w_eco13152, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13153(w_eco13153, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13154(w_eco13154, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13155(w_eco13155, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13156(w_eco13156, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13157(w_eco13157, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13158(w_eco13158, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13159(w_eco13159, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13160(w_eco13160, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13161(w_eco13161, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13162(w_eco13162, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13163(w_eco13163, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13164(w_eco13164, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13165(w_eco13165, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13166(w_eco13166, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13167(w_eco13167, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13168(w_eco13168, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13169(w_eco13169, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13170(w_eco13170, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13171(w_eco13171, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13172(w_eco13172, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13173(w_eco13173, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13174(w_eco13174, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13175(w_eco13175, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13176(w_eco13176, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13177(w_eco13177, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13178(w_eco13178, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13179(w_eco13179, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13180(w_eco13180, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13181(w_eco13181, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13182(w_eco13182, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13183(w_eco13183, !prev_cnt[14], !prev_cnt[1], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13184(w_eco13184, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13185(w_eco13185, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13186(w_eco13186, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13187(w_eco13187, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13188(w_eco13188, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13189(w_eco13189, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13190(w_eco13190, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13191(w_eco13191, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13192(w_eco13192, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13193(w_eco13193, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13194(w_eco13194, !prev_cnt[14], !prev_cnt[1], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13195(w_eco13195, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13196(w_eco13196, !Tgate[15], prev_cnt[1], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13197(w_eco13197, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13198(w_eco13198, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13199(w_eco13199, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13200(w_eco13200, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13201(w_eco13201, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13202(w_eco13202, !prev_cnt[14], prev_cnt[0], !prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13203(w_eco13203, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13204(w_eco13204, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13205(w_eco13205, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13206(w_eco13206, !prev_cnt[14], !prev_cnt[1], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13207(w_eco13207, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13208(w_eco13208, !prev_cnt[14], !prev_cnt[1], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13209(w_eco13209, !prev_cnt[14], !prev_cnt[1], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, prev_state[1], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_13210(w_eco13210, w_eco12797, w_eco12798, w_eco12799, w_eco12800, w_eco12801, w_eco12802, w_eco12803, w_eco12804, w_eco12805, w_eco12806, w_eco12807, w_eco12808, w_eco12809, w_eco12810, w_eco12811, w_eco12812, w_eco12813, w_eco12814, w_eco12815, w_eco12816, w_eco12817, w_eco12818, w_eco12819, w_eco12820, w_eco12821, w_eco12822, w_eco12823, w_eco12824, w_eco12825, w_eco12826, w_eco12827, w_eco12828, w_eco12829, w_eco12830, w_eco12831, w_eco12832, w_eco12833, w_eco12834, w_eco12835, w_eco12836, w_eco12837, w_eco12838, w_eco12839, w_eco12840, w_eco12841, w_eco12842, w_eco12843, w_eco12844, w_eco12845, w_eco12846, w_eco12847, w_eco12848, w_eco12849, w_eco12850, w_eco12851, w_eco12852, w_eco12853, w_eco12854, w_eco12855, w_eco12856, w_eco12857, w_eco12858, w_eco12859, w_eco12860, w_eco12861, w_eco12862, w_eco12863, w_eco12864, w_eco12865, w_eco12866, w_eco12867, w_eco12868, w_eco12869, w_eco12870, w_eco12871, w_eco12872, w_eco12873, w_eco12874, w_eco12875, w_eco12876, w_eco12877, w_eco12878, w_eco12879, w_eco12880, w_eco12881, w_eco12882, w_eco12883, w_eco12884, w_eco12885, w_eco12886, w_eco12887, w_eco12888, w_eco12889, w_eco12890, w_eco12891, w_eco12892, w_eco12893, w_eco12894, w_eco12895, w_eco12896, w_eco12897, w_eco12898, w_eco12899, w_eco12900, w_eco12901, w_eco12902, w_eco12903, w_eco12904, w_eco12905, w_eco12906, w_eco12907, w_eco12908, w_eco12909, w_eco12910, w_eco12911, w_eco12912, w_eco12913, w_eco12914, w_eco12915, w_eco12916, w_eco12917, w_eco12918, w_eco12919, w_eco12920, w_eco12921, w_eco12922, w_eco12923, w_eco12924, w_eco12925, w_eco12926, w_eco12927, w_eco12928, w_eco12929, w_eco12930, w_eco12931, w_eco12932, w_eco12933, w_eco12934, w_eco12935, w_eco12936, w_eco12937, w_eco12938, w_eco12939, w_eco12940, w_eco12941, w_eco12942, w_eco12943, w_eco12944, w_eco12945, w_eco12946, w_eco12947, w_eco12948, w_eco12949, w_eco12950, w_eco12951, w_eco12952, w_eco12953, w_eco12954, w_eco12955, w_eco12956, w_eco12957, w_eco12958, w_eco12959, w_eco12960, w_eco12961, w_eco12962, w_eco12963, w_eco12964, w_eco12965, w_eco12966, w_eco12967, w_eco12968, w_eco12969, w_eco12970, w_eco12971, w_eco12972, w_eco12973, w_eco12974, w_eco12975, w_eco12976, w_eco12977, w_eco12978, w_eco12979, w_eco12980, w_eco12981, w_eco12982, w_eco12983, w_eco12984, w_eco12985, w_eco12986, w_eco12987, w_eco12988, w_eco12989, w_eco12990, w_eco12991, w_eco12992, w_eco12993, w_eco12994, w_eco12995, w_eco12996, w_eco12997, w_eco12998, w_eco12999, w_eco13000, w_eco13001, w_eco13002, w_eco13003, w_eco13004, w_eco13005, w_eco13006, w_eco13007, w_eco13008, w_eco13009, w_eco13010, w_eco13011, w_eco13012, w_eco13013, w_eco13014, w_eco13015, w_eco13016, w_eco13017, w_eco13018, w_eco13019, w_eco13020, w_eco13021, w_eco13022, w_eco13023, w_eco13024, w_eco13025, w_eco13026, w_eco13027, w_eco13028, w_eco13029, w_eco13030, w_eco13031, w_eco13032, w_eco13033, w_eco13034, w_eco13035, w_eco13036, w_eco13037, w_eco13038, w_eco13039, w_eco13040, w_eco13041, w_eco13042, w_eco13043, w_eco13044, w_eco13045, w_eco13046, w_eco13047, w_eco13048, w_eco13049, w_eco13050, w_eco13051, w_eco13052, w_eco13053, w_eco13054, w_eco13055, w_eco13056, w_eco13057, w_eco13058, w_eco13059, w_eco13060, w_eco13061, w_eco13062, w_eco13063, w_eco13064, w_eco13065, w_eco13066, w_eco13067, w_eco13068, w_eco13069, w_eco13070, w_eco13071, w_eco13072, w_eco13073, w_eco13074, w_eco13075, w_eco13076, w_eco13077, w_eco13078, w_eco13079, w_eco13080, w_eco13081, w_eco13082, w_eco13083, w_eco13084, w_eco13085, w_eco13086, w_eco13087, w_eco13088, w_eco13089, w_eco13090, w_eco13091, w_eco13092, w_eco13093, w_eco13094, w_eco13095, w_eco13096, w_eco13097, w_eco13098, w_eco13099, w_eco13100, w_eco13101, w_eco13102, w_eco13103, w_eco13104, w_eco13105, w_eco13106, w_eco13107, w_eco13108, w_eco13109, w_eco13110, w_eco13111, w_eco13112, w_eco13113, w_eco13114, w_eco13115, w_eco13116, w_eco13117, w_eco13118, w_eco13119, w_eco13120, w_eco13121, w_eco13122, w_eco13123, w_eco13124, w_eco13125, w_eco13126, w_eco13127, w_eco13128, w_eco13129, w_eco13130, w_eco13131, w_eco13132, w_eco13133, w_eco13134, w_eco13135, w_eco13136, w_eco13137, w_eco13138, w_eco13139, w_eco13140, w_eco13141, w_eco13142, w_eco13143, w_eco13144, w_eco13145, w_eco13146, w_eco13147, w_eco13148, w_eco13149, w_eco13150, w_eco13151, w_eco13152, w_eco13153, w_eco13154, w_eco13155, w_eco13156, w_eco13157, w_eco13158, w_eco13159, w_eco13160, w_eco13161, w_eco13162, w_eco13163, w_eco13164, w_eco13165, w_eco13166, w_eco13167, w_eco13168, w_eco13169, w_eco13170, w_eco13171, w_eco13172, w_eco13173, w_eco13174, w_eco13175, w_eco13176, w_eco13177, w_eco13178, w_eco13179, w_eco13180, w_eco13181, w_eco13182, w_eco13183, w_eco13184, w_eco13185, w_eco13186, w_eco13187, w_eco13188, w_eco13189, w_eco13190, w_eco13191, w_eco13192, w_eco13193, w_eco13194, w_eco13195, w_eco13196, w_eco13197, w_eco13198, w_eco13199, w_eco13200, w_eco13201, w_eco13202, w_eco13203, w_eco13204, w_eco13205, w_eco13206, w_eco13207, w_eco13208, w_eco13209);
	xor _ECO_out10(cnt[15], sub_wire10, w_eco13210);
	and _ECO_13211(w_eco13211, prev_cnt[14], rst);
	and _ECO_13212(w_eco13212, prev_cnt[14], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13213(w_eco13213, prev_cnt[14], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13214(w_eco13214, prev_cnt[14], prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13215(w_eco13215, prev_cnt[14], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13216(w_eco13216, prev_cnt[14], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13217(w_eco13217, prev_cnt[14], prev_cnt[12], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13218(w_eco13218, prev_cnt[14], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13219(w_eco13219, Tgate[14], prev_cnt[14], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13220(w_eco13220, prev_cnt[14], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13221(w_eco13221, Tgate[14], prev_cnt[14], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13222(w_eco13222, prev_cnt[14], prev_cnt[12], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13223(w_eco13223, prev_cnt[14], prev_cnt[13], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13224(w_eco13224, prev_cnt[14], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13225(w_eco13225, prev_cnt[14], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13226(w_eco13226, prev_cnt[14], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13227(w_eco13227, prev_cnt[14], prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13228(w_eco13228, prev_cnt[14], prev_cnt[6], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13229(w_eco13229, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13230(w_eco13230, prev_cnt[14], prev_cnt[9], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13231(w_eco13231, prev_cnt[14], prev_cnt[6], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13232(w_eco13232, prev_cnt[14], prev_cnt[6], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13233(w_eco13233, prev_cnt[14], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13234(w_eco13234, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13235(w_eco13235, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13236(w_eco13236, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13237(w_eco13237, prev_cnt[14], prev_cnt[6], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13238(w_eco13238, prev_cnt[14], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13239(w_eco13239, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13240(w_eco13240, prev_cnt[14], prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13241(w_eco13241, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13242(w_eco13242, prev_cnt[14], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13243(w_eco13243, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13244(w_eco13244, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13245(w_eco13245, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13246(w_eco13246, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13247(w_eco13247, prev_cnt[14], prev_cnt[8], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13248(w_eco13248, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13249(w_eco13249, prev_cnt[14], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13250(w_eco13250, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13251(w_eco13251, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13252(w_eco13252, prev_cnt[14], prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13253(w_eco13253, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13254(w_eco13254, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13255(w_eco13255, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13256(w_eco13256, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13257(w_eco13257, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13258(w_eco13258, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13259(w_eco13259, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13260(w_eco13260, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13261(w_eco13261, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13262(w_eco13262, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13263(w_eco13263, prev_cnt[14], prev_cnt[10], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13264(w_eco13264, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13265(w_eco13265, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13266(w_eco13266, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13267(w_eco13267, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13268(w_eco13268, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13269(w_eco13269, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13270(w_eco13270, prev_cnt[14], prev_cnt[13], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13271(w_eco13271, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13272(w_eco13272, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13273(w_eco13273, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13274(w_eco13274, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13275(w_eco13275, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13276(w_eco13276, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13277(w_eco13277, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13278(w_eco13278, Tgate[14], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13279(w_eco13279, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13280(w_eco13280, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13281(w_eco13281, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13282(w_eco13282, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13283(w_eco13283, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13284(w_eco13284, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13285(w_eco13285, Tgate[14], prev_cnt[14], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13286(w_eco13286, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13287(w_eco13287, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13288(w_eco13288, prev_cnt[14], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13289(w_eco13289, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13290(w_eco13290, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13291(w_eco13291, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13292(w_eco13292, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13293(w_eco13293, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13294(w_eco13294, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13295(w_eco13295, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13296(w_eco13296, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13297(w_eco13297, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13298(w_eco13298, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13299(w_eco13299, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13300(w_eco13300, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13301(w_eco13301, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13302(w_eco13302, Tgate[14], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13303(w_eco13303, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13304(w_eco13304, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13305(w_eco13305, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13306(w_eco13306, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13307(w_eco13307, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13308(w_eco13308, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13309(w_eco13309, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13310(w_eco13310, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13311(w_eco13311, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13312(w_eco13312, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13313(w_eco13313, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13314(w_eco13314, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13315(w_eco13315, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13316(w_eco13316, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13317(w_eco13317, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13318(w_eco13318, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13319(w_eco13319, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13320(w_eco13320, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13321(w_eco13321, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13322(w_eco13322, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13323(w_eco13323, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13324(w_eco13324, Tgate[14], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13325(w_eco13325, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13326(w_eco13326, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13327(w_eco13327, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13328(w_eco13328, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13329(w_eco13329, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13330(w_eco13330, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13331(w_eco13331, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13332(w_eco13332, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13333(w_eco13333, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13334(w_eco13334, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13335(w_eco13335, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13336(w_eco13336, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13337(w_eco13337, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13338(w_eco13338, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13339(w_eco13339, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13340(w_eco13340, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13341(w_eco13341, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13342(w_eco13342, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13343(w_eco13343, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13344(w_eco13344, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13345(w_eco13345, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13346(w_eco13346, Tgate[14], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13347(w_eco13347, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13348(w_eco13348, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13349(w_eco13349, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !ena, !rst);
	and _ECO_13350(w_eco13350, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13351(w_eco13351, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], !prev_state[2]);
	and _ECO_13352(w_eco13352, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13353(w_eco13353, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13354(w_eco13354, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13355(w_eco13355, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[3], !prev_state[2]);
	and _ECO_13356(w_eco13356, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13357(w_eco13357, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13358(w_eco13358, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13359(w_eco13359, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13360(w_eco13360, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13361(w_eco13361, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13362(w_eco13362, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13363(w_eco13363, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13364(w_eco13364, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13365(w_eco13365, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13366(w_eco13366, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13367(w_eco13367, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena, !rst);
	and _ECO_13368(w_eco13368, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13369(w_eco13369, Tgate[14], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13370(w_eco13370, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13371(w_eco13371, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13372(w_eco13372, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13373(w_eco13373, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_state[1]);
	and _ECO_13374(w_eco13374, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13375(w_eco13375, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13376(w_eco13376, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13377(w_eco13377, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13378(w_eco13378, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13379(w_eco13379, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13380(w_eco13380, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13381(w_eco13381, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13382(w_eco13382, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13383(w_eco13383, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13384(w_eco13384, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13385(w_eco13385, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13386(w_eco13386, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], ena, !rst, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13387(w_eco13387, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13388(w_eco13388, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13389(w_eco13389, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13390(w_eco13390, Tgate[14], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13391(w_eco13391, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13392(w_eco13392, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !ena);
	and _ECO_13393(w_eco13393, prev_cnt[14], !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13394(w_eco13394, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13395(w_eco13395, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13396(w_eco13396, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13397(w_eco13397, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13398(w_eco13398, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13399(w_eco13399, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13400(w_eco13400, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13401(w_eco13401, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13402(w_eco13402, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13403(w_eco13403, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13404(w_eco13404, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13405(w_eco13405, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13406(w_eco13406, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13407(w_eco13407, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13408(w_eco13408, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13409(w_eco13409, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13410(w_eco13410, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13411(w_eco13411, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13412(w_eco13412, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13413(w_eco13413, Tgate[14], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13414(w_eco13414, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13415(w_eco13415, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13416(w_eco13416, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13417(w_eco13417, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13418(w_eco13418, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13419(w_eco13419, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13420(w_eco13420, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13421(w_eco13421, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13422(w_eco13422, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13423(w_eco13423, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13424(w_eco13424, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13425(w_eco13425, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13426(w_eco13426, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13427(w_eco13427, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13428(w_eco13428, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13429(w_eco13429, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13430(w_eco13430, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13431(w_eco13431, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13432(w_eco13432, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13433(w_eco13433, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13434(w_eco13434, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13435(w_eco13435, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13436(w_eco13436, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13437(w_eco13437, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13438(w_eco13438, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13439(w_eco13439, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13440(w_eco13440, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13441(w_eco13441, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13442(w_eco13442, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13443(w_eco13443, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13444(w_eco13444, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13445(w_eco13445, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13446(w_eco13446, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13447(w_eco13447, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13448(w_eco13448, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13449(w_eco13449, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13450(w_eco13450, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13451(w_eco13451, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13452(w_eco13452, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13453(w_eco13453, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13454(w_eco13454, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13455(w_eco13455, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13456(w_eco13456, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13457(w_eco13457, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13458(w_eco13458, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13459(w_eco13459, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13460(w_eco13460, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13461(w_eco13461, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13462(w_eco13462, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13463(w_eco13463, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13464(w_eco13464, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13465(w_eco13465, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13466(w_eco13466, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13467(w_eco13467, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13468(w_eco13468, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13469(w_eco13469, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13470(w_eco13470, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13471(w_eco13471, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13472(w_eco13472, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13473(w_eco13473, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13474(w_eco13474, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13475(w_eco13475, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13476(w_eco13476, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13477(w_eco13477, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13478(w_eco13478, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13479(w_eco13479, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13480(w_eco13480, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13481(w_eco13481, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13482(w_eco13482, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13483(w_eco13483, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13484(w_eco13484, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13485(w_eco13485, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13486(w_eco13486, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13487(w_eco13487, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13488(w_eco13488, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13489(w_eco13489, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13490(w_eco13490, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13491(w_eco13491, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13492(w_eco13492, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13493(w_eco13493, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13494(w_eco13494, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13495(w_eco13495, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13496(w_eco13496, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13497(w_eco13497, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13498(w_eco13498, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13499(w_eco13499, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13500(w_eco13500, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13501(w_eco13501, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13502(w_eco13502, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13503(w_eco13503, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13504(w_eco13504, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13505(w_eco13505, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13506(w_eco13506, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13507(w_eco13507, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13508(w_eco13508, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13509(w_eco13509, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13510(w_eco13510, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13511(w_eco13511, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13512(w_eco13512, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13513(w_eco13513, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13514(w_eco13514, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13515(w_eco13515, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13516(w_eco13516, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13517(w_eco13517, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13518(w_eco13518, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13519(w_eco13519, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13520(w_eco13520, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13521(w_eco13521, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13522(w_eco13522, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13523(w_eco13523, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13524(w_eco13524, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13525(w_eco13525, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13526(w_eco13526, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13527(w_eco13527, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13528(w_eco13528, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13529(w_eco13529, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13530(w_eco13530, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13531(w_eco13531, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13532(w_eco13532, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13533(w_eco13533, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13534(w_eco13534, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13535(w_eco13535, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13536(w_eco13536, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13537(w_eco13537, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13538(w_eco13538, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13539(w_eco13539, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13540(w_eco13540, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13541(w_eco13541, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13542(w_eco13542, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13543(w_eco13543, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13544(w_eco13544, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13545(w_eco13545, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13546(w_eco13546, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13547(w_eco13547, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13548(w_eco13548, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13549(w_eco13549, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13550(w_eco13550, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13551(w_eco13551, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13552(w_eco13552, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13553(w_eco13553, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13554(w_eco13554, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13555(w_eco13555, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13556(w_eco13556, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13557(w_eco13557, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13558(w_eco13558, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13559(w_eco13559, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13560(w_eco13560, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13561(w_eco13561, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13562(w_eco13562, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13563(w_eco13563, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13564(w_eco13564, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13565(w_eco13565, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13566(w_eco13566, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13567(w_eco13567, !Tgate[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13568(w_eco13568, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13569(w_eco13569, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13570(w_eco13570, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13571(w_eco13571, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13572(w_eco13572, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13573(w_eco13573, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13574(w_eco13574, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13575(w_eco13575, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13576(w_eco13576, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13577(w_eco13577, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13578(w_eco13578, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13579(w_eco13579, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13580(w_eco13580, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13581(w_eco13581, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13582(w_eco13582, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13583(w_eco13583, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13584(w_eco13584, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13585(w_eco13585, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13586(w_eco13586, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13587(w_eco13587, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13588(w_eco13588, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13589(w_eco13589, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13590(w_eco13590, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13591(w_eco13591, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13592(w_eco13592, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13593(w_eco13593, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13594(w_eco13594, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13595(w_eco13595, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13596(w_eco13596, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13597(w_eco13597, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13598(w_eco13598, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13599(w_eco13599, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13600(w_eco13600, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13601(w_eco13601, !Tgate[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13602(w_eco13602, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13603(w_eco13603, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13604(w_eco13604, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13605(w_eco13605, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13606(w_eco13606, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13607(w_eco13607, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13608(w_eco13608, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13609(w_eco13609, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13610(w_eco13610, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13611(w_eco13611, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13612(w_eco13612, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13613(w_eco13613, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13614(w_eco13614, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13615(w_eco13615, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13616(w_eco13616, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13617(w_eco13617, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13618(w_eco13618, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13619(w_eco13619, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13620(w_eco13620, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13621(w_eco13621, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13622(w_eco13622, !Tgate[14], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13623(w_eco13623, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13624(w_eco13624, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13625(w_eco13625, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13626(w_eco13626, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13627(w_eco13627, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13628(w_eco13628, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13629(w_eco13629, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13630(w_eco13630, !Tgate[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13631(w_eco13631, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13632(w_eco13632, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13633(w_eco13633, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13634(w_eco13634, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13635(w_eco13635, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13636(w_eco13636, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13637(w_eco13637, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13638(w_eco13638, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13639(w_eco13639, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13640(w_eco13640, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13641(w_eco13641, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13642(w_eco13642, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13643(w_eco13643, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13644(w_eco13644, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13645(w_eco13645, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13646(w_eco13646, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13647(w_eco13647, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13648(w_eco13648, !Tgate[14], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13649(w_eco13649, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13650(w_eco13650, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13651(w_eco13651, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13652(w_eco13652, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13653(w_eco13653, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13654(w_eco13654, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13655(w_eco13655, !Tgate[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13656(w_eco13656, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13657(w_eco13657, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13658(w_eco13658, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13659(w_eco13659, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13660(w_eco13660, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13661(w_eco13661, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13662(w_eco13662, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13663(w_eco13663, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13664(w_eco13664, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13665(w_eco13665, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13666(w_eco13666, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13667(w_eco13667, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13668(w_eco13668, !Tgate[14], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13669(w_eco13669, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13670(w_eco13670, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13671(w_eco13671, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13672(w_eco13672, !Tgate[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13673(w_eco13673, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13674(w_eco13674, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13675(w_eco13675, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13676(w_eco13676, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13677(w_eco13677, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13678(w_eco13678, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13679(w_eco13679, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13680(w_eco13680, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13681(w_eco13681, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13682(w_eco13682, !Tgate[14], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13683(w_eco13683, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13684(w_eco13684, !Tgate[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13685(w_eco13685, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13686(w_eco13686, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13687(w_eco13687, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13688(w_eco13688, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13689(w_eco13689, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13690(w_eco13690, !Tgate[14], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13691(w_eco13691, !Tgate[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13692(w_eco13692, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13693(w_eco13693, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13694(w_eco13694, !Tgate[14], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13695(w_eco13695, !Tgate[14], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_13696(w_eco13696, w_eco13211, w_eco13212, w_eco13213, w_eco13214, w_eco13215, w_eco13216, w_eco13217, w_eco13218, w_eco13219, w_eco13220, w_eco13221, w_eco13222, w_eco13223, w_eco13224, w_eco13225, w_eco13226, w_eco13227, w_eco13228, w_eco13229, w_eco13230, w_eco13231, w_eco13232, w_eco13233, w_eco13234, w_eco13235, w_eco13236, w_eco13237, w_eco13238, w_eco13239, w_eco13240, w_eco13241, w_eco13242, w_eco13243, w_eco13244, w_eco13245, w_eco13246, w_eco13247, w_eco13248, w_eco13249, w_eco13250, w_eco13251, w_eco13252, w_eco13253, w_eco13254, w_eco13255, w_eco13256, w_eco13257, w_eco13258, w_eco13259, w_eco13260, w_eco13261, w_eco13262, w_eco13263, w_eco13264, w_eco13265, w_eco13266, w_eco13267, w_eco13268, w_eco13269, w_eco13270, w_eco13271, w_eco13272, w_eco13273, w_eco13274, w_eco13275, w_eco13276, w_eco13277, w_eco13278, w_eco13279, w_eco13280, w_eco13281, w_eco13282, w_eco13283, w_eco13284, w_eco13285, w_eco13286, w_eco13287, w_eco13288, w_eco13289, w_eco13290, w_eco13291, w_eco13292, w_eco13293, w_eco13294, w_eco13295, w_eco13296, w_eco13297, w_eco13298, w_eco13299, w_eco13300, w_eco13301, w_eco13302, w_eco13303, w_eco13304, w_eco13305, w_eco13306, w_eco13307, w_eco13308, w_eco13309, w_eco13310, w_eco13311, w_eco13312, w_eco13313, w_eco13314, w_eco13315, w_eco13316, w_eco13317, w_eco13318, w_eco13319, w_eco13320, w_eco13321, w_eco13322, w_eco13323, w_eco13324, w_eco13325, w_eco13326, w_eco13327, w_eco13328, w_eco13329, w_eco13330, w_eco13331, w_eco13332, w_eco13333, w_eco13334, w_eco13335, w_eco13336, w_eco13337, w_eco13338, w_eco13339, w_eco13340, w_eco13341, w_eco13342, w_eco13343, w_eco13344, w_eco13345, w_eco13346, w_eco13347, w_eco13348, w_eco13349, w_eco13350, w_eco13351, w_eco13352, w_eco13353, w_eco13354, w_eco13355, w_eco13356, w_eco13357, w_eco13358, w_eco13359, w_eco13360, w_eco13361, w_eco13362, w_eco13363, w_eco13364, w_eco13365, w_eco13366, w_eco13367, w_eco13368, w_eco13369, w_eco13370, w_eco13371, w_eco13372, w_eco13373, w_eco13374, w_eco13375, w_eco13376, w_eco13377, w_eco13378, w_eco13379, w_eco13380, w_eco13381, w_eco13382, w_eco13383, w_eco13384, w_eco13385, w_eco13386, w_eco13387, w_eco13388, w_eco13389, w_eco13390, w_eco13391, w_eco13392, w_eco13393, w_eco13394, w_eco13395, w_eco13396, w_eco13397, w_eco13398, w_eco13399, w_eco13400, w_eco13401, w_eco13402, w_eco13403, w_eco13404, w_eco13405, w_eco13406, w_eco13407, w_eco13408, w_eco13409, w_eco13410, w_eco13411, w_eco13412, w_eco13413, w_eco13414, w_eco13415, w_eco13416, w_eco13417, w_eco13418, w_eco13419, w_eco13420, w_eco13421, w_eco13422, w_eco13423, w_eco13424, w_eco13425, w_eco13426, w_eco13427, w_eco13428, w_eco13429, w_eco13430, w_eco13431, w_eco13432, w_eco13433, w_eco13434, w_eco13435, w_eco13436, w_eco13437, w_eco13438, w_eco13439, w_eco13440, w_eco13441, w_eco13442, w_eco13443, w_eco13444, w_eco13445, w_eco13446, w_eco13447, w_eco13448, w_eco13449, w_eco13450, w_eco13451, w_eco13452, w_eco13453, w_eco13454, w_eco13455, w_eco13456, w_eco13457, w_eco13458, w_eco13459, w_eco13460, w_eco13461, w_eco13462, w_eco13463, w_eco13464, w_eco13465, w_eco13466, w_eco13467, w_eco13468, w_eco13469, w_eco13470, w_eco13471, w_eco13472, w_eco13473, w_eco13474, w_eco13475, w_eco13476, w_eco13477, w_eco13478, w_eco13479, w_eco13480, w_eco13481, w_eco13482, w_eco13483, w_eco13484, w_eco13485, w_eco13486, w_eco13487, w_eco13488, w_eco13489, w_eco13490, w_eco13491, w_eco13492, w_eco13493, w_eco13494, w_eco13495, w_eco13496, w_eco13497, w_eco13498, w_eco13499, w_eco13500, w_eco13501, w_eco13502, w_eco13503, w_eco13504, w_eco13505, w_eco13506, w_eco13507, w_eco13508, w_eco13509, w_eco13510, w_eco13511, w_eco13512, w_eco13513, w_eco13514, w_eco13515, w_eco13516, w_eco13517, w_eco13518, w_eco13519, w_eco13520, w_eco13521, w_eco13522, w_eco13523, w_eco13524, w_eco13525, w_eco13526, w_eco13527, w_eco13528, w_eco13529, w_eco13530, w_eco13531, w_eco13532, w_eco13533, w_eco13534, w_eco13535, w_eco13536, w_eco13537, w_eco13538, w_eco13539, w_eco13540, w_eco13541, w_eco13542, w_eco13543, w_eco13544, w_eco13545, w_eco13546, w_eco13547, w_eco13548, w_eco13549, w_eco13550, w_eco13551, w_eco13552, w_eco13553, w_eco13554, w_eco13555, w_eco13556, w_eco13557, w_eco13558, w_eco13559, w_eco13560, w_eco13561, w_eco13562, w_eco13563, w_eco13564, w_eco13565, w_eco13566, w_eco13567, w_eco13568, w_eco13569, w_eco13570, w_eco13571, w_eco13572, w_eco13573, w_eco13574, w_eco13575, w_eco13576, w_eco13577, w_eco13578, w_eco13579, w_eco13580, w_eco13581, w_eco13582, w_eco13583, w_eco13584, w_eco13585, w_eco13586, w_eco13587, w_eco13588, w_eco13589, w_eco13590, w_eco13591, w_eco13592, w_eco13593, w_eco13594, w_eco13595, w_eco13596, w_eco13597, w_eco13598, w_eco13599, w_eco13600, w_eco13601, w_eco13602, w_eco13603, w_eco13604, w_eco13605, w_eco13606, w_eco13607, w_eco13608, w_eco13609, w_eco13610, w_eco13611, w_eco13612, w_eco13613, w_eco13614, w_eco13615, w_eco13616, w_eco13617, w_eco13618, w_eco13619, w_eco13620, w_eco13621, w_eco13622, w_eco13623, w_eco13624, w_eco13625, w_eco13626, w_eco13627, w_eco13628, w_eco13629, w_eco13630, w_eco13631, w_eco13632, w_eco13633, w_eco13634, w_eco13635, w_eco13636, w_eco13637, w_eco13638, w_eco13639, w_eco13640, w_eco13641, w_eco13642, w_eco13643, w_eco13644, w_eco13645, w_eco13646, w_eco13647, w_eco13648, w_eco13649, w_eco13650, w_eco13651, w_eco13652, w_eco13653, w_eco13654, w_eco13655, w_eco13656, w_eco13657, w_eco13658, w_eco13659, w_eco13660, w_eco13661, w_eco13662, w_eco13663, w_eco13664, w_eco13665, w_eco13666, w_eco13667, w_eco13668, w_eco13669, w_eco13670, w_eco13671, w_eco13672, w_eco13673, w_eco13674, w_eco13675, w_eco13676, w_eco13677, w_eco13678, w_eco13679, w_eco13680, w_eco13681, w_eco13682, w_eco13683, w_eco13684, w_eco13685, w_eco13686, w_eco13687, w_eco13688, w_eco13689, w_eco13690, w_eco13691, w_eco13692, w_eco13693, w_eco13694, w_eco13695);
	xor _ECO_out11(cnt[14], sub_wire11, w_eco13696);
	and _ECO_13697(w_eco13697, prev_cnt[13], rst);
	and _ECO_13698(w_eco13698, prev_cnt[11], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13699(w_eco13699, prev_cnt[11], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13700(w_eco13700, prev_cnt[11], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13701(w_eco13701, prev_cnt[13], prev_cnt[15], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13702(w_eco13702, prev_cnt[11], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13703(w_eco13703, prev_cnt[12], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1], prev_state[0]);
	and _ECO_13704(w_eco13704, prev_cnt[12], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13705(w_eco13705, prev_cnt[9], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13706(w_eco13706, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13707(w_eco13707, prev_cnt[9], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13708(w_eco13708, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13709(w_eco13709, !prev_cnt[12], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13710(w_eco13710, !prev_cnt[14], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13711(w_eco13711, prev_cnt[12], prev_cnt[13], prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13712(w_eco13712, Tgate[13], prev_cnt[14], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13713(w_eco13713, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13714(w_eco13714, prev_cnt[6], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13715(w_eco13715, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13716(w_eco13716, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13717(w_eco13717, prev_cnt[6], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13718(w_eco13718, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13719(w_eco13719, prev_cnt[9], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13720(w_eco13720, prev_cnt[9], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13721(w_eco13721, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13722(w_eco13722, prev_cnt[8], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13723(w_eco13723, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13724(w_eco13724, Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13725(w_eco13725, Tgate[13], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13726(w_eco13726, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13727(w_eco13727, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13728(w_eco13728, prev_cnt[8], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13729(w_eco13729, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13730(w_eco13730, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13731(w_eco13731, prev_cnt[6], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13732(w_eco13732, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13733(w_eco13733, prev_cnt[6], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13734(w_eco13734, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13735(w_eco13735, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13736(w_eco13736, prev_cnt[10], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13737(w_eco13737, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13738(w_eco13738, Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13739(w_eco13739, Tgate[13], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13740(w_eco13740, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13741(w_eco13741, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13742(w_eco13742, prev_cnt[10], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13743(w_eco13743, Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13744(w_eco13744, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13745(w_eco13745, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13746(w_eco13746, prev_cnt[8], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13747(w_eco13747, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13748(w_eco13748, prev_cnt[8], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13749(w_eco13749, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13750(w_eco13750, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13751(w_eco13751, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13752(w_eco13752, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13753(w_eco13753, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13754(w_eco13754, Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13755(w_eco13755, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13756(w_eco13756, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13757(w_eco13757, Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13758(w_eco13758, Tgate[13], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13759(w_eco13759, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13760(w_eco13760, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13761(w_eco13761, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13762(w_eco13762, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13763(w_eco13763, prev_cnt[12], prev_cnt[13], prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13764(w_eco13764, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13765(w_eco13765, Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13766(w_eco13766, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13767(w_eco13767, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13768(w_eco13768, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13769(w_eco13769, prev_cnt[10], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13770(w_eco13770, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13771(w_eco13771, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13772(w_eco13772, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13773(w_eco13773, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13774(w_eco13774, prev_cnt[10], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13775(w_eco13775, Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13776(w_eco13776, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13777(w_eco13777, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13778(w_eco13778, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13779(w_eco13779, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13780(w_eco13780, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13781(w_eco13781, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13782(w_eco13782, !prev_cnt[14], prev_cnt[12], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13783(w_eco13783, Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13784(w_eco13784, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13785(w_eco13785, Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13786(w_eco13786, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13787(w_eco13787, Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13788(w_eco13788, Tgate[13], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13789(w_eco13789, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13790(w_eco13790, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13791(w_eco13791, Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13792(w_eco13792, Tgate[13], prev_cnt[14], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13793(w_eco13793, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13794(w_eco13794, !prev_cnt[14], prev_cnt[12], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13795(w_eco13795, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13796(w_eco13796, Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13797(w_eco13797, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13798(w_eco13798, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13799(w_eco13799, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13800(w_eco13800, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13801(w_eco13801, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13802(w_eco13802, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13803(w_eco13803, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13804(w_eco13804, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13805(w_eco13805, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13806(w_eco13806, Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13807(w_eco13807, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13808(w_eco13808, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13809(w_eco13809, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13810(w_eco13810, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13811(w_eco13811, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13812(w_eco13812, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13813(w_eco13813, Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13814(w_eco13814, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13815(w_eco13815, Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13816(w_eco13816, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13817(w_eco13817, Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13818(w_eco13818, Tgate[13], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13819(w_eco13819, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13820(w_eco13820, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_13821(w_eco13821, Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13822(w_eco13822, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13823(w_eco13823, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13824(w_eco13824, Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13825(w_eco13825, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_13826(w_eco13826, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13827(w_eco13827, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13828(w_eco13828, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13829(w_eco13829, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13830(w_eco13830, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13831(w_eco13831, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13832(w_eco13832, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13833(w_eco13833, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13834(w_eco13834, Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13835(w_eco13835, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13836(w_eco13836, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13837(w_eco13837, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13838(w_eco13838, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13839(w_eco13839, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13840(w_eco13840, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13841(w_eco13841, Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13842(w_eco13842, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13843(w_eco13843, Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13844(w_eco13844, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13845(w_eco13845, Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13846(w_eco13846, Tgate[13], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13847(w_eco13847, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13848(w_eco13848, Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13849(w_eco13849, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13850(w_eco13850, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13851(w_eco13851, Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13852(w_eco13852, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13853(w_eco13853, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13854(w_eco13854, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13855(w_eco13855, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13856(w_eco13856, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13857(w_eco13857, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13858(w_eco13858, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13859(w_eco13859, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13860(w_eco13860, Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13861(w_eco13861, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13862(w_eco13862, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13863(w_eco13863, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13864(w_eco13864, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13865(w_eco13865, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13866(w_eco13866, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13867(w_eco13867, Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13868(w_eco13868, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13869(w_eco13869, Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13870(w_eco13870, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13871(w_eco13871, Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[1]);
	and _ECO_13872(w_eco13872, Tgate[13], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1]);
	and _ECO_13873(w_eco13873, Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13874(w_eco13874, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13875(w_eco13875, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13876(w_eco13876, Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13877(w_eco13877, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13878(w_eco13878, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13879(w_eco13879, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_13880(w_eco13880, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13881(w_eco13881, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !ena, !rst);
	and _ECO_13882(w_eco13882, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13883(w_eco13883, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13884(w_eco13884, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, !prev_state[3], prev_state[0]);
	and _ECO_13885(w_eco13885, Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13886(w_eco13886, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13887(w_eco13887, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13888(w_eco13888, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_state[0]);
	and _ECO_13889(w_eco13889, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13890(w_eco13890, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13891(w_eco13891, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13892(w_eco13892, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13893(w_eco13893, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !rst, prev_state[0]);
	and _ECO_13894(w_eco13894, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13895(w_eco13895, Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13896(w_eco13896, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13897(w_eco13897, Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13898(w_eco13898, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13899(w_eco13899, Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13900(w_eco13900, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_13901(w_eco13901, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13902(w_eco13902, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13903(w_eco13903, Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_13904(w_eco13904, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13905(w_eco13905, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13906(w_eco13906, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_13907(w_eco13907, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13908(w_eco13908, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13909(w_eco13909, Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13910(w_eco13910, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13911(w_eco13911, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13912(w_eco13912, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13913(w_eco13913, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_13914(w_eco13914, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13915(w_eco13915, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_13916(w_eco13916, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13917(w_eco13917, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13918(w_eco13918, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13919(w_eco13919, Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13920(w_eco13920, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13921(w_eco13921, Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !ena, !rst);
	and _ECO_13922(w_eco13922, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_13923(w_eco13923, Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13924(w_eco13924, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13925(w_eco13925, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_13926(w_eco13926, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13927(w_eco13927, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_13928(w_eco13928, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13929(w_eco13929, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13930(w_eco13930, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_13931(w_eco13931, Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_13932(w_eco13932, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[13], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13933(w_eco13933, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_13934(w_eco13934, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_13935(w_eco13935, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13936(w_eco13936, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13937(w_eco13937, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_13938(w_eco13938, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13939(w_eco13939, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13940(w_eco13940, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13941(w_eco13941, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13942(w_eco13942, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13943(w_eco13943, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13944(w_eco13944, Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_13945(w_eco13945, Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[13], !prev_cnt[15], !rst, prev_state[0]);
	and _ECO_13946(w_eco13946, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[4], !prev_state[2]);
	and _ECO_13947(w_eco13947, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13948(w_eco13948, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13949(w_eco13949, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_13950(w_eco13950, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13951(w_eco13951, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13952(w_eco13952, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13953(w_eco13953, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13954(w_eco13954, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13955(w_eco13955, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13956(w_eco13956, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13957(w_eco13957, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13958(w_eco13958, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !prev_state[3], prev_state[0]);
	and _ECO_13959(w_eco13959, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13960(w_eco13960, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13961(w_eco13961, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13962(w_eco13962, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13963(w_eco13963, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13964(w_eco13964, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13965(w_eco13965, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13966(w_eco13966, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_13967(w_eco13967, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13968(w_eco13968, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13969(w_eco13969, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13970(w_eco13970, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13971(w_eco13971, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13972(w_eco13972, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13973(w_eco13973, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13974(w_eco13974, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13975(w_eco13975, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13976(w_eco13976, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13977(w_eco13977, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13978(w_eco13978, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13979(w_eco13979, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13980(w_eco13980, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13981(w_eco13981, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13982(w_eco13982, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13983(w_eco13983, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13984(w_eco13984, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13985(w_eco13985, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_13986(w_eco13986, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13987(w_eco13987, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_13988(w_eco13988, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13989(w_eco13989, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13990(w_eco13990, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13991(w_eco13991, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_13992(w_eco13992, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13993(w_eco13993, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_13994(w_eco13994, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13995(w_eco13995, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13996(w_eco13996, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_13997(w_eco13997, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_13998(w_eco13998, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_13999(w_eco13999, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14000(w_eco14000, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14001(w_eco14001, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14002(w_eco14002, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14003(w_eco14003, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14004(w_eco14004, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14005(w_eco14005, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14006(w_eco14006, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14007(w_eco14007, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14008(w_eco14008, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14009(w_eco14009, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14010(w_eco14010, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14011(w_eco14011, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14012(w_eco14012, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14013(w_eco14013, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14014(w_eco14014, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14015(w_eco14015, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14016(w_eco14016, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_14017(w_eco14017, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14018(w_eco14018, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14019(w_eco14019, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14020(w_eco14020, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14021(w_eco14021, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14022(w_eco14022, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14023(w_eco14023, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14024(w_eco14024, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14025(w_eco14025, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14026(w_eco14026, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14027(w_eco14027, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14028(w_eco14028, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14029(w_eco14029, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14030(w_eco14030, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14031(w_eco14031, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14032(w_eco14032, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14033(w_eco14033, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14034(w_eco14034, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14035(w_eco14035, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14036(w_eco14036, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14037(w_eco14037, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14038(w_eco14038, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14039(w_eco14039, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14040(w_eco14040, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14041(w_eco14041, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14042(w_eco14042, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14043(w_eco14043, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14044(w_eco14044, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14045(w_eco14045, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14046(w_eco14046, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14047(w_eco14047, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], prev_state[1]);
	and _ECO_14048(w_eco14048, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14049(w_eco14049, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14050(w_eco14050, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14051(w_eco14051, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14052(w_eco14052, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14053(w_eco14053, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14054(w_eco14054, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14055(w_eco14055, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14056(w_eco14056, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14057(w_eco14057, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14058(w_eco14058, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14059(w_eco14059, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14060(w_eco14060, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14061(w_eco14061, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14062(w_eco14062, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14063(w_eco14063, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14064(w_eco14064, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14065(w_eco14065, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14066(w_eco14066, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14067(w_eco14067, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14068(w_eco14068, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14069(w_eco14069, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14070(w_eco14070, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14071(w_eco14071, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14072(w_eco14072, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14073(w_eco14073, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14074(w_eco14074, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14075(w_eco14075, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14076(w_eco14076, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14077(w_eco14077, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14078(w_eco14078, !Tgate[13], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14079(w_eco14079, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14080(w_eco14080, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14081(w_eco14081, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14082(w_eco14082, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14083(w_eco14083, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14084(w_eco14084, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14085(w_eco14085, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14086(w_eco14086, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14087(w_eco14087, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14088(w_eco14088, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14089(w_eco14089, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14090(w_eco14090, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14091(w_eco14091, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14092(w_eco14092, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14093(w_eco14093, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14094(w_eco14094, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14095(w_eco14095, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14096(w_eco14096, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14097(w_eco14097, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14098(w_eco14098, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14099(w_eco14099, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14100(w_eco14100, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14101(w_eco14101, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14102(w_eco14102, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14103(w_eco14103, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14104(w_eco14104, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14105(w_eco14105, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14106(w_eco14106, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14107(w_eco14107, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14108(w_eco14108, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14109(w_eco14109, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14110(w_eco14110, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14111(w_eco14111, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14112(w_eco14112, !Tgate[13], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14113(w_eco14113, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14114(w_eco14114, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14115(w_eco14115, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14116(w_eco14116, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14117(w_eco14117, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14118(w_eco14118, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14119(w_eco14119, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14120(w_eco14120, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14121(w_eco14121, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14122(w_eco14122, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14123(w_eco14123, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14124(w_eco14124, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14125(w_eco14125, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14126(w_eco14126, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14127(w_eco14127, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14128(w_eco14128, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14129(w_eco14129, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14130(w_eco14130, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14131(w_eco14131, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14132(w_eco14132, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14133(w_eco14133, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14134(w_eco14134, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14135(w_eco14135, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14136(w_eco14136, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14137(w_eco14137, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14138(w_eco14138, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14139(w_eco14139, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14140(w_eco14140, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14141(w_eco14141, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14142(w_eco14142, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14143(w_eco14143, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14144(w_eco14144, !Tgate[13], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14145(w_eco14145, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14146(w_eco14146, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14147(w_eco14147, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14148(w_eco14148, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14149(w_eco14149, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14150(w_eco14150, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14151(w_eco14151, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14152(w_eco14152, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14153(w_eco14153, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14154(w_eco14154, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14155(w_eco14155, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14156(w_eco14156, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14157(w_eco14157, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14158(w_eco14158, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14159(w_eco14159, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14160(w_eco14160, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14161(w_eco14161, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14162(w_eco14162, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14163(w_eco14163, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14164(w_eco14164, !Tgate[13], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14165(w_eco14165, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14166(w_eco14166, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14167(w_eco14167, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14168(w_eco14168, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14169(w_eco14169, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14170(w_eco14170, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14171(w_eco14171, !Tgate[13], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14172(w_eco14172, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14173(w_eco14173, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14174(w_eco14174, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14175(w_eco14175, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14176(w_eco14176, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14177(w_eco14177, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14178(w_eco14178, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14179(w_eco14179, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14180(w_eco14180, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14181(w_eco14181, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14182(w_eco14182, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14183(w_eco14183, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14184(w_eco14184, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14185(w_eco14185, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14186(w_eco14186, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14187(w_eco14187, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14188(w_eco14188, !Tgate[13], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14189(w_eco14189, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14190(w_eco14190, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14191(w_eco14191, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14192(w_eco14192, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14193(w_eco14193, !Tgate[13], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14194(w_eco14194, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14195(w_eco14195, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14196(w_eco14196, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14197(w_eco14197, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14198(w_eco14198, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14199(w_eco14199, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14200(w_eco14200, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14201(w_eco14201, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14202(w_eco14202, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14203(w_eco14203, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14204(w_eco14204, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14205(w_eco14205, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14206(w_eco14206, !Tgate[13], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14207(w_eco14207, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14208(w_eco14208, !Tgate[13], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14209(w_eco14209, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14210(w_eco14210, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14211(w_eco14211, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14212(w_eco14212, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14213(w_eco14213, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14214(w_eco14214, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14215(w_eco14215, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14216(w_eco14216, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14217(w_eco14217, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14218(w_eco14218, !Tgate[13], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14219(w_eco14219, !Tgate[13], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14220(w_eco14220, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14221(w_eco14221, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14222(w_eco14222, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14223(w_eco14223, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14224(w_eco14224, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_14225(w_eco14225, !Tgate[13], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14226(w_eco14226, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, prev_state[2], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14227(w_eco14227, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14228(w_eco14228, !Tgate[13], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_14229(w_eco14229, !Tgate[13], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !prev_cnt[15], ena, !prev_state[4], !prev_state[3], prev_state[1], !prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_14230(w_eco14230, w_eco13697, w_eco13698, w_eco13699, w_eco13700, w_eco13701, w_eco13702, w_eco13703, w_eco13704, w_eco13705, w_eco13706, w_eco13707, w_eco13708, w_eco13709, w_eco13710, w_eco13711, w_eco13712, w_eco13713, w_eco13714, w_eco13715, w_eco13716, w_eco13717, w_eco13718, w_eco13719, w_eco13720, w_eco13721, w_eco13722, w_eco13723, w_eco13724, w_eco13725, w_eco13726, w_eco13727, w_eco13728, w_eco13729, w_eco13730, w_eco13731, w_eco13732, w_eco13733, w_eco13734, w_eco13735, w_eco13736, w_eco13737, w_eco13738, w_eco13739, w_eco13740, w_eco13741, w_eco13742, w_eco13743, w_eco13744, w_eco13745, w_eco13746, w_eco13747, w_eco13748, w_eco13749, w_eco13750, w_eco13751, w_eco13752, w_eco13753, w_eco13754, w_eco13755, w_eco13756, w_eco13757, w_eco13758, w_eco13759, w_eco13760, w_eco13761, w_eco13762, w_eco13763, w_eco13764, w_eco13765, w_eco13766, w_eco13767, w_eco13768, w_eco13769, w_eco13770, w_eco13771, w_eco13772, w_eco13773, w_eco13774, w_eco13775, w_eco13776, w_eco13777, w_eco13778, w_eco13779, w_eco13780, w_eco13781, w_eco13782, w_eco13783, w_eco13784, w_eco13785, w_eco13786, w_eco13787, w_eco13788, w_eco13789, w_eco13790, w_eco13791, w_eco13792, w_eco13793, w_eco13794, w_eco13795, w_eco13796, w_eco13797, w_eco13798, w_eco13799, w_eco13800, w_eco13801, w_eco13802, w_eco13803, w_eco13804, w_eco13805, w_eco13806, w_eco13807, w_eco13808, w_eco13809, w_eco13810, w_eco13811, w_eco13812, w_eco13813, w_eco13814, w_eco13815, w_eco13816, w_eco13817, w_eco13818, w_eco13819, w_eco13820, w_eco13821, w_eco13822, w_eco13823, w_eco13824, w_eco13825, w_eco13826, w_eco13827, w_eco13828, w_eco13829, w_eco13830, w_eco13831, w_eco13832, w_eco13833, w_eco13834, w_eco13835, w_eco13836, w_eco13837, w_eco13838, w_eco13839, w_eco13840, w_eco13841, w_eco13842, w_eco13843, w_eco13844, w_eco13845, w_eco13846, w_eco13847, w_eco13848, w_eco13849, w_eco13850, w_eco13851, w_eco13852, w_eco13853, w_eco13854, w_eco13855, w_eco13856, w_eco13857, w_eco13858, w_eco13859, w_eco13860, w_eco13861, w_eco13862, w_eco13863, w_eco13864, w_eco13865, w_eco13866, w_eco13867, w_eco13868, w_eco13869, w_eco13870, w_eco13871, w_eco13872, w_eco13873, w_eco13874, w_eco13875, w_eco13876, w_eco13877, w_eco13878, w_eco13879, w_eco13880, w_eco13881, w_eco13882, w_eco13883, w_eco13884, w_eco13885, w_eco13886, w_eco13887, w_eco13888, w_eco13889, w_eco13890, w_eco13891, w_eco13892, w_eco13893, w_eco13894, w_eco13895, w_eco13896, w_eco13897, w_eco13898, w_eco13899, w_eco13900, w_eco13901, w_eco13902, w_eco13903, w_eco13904, w_eco13905, w_eco13906, w_eco13907, w_eco13908, w_eco13909, w_eco13910, w_eco13911, w_eco13912, w_eco13913, w_eco13914, w_eco13915, w_eco13916, w_eco13917, w_eco13918, w_eco13919, w_eco13920, w_eco13921, w_eco13922, w_eco13923, w_eco13924, w_eco13925, w_eco13926, w_eco13927, w_eco13928, w_eco13929, w_eco13930, w_eco13931, w_eco13932, w_eco13933, w_eco13934, w_eco13935, w_eco13936, w_eco13937, w_eco13938, w_eco13939, w_eco13940, w_eco13941, w_eco13942, w_eco13943, w_eco13944, w_eco13945, w_eco13946, w_eco13947, w_eco13948, w_eco13949, w_eco13950, w_eco13951, w_eco13952, w_eco13953, w_eco13954, w_eco13955, w_eco13956, w_eco13957, w_eco13958, w_eco13959, w_eco13960, w_eco13961, w_eco13962, w_eco13963, w_eco13964, w_eco13965, w_eco13966, w_eco13967, w_eco13968, w_eco13969, w_eco13970, w_eco13971, w_eco13972, w_eco13973, w_eco13974, w_eco13975, w_eco13976, w_eco13977, w_eco13978, w_eco13979, w_eco13980, w_eco13981, w_eco13982, w_eco13983, w_eco13984, w_eco13985, w_eco13986, w_eco13987, w_eco13988, w_eco13989, w_eco13990, w_eco13991, w_eco13992, w_eco13993, w_eco13994, w_eco13995, w_eco13996, w_eco13997, w_eco13998, w_eco13999, w_eco14000, w_eco14001, w_eco14002, w_eco14003, w_eco14004, w_eco14005, w_eco14006, w_eco14007, w_eco14008, w_eco14009, w_eco14010, w_eco14011, w_eco14012, w_eco14013, w_eco14014, w_eco14015, w_eco14016, w_eco14017, w_eco14018, w_eco14019, w_eco14020, w_eco14021, w_eco14022, w_eco14023, w_eco14024, w_eco14025, w_eco14026, w_eco14027, w_eco14028, w_eco14029, w_eco14030, w_eco14031, w_eco14032, w_eco14033, w_eco14034, w_eco14035, w_eco14036, w_eco14037, w_eco14038, w_eco14039, w_eco14040, w_eco14041, w_eco14042, w_eco14043, w_eco14044, w_eco14045, w_eco14046, w_eco14047, w_eco14048, w_eco14049, w_eco14050, w_eco14051, w_eco14052, w_eco14053, w_eco14054, w_eco14055, w_eco14056, w_eco14057, w_eco14058, w_eco14059, w_eco14060, w_eco14061, w_eco14062, w_eco14063, w_eco14064, w_eco14065, w_eco14066, w_eco14067, w_eco14068, w_eco14069, w_eco14070, w_eco14071, w_eco14072, w_eco14073, w_eco14074, w_eco14075, w_eco14076, w_eco14077, w_eco14078, w_eco14079, w_eco14080, w_eco14081, w_eco14082, w_eco14083, w_eco14084, w_eco14085, w_eco14086, w_eco14087, w_eco14088, w_eco14089, w_eco14090, w_eco14091, w_eco14092, w_eco14093, w_eco14094, w_eco14095, w_eco14096, w_eco14097, w_eco14098, w_eco14099, w_eco14100, w_eco14101, w_eco14102, w_eco14103, w_eco14104, w_eco14105, w_eco14106, w_eco14107, w_eco14108, w_eco14109, w_eco14110, w_eco14111, w_eco14112, w_eco14113, w_eco14114, w_eco14115, w_eco14116, w_eco14117, w_eco14118, w_eco14119, w_eco14120, w_eco14121, w_eco14122, w_eco14123, w_eco14124, w_eco14125, w_eco14126, w_eco14127, w_eco14128, w_eco14129, w_eco14130, w_eco14131, w_eco14132, w_eco14133, w_eco14134, w_eco14135, w_eco14136, w_eco14137, w_eco14138, w_eco14139, w_eco14140, w_eco14141, w_eco14142, w_eco14143, w_eco14144, w_eco14145, w_eco14146, w_eco14147, w_eco14148, w_eco14149, w_eco14150, w_eco14151, w_eco14152, w_eco14153, w_eco14154, w_eco14155, w_eco14156, w_eco14157, w_eco14158, w_eco14159, w_eco14160, w_eco14161, w_eco14162, w_eco14163, w_eco14164, w_eco14165, w_eco14166, w_eco14167, w_eco14168, w_eco14169, w_eco14170, w_eco14171, w_eco14172, w_eco14173, w_eco14174, w_eco14175, w_eco14176, w_eco14177, w_eco14178, w_eco14179, w_eco14180, w_eco14181, w_eco14182, w_eco14183, w_eco14184, w_eco14185, w_eco14186, w_eco14187, w_eco14188, w_eco14189, w_eco14190, w_eco14191, w_eco14192, w_eco14193, w_eco14194, w_eco14195, w_eco14196, w_eco14197, w_eco14198, w_eco14199, w_eco14200, w_eco14201, w_eco14202, w_eco14203, w_eco14204, w_eco14205, w_eco14206, w_eco14207, w_eco14208, w_eco14209, w_eco14210, w_eco14211, w_eco14212, w_eco14213, w_eco14214, w_eco14215, w_eco14216, w_eco14217, w_eco14218, w_eco14219, w_eco14220, w_eco14221, w_eco14222, w_eco14223, w_eco14224, w_eco14225, w_eco14226, w_eco14227, w_eco14228, w_eco14229);
	xor _ECO_out12(cnt[13], sub_wire12, w_eco14230);
	and _ECO_14231(w_eco14231, prev_cnt[12], rst);
	and _ECO_14232(w_eco14232, prev_cnt[12], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14233(w_eco14233, prev_cnt[11], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14234(w_eco14234, prev_cnt[11], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14235(w_eco14235, prev_cnt[11], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14236(w_eco14236, prev_cnt[9], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14237(w_eco14237, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14238(w_eco14238, prev_cnt[9], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14239(w_eco14239, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14240(w_eco14240, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14241(w_eco14241, prev_cnt[6], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14242(w_eco14242, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14243(w_eco14243, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14244(w_eco14244, prev_cnt[6], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14245(w_eco14245, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14246(w_eco14246, prev_cnt[9], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14247(w_eco14247, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14248(w_eco14248, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14249(w_eco14249, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14250(w_eco14250, prev_cnt[8], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14251(w_eco14251, Tgate[12], !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14252(w_eco14252, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14253(w_eco14253, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14254(w_eco14254, prev_cnt[8], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14255(w_eco14255, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14256(w_eco14256, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14257(w_eco14257, prev_cnt[6], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14258(w_eco14258, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14259(w_eco14259, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14260(w_eco14260, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14261(w_eco14261, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14262(w_eco14262, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14263(w_eco14263, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14264(w_eco14264, prev_cnt[10], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14265(w_eco14265, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14266(w_eco14266, prev_cnt[10], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14267(w_eco14267, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14268(w_eco14268, prev_cnt[8], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14269(w_eco14269, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14270(w_eco14270, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14271(w_eco14271, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14272(w_eco14272, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14273(w_eco14273, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14274(w_eco14274, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14275(w_eco14275, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14276(w_eco14276, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14277(w_eco14277, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14278(w_eco14278, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14279(w_eco14279, Tgate[12], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14280(w_eco14280, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14281(w_eco14281, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14282(w_eco14282, Tgate[12], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14283(w_eco14283, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14284(w_eco14284, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14285(w_eco14285, prev_cnt[10], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14286(w_eco14286, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14287(w_eco14287, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14288(w_eco14288, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14289(w_eco14289, Tgate[12], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14290(w_eco14290, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14291(w_eco14291, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14292(w_eco14292, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14293(w_eco14293, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14294(w_eco14294, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14295(w_eco14295, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14296(w_eco14296, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14297(w_eco14297, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14298(w_eco14298, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14299(w_eco14299, Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14300(w_eco14300, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14301(w_eco14301, Tgate[12], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14302(w_eco14302, Tgate[12], !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14303(w_eco14303, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14304(w_eco14304, Tgate[12], prev_cnt[14], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14305(w_eco14305, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14306(w_eco14306, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14307(w_eco14307, Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14308(w_eco14308, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14309(w_eco14309, Tgate[12], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14310(w_eco14310, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14311(w_eco14311, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14312(w_eco14312, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14313(w_eco14313, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14314(w_eco14314, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14315(w_eco14315, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14316(w_eco14316, Tgate[12], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14317(w_eco14317, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14318(w_eco14318, Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14319(w_eco14319, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14320(w_eco14320, Tgate[12], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14321(w_eco14321, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14322(w_eco14322, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14323(w_eco14323, Tgate[12], !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14324(w_eco14324, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14325(w_eco14325, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14326(w_eco14326, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14327(w_eco14327, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14328(w_eco14328, Tgate[12], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14329(w_eco14329, Tgate[12], !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14330(w_eco14330, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14331(w_eco14331, Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14332(w_eco14332, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14333(w_eco14333, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14334(w_eco14334, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14335(w_eco14335, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14336(w_eco14336, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14337(w_eco14337, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14338(w_eco14338, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14339(w_eco14339, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14340(w_eco14340, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14341(w_eco14341, Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14342(w_eco14342, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14343(w_eco14343, Tgate[12], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], ena, !rst, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14344(w_eco14344, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14345(w_eco14345, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14346(w_eco14346, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14347(w_eco14347, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14348(w_eco14348, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_state[0]);
	and _ECO_14349(w_eco14349, Tgate[12], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14350(w_eco14350, Tgate[12], !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14351(w_eco14351, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14352(w_eco14352, Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14353(w_eco14353, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14354(w_eco14354, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14355(w_eco14355, Tgate[12], prev_cnt[14], prev_cnt[12], !prev_cnt[15], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14356(w_eco14356, Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14357(w_eco14357, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14358(w_eco14358, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14359(w_eco14359, Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14360(w_eco14360, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14361(w_eco14361, Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14362(w_eco14362, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14363(w_eco14363, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14364(w_eco14364, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14365(w_eco14365, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14366(w_eco14366, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14367(w_eco14367, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14368(w_eco14368, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_14369(w_eco14369, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14370(w_eco14370, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14371(w_eco14371, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14372(w_eco14372, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14373(w_eco14373, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14374(w_eco14374, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !ena, !rst);
	and _ECO_14375(w_eco14375, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14376(w_eco14376, Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14377(w_eco14377, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14378(w_eco14378, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14379(w_eco14379, Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14380(w_eco14380, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14381(w_eco14381, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14382(w_eco14382, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14383(w_eco14383, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14384(w_eco14384, Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14385(w_eco14385, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14386(w_eco14386, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14387(w_eco14387, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14388(w_eco14388, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14389(w_eco14389, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14390(w_eco14390, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14391(w_eco14391, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14392(w_eco14392, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14393(w_eco14393, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_14394(w_eco14394, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14395(w_eco14395, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14396(w_eco14396, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14397(w_eco14397, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14398(w_eco14398, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14399(w_eco14399, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14400(w_eco14400, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14401(w_eco14401, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14402(w_eco14402, !Tgate[12], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14403(w_eco14403, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !ena, !rst);
	and _ECO_14404(w_eco14404, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[0]);
	and _ECO_14405(w_eco14405, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14406(w_eco14406, Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14407(w_eco14407, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14408(w_eco14408, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14409(w_eco14409, Tgate[12], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14410(w_eco14410, Tgate[12], !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14411(w_eco14411, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14412(w_eco14412, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14413(w_eco14413, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14414(w_eco14414, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14415(w_eco14415, Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14416(w_eco14416, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14417(w_eco14417, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14418(w_eco14418, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14419(w_eco14419, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14420(w_eco14420, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14421(w_eco14421, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_14422(w_eco14422, Tgate[12], prev_cnt[14], prev_cnt[12], !prev_cnt[15], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14423(w_eco14423, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[12], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14424(w_eco14424, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14425(w_eco14425, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14426(w_eco14426, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14427(w_eco14427, !Tgate[12], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14428(w_eco14428, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14429(w_eco14429, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14430(w_eco14430, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !ena);
	and _ECO_14431(w_eco14431, Tgate[12], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14432(w_eco14432, Tgate[12], !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14433(w_eco14433, Tgate[12], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst);
	and _ECO_14434(w_eco14434, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14435(w_eco14435, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14436(w_eco14436, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14437(w_eco14437, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[4], !prev_state[2]);
	and _ECO_14438(w_eco14438, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14439(w_eco14439, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_cnt[15], !prev_state[3], prev_state[0]);
	and _ECO_14440(w_eco14440, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14441(w_eco14441, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14442(w_eco14442, !Tgate[12], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14443(w_eco14443, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14444(w_eco14444, Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14445(w_eco14445, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14446(w_eco14446, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14447(w_eco14447, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14448(w_eco14448, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14449(w_eco14449, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[4], !prev_state[2]);
	and _ECO_14450(w_eco14450, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14451(w_eco14451, !Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14452(w_eco14452, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14453(w_eco14453, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14454(w_eco14454, Tgate[12], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14455(w_eco14455, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14456(w_eco14456, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !ena, !rst);
	and _ECO_14457(w_eco14457, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !prev_state[3], prev_state[0]);
	and _ECO_14458(w_eco14458, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14459(w_eco14459, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14460(w_eco14460, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14461(w_eco14461, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14462(w_eco14462, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14463(w_eco14463, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14464(w_eco14464, !Tgate[12], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14465(w_eco14465, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14466(w_eco14466, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14467(w_eco14467, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14468(w_eco14468, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14469(w_eco14469, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14470(w_eco14470, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14471(w_eco14471, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14472(w_eco14472, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14473(w_eco14473, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14474(w_eco14474, !Tgate[12], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14475(w_eco14475, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14476(w_eco14476, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14477(w_eco14477, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14478(w_eco14478, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14479(w_eco14479, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14480(w_eco14480, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14481(w_eco14481, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14482(w_eco14482, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14483(w_eco14483, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14484(w_eco14484, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14485(w_eco14485, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14486(w_eco14486, !Tgate[12], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], prev_state[1]);
	and _ECO_14487(w_eco14487, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14488(w_eco14488, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14489(w_eco14489, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14490(w_eco14490, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14491(w_eco14491, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14492(w_eco14492, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14493(w_eco14493, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14494(w_eco14494, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14495(w_eco14495, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14496(w_eco14496, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14497(w_eco14497, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14498(w_eco14498, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14499(w_eco14499, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14500(w_eco14500, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14501(w_eco14501, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14502(w_eco14502, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14503(w_eco14503, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14504(w_eco14504, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14505(w_eco14505, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14506(w_eco14506, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14507(w_eco14507, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14508(w_eco14508, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14509(w_eco14509, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14510(w_eco14510, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14511(w_eco14511, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14512(w_eco14512, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14513(w_eco14513, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14514(w_eco14514, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14515(w_eco14515, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14516(w_eco14516, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14517(w_eco14517, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14518(w_eco14518, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14519(w_eco14519, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14520(w_eco14520, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14521(w_eco14521, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14522(w_eco14522, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14523(w_eco14523, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14524(w_eco14524, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14525(w_eco14525, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14526(w_eco14526, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14527(w_eco14527, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14528(w_eco14528, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14529(w_eco14529, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14530(w_eco14530, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14531(w_eco14531, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14532(w_eco14532, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14533(w_eco14533, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14534(w_eco14534, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14535(w_eco14535, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14536(w_eco14536, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14537(w_eco14537, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14538(w_eco14538, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14539(w_eco14539, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14540(w_eco14540, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14541(w_eco14541, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14542(w_eco14542, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14543(w_eco14543, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14544(w_eco14544, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14545(w_eco14545, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14546(w_eco14546, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14547(w_eco14547, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14548(w_eco14548, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14549(w_eco14549, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14550(w_eco14550, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14551(w_eco14551, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14552(w_eco14552, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14553(w_eco14553, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14554(w_eco14554, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14555(w_eco14555, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14556(w_eco14556, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14557(w_eco14557, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14558(w_eco14558, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14559(w_eco14559, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14560(w_eco14560, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14561(w_eco14561, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14562(w_eco14562, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_14563(w_eco14563, w_eco14231, w_eco14232, w_eco14233, w_eco14234, w_eco14235, w_eco14236, w_eco14237, w_eco14238, w_eco14239, w_eco14240, w_eco14241, w_eco14242, w_eco14243, w_eco14244, w_eco14245, w_eco14246, w_eco14247, w_eco14248, w_eco14249, w_eco14250, w_eco14251, w_eco14252, w_eco14253, w_eco14254, w_eco14255, w_eco14256, w_eco14257, w_eco14258, w_eco14259, w_eco14260, w_eco14261, w_eco14262, w_eco14263, w_eco14264, w_eco14265, w_eco14266, w_eco14267, w_eco14268, w_eco14269, w_eco14270, w_eco14271, w_eco14272, w_eco14273, w_eco14274, w_eco14275, w_eco14276, w_eco14277, w_eco14278, w_eco14279, w_eco14280, w_eco14281, w_eco14282, w_eco14283, w_eco14284, w_eco14285, w_eco14286, w_eco14287, w_eco14288, w_eco14289, w_eco14290, w_eco14291, w_eco14292, w_eco14293, w_eco14294, w_eco14295, w_eco14296, w_eco14297, w_eco14298, w_eco14299, w_eco14300, w_eco14301, w_eco14302, w_eco14303, w_eco14304, w_eco14305, w_eco14306, w_eco14307, w_eco14308, w_eco14309, w_eco14310, w_eco14311, w_eco14312, w_eco14313, w_eco14314, w_eco14315, w_eco14316, w_eco14317, w_eco14318, w_eco14319, w_eco14320, w_eco14321, w_eco14322, w_eco14323, w_eco14324, w_eco14325, w_eco14326, w_eco14327, w_eco14328, w_eco14329, w_eco14330, w_eco14331, w_eco14332, w_eco14333, w_eco14334, w_eco14335, w_eco14336, w_eco14337, w_eco14338, w_eco14339, w_eco14340, w_eco14341, w_eco14342, w_eco14343, w_eco14344, w_eco14345, w_eco14346, w_eco14347, w_eco14348, w_eco14349, w_eco14350, w_eco14351, w_eco14352, w_eco14353, w_eco14354, w_eco14355, w_eco14356, w_eco14357, w_eco14358, w_eco14359, w_eco14360, w_eco14361, w_eco14362, w_eco14363, w_eco14364, w_eco14365, w_eco14366, w_eco14367, w_eco14368, w_eco14369, w_eco14370, w_eco14371, w_eco14372, w_eco14373, w_eco14374, w_eco14375, w_eco14376, w_eco14377, w_eco14378, w_eco14379, w_eco14380, w_eco14381, w_eco14382, w_eco14383, w_eco14384, w_eco14385, w_eco14386, w_eco14387, w_eco14388, w_eco14389, w_eco14390, w_eco14391, w_eco14392, w_eco14393, w_eco14394, w_eco14395, w_eco14396, w_eco14397, w_eco14398, w_eco14399, w_eco14400, w_eco14401, w_eco14402, w_eco14403, w_eco14404, w_eco14405, w_eco14406, w_eco14407, w_eco14408, w_eco14409, w_eco14410, w_eco14411, w_eco14412, w_eco14413, w_eco14414, w_eco14415, w_eco14416, w_eco14417, w_eco14418, w_eco14419, w_eco14420, w_eco14421, w_eco14422, w_eco14423, w_eco14424, w_eco14425, w_eco14426, w_eco14427, w_eco14428, w_eco14429, w_eco14430, w_eco14431, w_eco14432, w_eco14433, w_eco14434, w_eco14435, w_eco14436, w_eco14437, w_eco14438, w_eco14439, w_eco14440, w_eco14441, w_eco14442, w_eco14443, w_eco14444, w_eco14445, w_eco14446, w_eco14447, w_eco14448, w_eco14449, w_eco14450, w_eco14451, w_eco14452, w_eco14453, w_eco14454, w_eco14455, w_eco14456, w_eco14457, w_eco14458, w_eco14459, w_eco14460, w_eco14461, w_eco14462, w_eco14463, w_eco14464, w_eco14465, w_eco14466, w_eco14467, w_eco14468, w_eco14469, w_eco14470, w_eco14471, w_eco14472, w_eco14473, w_eco14474, w_eco14475, w_eco14476, w_eco14477, w_eco14478, w_eco14479, w_eco14480, w_eco14481, w_eco14482, w_eco14483, w_eco14484, w_eco14485, w_eco14486, w_eco14487, w_eco14488, w_eco14489, w_eco14490, w_eco14491, w_eco14492, w_eco14493, w_eco14494, w_eco14495, w_eco14496, w_eco14497, w_eco14498, w_eco14499, w_eco14500, w_eco14501, w_eco14502, w_eco14503, w_eco14504, w_eco14505, w_eco14506, w_eco14507, w_eco14508, w_eco14509, w_eco14510, w_eco14511, w_eco14512, w_eco14513, w_eco14514, w_eco14515, w_eco14516, w_eco14517, w_eco14518, w_eco14519, w_eco14520, w_eco14521, w_eco14522, w_eco14523, w_eco14524, w_eco14525, w_eco14526, w_eco14527, w_eco14528, w_eco14529, w_eco14530, w_eco14531, w_eco14532, w_eco14533, w_eco14534, w_eco14535, w_eco14536, w_eco14537, w_eco14538, w_eco14539, w_eco14540, w_eco14541, w_eco14542, w_eco14543, w_eco14544, w_eco14545, w_eco14546, w_eco14547, w_eco14548, w_eco14549, w_eco14550, w_eco14551, w_eco14552, w_eco14553, w_eco14554, w_eco14555, w_eco14556, w_eco14557, w_eco14558, w_eco14559, w_eco14560, w_eco14561, w_eco14562);
	xor _ECO_out13(cnt[12], sub_wire13, w_eco14563);
	and _ECO_14564(w_eco14564, prev_cnt[11], rst);
	and _ECO_14565(w_eco14565, prev_cnt[11], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14566(w_eco14566, prev_cnt[9], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14567(w_eco14567, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14568(w_eco14568, prev_cnt[9], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14569(w_eco14569, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14570(w_eco14570, prev_cnt[9], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14571(w_eco14571, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14572(w_eco14572, prev_cnt[6], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14573(w_eco14573, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14574(w_eco14574, prev_cnt[6], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14575(w_eco14575, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14576(w_eco14576, prev_cnt[6], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14577(w_eco14577, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14578(w_eco14578, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14579(w_eco14579, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14580(w_eco14580, prev_cnt[8], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14581(w_eco14581, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14582(w_eco14582, prev_cnt[8], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14583(w_eco14583, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14584(w_eco14584, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14585(w_eco14585, prev_cnt[8], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14586(w_eco14586, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14587(w_eco14587, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14588(w_eco14588, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14589(w_eco14589, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14590(w_eco14590, prev_cnt[10], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14591(w_eco14591, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14592(w_eco14592, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14593(w_eco14593, prev_cnt[10], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14594(w_eco14594, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14595(w_eco14595, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14596(w_eco14596, prev_cnt[10], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14597(w_eco14597, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14598(w_eco14598, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14599(w_eco14599, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14600(w_eco14600, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14601(w_eco14601, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14602(w_eco14602, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14603(w_eco14603, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14604(w_eco14604, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14605(w_eco14605, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14606(w_eco14606, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14607(w_eco14607, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14608(w_eco14608, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14609(w_eco14609, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14610(w_eco14610, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14611(w_eco14611, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14612(w_eco14612, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14613(w_eco14613, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14614(w_eco14614, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14615(w_eco14615, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14616(w_eco14616, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14617(w_eco14617, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14618(w_eco14618, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14619(w_eco14619, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14620(w_eco14620, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14621(w_eco14621, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14622(w_eco14622, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14623(w_eco14623, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14624(w_eco14624, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14625(w_eco14625, Tgate[11], prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14626(w_eco14626, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14627(w_eco14627, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14628(w_eco14628, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14629(w_eco14629, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14630(w_eco14630, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14631(w_eco14631, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14632(w_eco14632, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14633(w_eco14633, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14634(w_eco14634, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14635(w_eco14635, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14636(w_eco14636, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !ena, !rst);
	and _ECO_14637(w_eco14637, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14638(w_eco14638, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14639(w_eco14639, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14640(w_eco14640, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14641(w_eco14641, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14642(w_eco14642, Tgate[11], prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14643(w_eco14643, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14644(w_eco14644, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14645(w_eco14645, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14646(w_eco14646, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14647(w_eco14647, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14648(w_eco14648, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14649(w_eco14649, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14650(w_eco14650, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14651(w_eco14651, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_state[0]);
	and _ECO_14652(w_eco14652, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14653(w_eco14653, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14654(w_eco14654, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14655(w_eco14655, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14656(w_eco14656, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14657(w_eco14657, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14658(w_eco14658, Tgate[11], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14659(w_eco14659, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14660(w_eco14660, Tgate[11], prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14661(w_eco14661, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14662(w_eco14662, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14663(w_eco14663, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14664(w_eco14664, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14665(w_eco14665, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14666(w_eco14666, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14667(w_eco14667, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14668(w_eco14668, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14669(w_eco14669, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14670(w_eco14670, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14671(w_eco14671, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14672(w_eco14672, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14673(w_eco14673, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14674(w_eco14674, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !rst, prev_state[0]);
	and _ECO_14675(w_eco14675, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14676(w_eco14676, Tgate[11], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14677(w_eco14677, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14678(w_eco14678, Tgate[11], prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14679(w_eco14679, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14680(w_eco14680, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14681(w_eco14681, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14682(w_eco14682, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14683(w_eco14683, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14684(w_eco14684, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14685(w_eco14685, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14686(w_eco14686, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14687(w_eco14687, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14688(w_eco14688, Tgate[11], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14689(w_eco14689, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14690(w_eco14690, Tgate[11], prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14691(w_eco14691, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14692(w_eco14692, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14693(w_eco14693, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14694(w_eco14694, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14695(w_eco14695, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[11], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14696(w_eco14696, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14697(w_eco14697, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14698(w_eco14698, Tgate[11], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14699(w_eco14699, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14700(w_eco14700, Tgate[11], prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14701(w_eco14701, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14702(w_eco14702, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14703(w_eco14703, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14704(w_eco14704, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14705(w_eco14705, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14706(w_eco14706, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14707(w_eco14707, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14708(w_eco14708, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14709(w_eco14709, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14710(w_eco14710, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14711(w_eco14711, Tgate[11], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14712(w_eco14712, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14713(w_eco14713, Tgate[11], prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst);
	and _ECO_14714(w_eco14714, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14715(w_eco14715, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14716(w_eco14716, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14717(w_eco14717, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14718(w_eco14718, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14719(w_eco14719, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14720(w_eco14720, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14721(w_eco14721, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14722(w_eco14722, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14723(w_eco14723, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14724(w_eco14724, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14725(w_eco14725, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14726(w_eco14726, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14727(w_eco14727, Tgate[11], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14728(w_eco14728, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14729(w_eco14729, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14730(w_eco14730, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14731(w_eco14731, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14732(w_eco14732, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14733(w_eco14733, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14734(w_eco14734, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14735(w_eco14735, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14736(w_eco14736, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14737(w_eco14737, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14738(w_eco14738, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14739(w_eco14739, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], prev_state[1]);
	and _ECO_14740(w_eco14740, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14741(w_eco14741, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14742(w_eco14742, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14743(w_eco14743, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14744(w_eco14744, Tgate[11], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst);
	and _ECO_14745(w_eco14745, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14746(w_eco14746, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14747(w_eco14747, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14748(w_eco14748, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14749(w_eco14749, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14750(w_eco14750, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14751(w_eco14751, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14752(w_eco14752, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14753(w_eco14753, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14754(w_eco14754, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14755(w_eco14755, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14756(w_eco14756, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14757(w_eco14757, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14758(w_eco14758, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14759(w_eco14759, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14760(w_eco14760, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14761(w_eco14761, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14762(w_eco14762, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14763(w_eco14763, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14764(w_eco14764, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_14765(w_eco14765, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14766(w_eco14766, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14767(w_eco14767, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14768(w_eco14768, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14769(w_eco14769, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14770(w_eco14770, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14771(w_eco14771, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14772(w_eco14772, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14773(w_eco14773, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14774(w_eco14774, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14775(w_eco14775, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14776(w_eco14776, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14777(w_eco14777, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14778(w_eco14778, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14779(w_eco14779, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14780(w_eco14780, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14781(w_eco14781, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14782(w_eco14782, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14783(w_eco14783, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14784(w_eco14784, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14785(w_eco14785, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14786(w_eco14786, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14787(w_eco14787, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14788(w_eco14788, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14789(w_eco14789, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14790(w_eco14790, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_14791(w_eco14791, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14792(w_eco14792, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14793(w_eco14793, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14794(w_eco14794, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14795(w_eco14795, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14796(w_eco14796, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14797(w_eco14797, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14798(w_eco14798, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14799(w_eco14799, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14800(w_eco14800, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14801(w_eco14801, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14802(w_eco14802, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14803(w_eco14803, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_14804(w_eco14804, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14805(w_eco14805, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14806(w_eco14806, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14807(w_eco14807, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14808(w_eco14808, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_14809(w_eco14809, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14810(w_eco14810, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14811(w_eco14811, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14812(w_eco14812, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14813(w_eco14813, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14814(w_eco14814, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14815(w_eco14815, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14816(w_eco14816, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14817(w_eco14817, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14818(w_eco14818, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14819(w_eco14819, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14820(w_eco14820, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14821(w_eco14821, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14822(w_eco14822, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14823(w_eco14823, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14824(w_eco14824, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14825(w_eco14825, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14826(w_eco14826, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14827(w_eco14827, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14828(w_eco14828, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14829(w_eco14829, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14830(w_eco14830, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14831(w_eco14831, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14832(w_eco14832, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14833(w_eco14833, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14834(w_eco14834, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14835(w_eco14835, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14836(w_eco14836, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14837(w_eco14837, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14838(w_eco14838, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14839(w_eco14839, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14840(w_eco14840, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14841(w_eco14841, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14842(w_eco14842, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_14843(w_eco14843, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14844(w_eco14844, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14845(w_eco14845, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_14846(w_eco14846, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_14847(w_eco14847, w_eco14564, w_eco14565, w_eco14566, w_eco14567, w_eco14568, w_eco14569, w_eco14570, w_eco14571, w_eco14572, w_eco14573, w_eco14574, w_eco14575, w_eco14576, w_eco14577, w_eco14578, w_eco14579, w_eco14580, w_eco14581, w_eco14582, w_eco14583, w_eco14584, w_eco14585, w_eco14586, w_eco14587, w_eco14588, w_eco14589, w_eco14590, w_eco14591, w_eco14592, w_eco14593, w_eco14594, w_eco14595, w_eco14596, w_eco14597, w_eco14598, w_eco14599, w_eco14600, w_eco14601, w_eco14602, w_eco14603, w_eco14604, w_eco14605, w_eco14606, w_eco14607, w_eco14608, w_eco14609, w_eco14610, w_eco14611, w_eco14612, w_eco14613, w_eco14614, w_eco14615, w_eco14616, w_eco14617, w_eco14618, w_eco14619, w_eco14620, w_eco14621, w_eco14622, w_eco14623, w_eco14624, w_eco14625, w_eco14626, w_eco14627, w_eco14628, w_eco14629, w_eco14630, w_eco14631, w_eco14632, w_eco14633, w_eco14634, w_eco14635, w_eco14636, w_eco14637, w_eco14638, w_eco14639, w_eco14640, w_eco14641, w_eco14642, w_eco14643, w_eco14644, w_eco14645, w_eco14646, w_eco14647, w_eco14648, w_eco14649, w_eco14650, w_eco14651, w_eco14652, w_eco14653, w_eco14654, w_eco14655, w_eco14656, w_eco14657, w_eco14658, w_eco14659, w_eco14660, w_eco14661, w_eco14662, w_eco14663, w_eco14664, w_eco14665, w_eco14666, w_eco14667, w_eco14668, w_eco14669, w_eco14670, w_eco14671, w_eco14672, w_eco14673, w_eco14674, w_eco14675, w_eco14676, w_eco14677, w_eco14678, w_eco14679, w_eco14680, w_eco14681, w_eco14682, w_eco14683, w_eco14684, w_eco14685, w_eco14686, w_eco14687, w_eco14688, w_eco14689, w_eco14690, w_eco14691, w_eco14692, w_eco14693, w_eco14694, w_eco14695, w_eco14696, w_eco14697, w_eco14698, w_eco14699, w_eco14700, w_eco14701, w_eco14702, w_eco14703, w_eco14704, w_eco14705, w_eco14706, w_eco14707, w_eco14708, w_eco14709, w_eco14710, w_eco14711, w_eco14712, w_eco14713, w_eco14714, w_eco14715, w_eco14716, w_eco14717, w_eco14718, w_eco14719, w_eco14720, w_eco14721, w_eco14722, w_eco14723, w_eco14724, w_eco14725, w_eco14726, w_eco14727, w_eco14728, w_eco14729, w_eco14730, w_eco14731, w_eco14732, w_eco14733, w_eco14734, w_eco14735, w_eco14736, w_eco14737, w_eco14738, w_eco14739, w_eco14740, w_eco14741, w_eco14742, w_eco14743, w_eco14744, w_eco14745, w_eco14746, w_eco14747, w_eco14748, w_eco14749, w_eco14750, w_eco14751, w_eco14752, w_eco14753, w_eco14754, w_eco14755, w_eco14756, w_eco14757, w_eco14758, w_eco14759, w_eco14760, w_eco14761, w_eco14762, w_eco14763, w_eco14764, w_eco14765, w_eco14766, w_eco14767, w_eco14768, w_eco14769, w_eco14770, w_eco14771, w_eco14772, w_eco14773, w_eco14774, w_eco14775, w_eco14776, w_eco14777, w_eco14778, w_eco14779, w_eco14780, w_eco14781, w_eco14782, w_eco14783, w_eco14784, w_eco14785, w_eco14786, w_eco14787, w_eco14788, w_eco14789, w_eco14790, w_eco14791, w_eco14792, w_eco14793, w_eco14794, w_eco14795, w_eco14796, w_eco14797, w_eco14798, w_eco14799, w_eco14800, w_eco14801, w_eco14802, w_eco14803, w_eco14804, w_eco14805, w_eco14806, w_eco14807, w_eco14808, w_eco14809, w_eco14810, w_eco14811, w_eco14812, w_eco14813, w_eco14814, w_eco14815, w_eco14816, w_eco14817, w_eco14818, w_eco14819, w_eco14820, w_eco14821, w_eco14822, w_eco14823, w_eco14824, w_eco14825, w_eco14826, w_eco14827, w_eco14828, w_eco14829, w_eco14830, w_eco14831, w_eco14832, w_eco14833, w_eco14834, w_eco14835, w_eco14836, w_eco14837, w_eco14838, w_eco14839, w_eco14840, w_eco14841, w_eco14842, w_eco14843, w_eco14844, w_eco14845, w_eco14846);
	xor _ECO_out14(cnt[11], sub_wire14, w_eco14847);
	and _ECO_14848(w_eco14848, prev_cnt[10], rst);
	and _ECO_14849(w_eco14849, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14850(w_eco14850, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14851(w_eco14851, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14852(w_eco14852, prev_cnt[9], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14853(w_eco14853, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14854(w_eco14854, prev_cnt[9], prev_cnt[10], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14855(w_eco14855, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14856(w_eco14856, prev_cnt[10], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14857(w_eco14857, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14858(w_eco14858, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14859(w_eco14859, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14860(w_eco14860, prev_cnt[6], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14861(w_eco14861, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14862(w_eco14862, prev_cnt[6], prev_cnt[10], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14863(w_eco14863, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14864(w_eco14864, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14865(w_eco14865, prev_cnt[9], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14866(w_eco14866, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14867(w_eco14867, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14868(w_eco14868, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14869(w_eco14869, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14870(w_eco14870, prev_cnt[8], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14871(w_eco14871, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14872(w_eco14872, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14873(w_eco14873, prev_cnt[8], prev_cnt[10], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14874(w_eco14874, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14875(w_eco14875, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14876(w_eco14876, prev_cnt[6], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14877(w_eco14877, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14878(w_eco14878, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14879(w_eco14879, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14880(w_eco14880, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14881(w_eco14881, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14882(w_eco14882, Tgate[10], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14883(w_eco14883, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14884(w_eco14884, Tgate[10], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14885(w_eco14885, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14886(w_eco14886, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14887(w_eco14887, prev_cnt[8], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14888(w_eco14888, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14889(w_eco14889, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14890(w_eco14890, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14891(w_eco14891, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14892(w_eco14892, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14893(w_eco14893, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14894(w_eco14894, Tgate[10], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14895(w_eco14895, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14896(w_eco14896, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14897(w_eco14897, Tgate[10], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14898(w_eco14898, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14899(w_eco14899, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14900(w_eco14900, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14901(w_eco14901, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14902(w_eco14902, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14903(w_eco14903, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14904(w_eco14904, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14905(w_eco14905, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14906(w_eco14906, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14907(w_eco14907, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14908(w_eco14908, Tgate[10], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14909(w_eco14909, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_14910(w_eco14910, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14911(w_eco14911, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14912(w_eco14912, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14913(w_eco14913, Tgate[10], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14914(w_eco14914, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_14915(w_eco14915, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14916(w_eco14916, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14917(w_eco14917, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14918(w_eco14918, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14919(w_eco14919, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !ena, !rst);
	and _ECO_14920(w_eco14920, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14921(w_eco14921, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14922(w_eco14922, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14923(w_eco14923, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14924(w_eco14924, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14925(w_eco14925, Tgate[10], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14926(w_eco14926, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14927(w_eco14927, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14928(w_eco14928, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14929(w_eco14929, Tgate[10], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14930(w_eco14930, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14931(w_eco14931, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_state[0]);
	and _ECO_14932(w_eco14932, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14933(w_eco14933, Tgate[10], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_14934(w_eco14934, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14935(w_eco14935, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[3], prev_state[0]);
	and _ECO_14936(w_eco14936, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14937(w_eco14937, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14938(w_eco14938, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14939(w_eco14939, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14940(w_eco14940, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14941(w_eco14941, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14942(w_eco14942, Tgate[10], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14943(w_eco14943, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14944(w_eco14944, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14945(w_eco14945, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14946(w_eco14946, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14947(w_eco14947, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14948(w_eco14948, Tgate[10], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14949(w_eco14949, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_14950(w_eco14950, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_14951(w_eco14951, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_14952(w_eco14952, Tgate[10], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_14953(w_eco14953, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14954(w_eco14954, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14955(w_eco14955, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14956(w_eco14956, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[0]);
	and _ECO_14957(w_eco14957, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_14958(w_eco14958, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14959(w_eco14959, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14960(w_eco14960, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14961(w_eco14961, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14962(w_eco14962, Tgate[10], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14963(w_eco14963, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_14964(w_eco14964, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14965(w_eco14965, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14966(w_eco14966, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14967(w_eco14967, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14968(w_eco14968, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14969(w_eco14969, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14970(w_eco14970, Tgate[10], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14971(w_eco14971, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_14972(w_eco14972, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14973(w_eco14973, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_14974(w_eco14974, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14975(w_eco14975, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14976(w_eco14976, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14977(w_eco14977, Tgate[10], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_14978(w_eco14978, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14979(w_eco14979, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14980(w_eco14980, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[10], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_14981(w_eco14981, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_14982(w_eco14982, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14983(w_eco14983, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14984(w_eco14984, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_14985(w_eco14985, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_14986(w_eco14986, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14987(w_eco14987, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_14988(w_eco14988, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_14989(w_eco14989, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_14990(w_eco14990, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_14991(w_eco14991, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_14992(w_eco14992, Tgate[10], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_14993(w_eco14993, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_14994(w_eco14994, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14995(w_eco14995, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_14996(w_eco14996, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_14997(w_eco14997, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_14998(w_eco14998, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_14999(w_eco14999, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15000(w_eco15000, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15001(w_eco15001, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15002(w_eco15002, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15003(w_eco15003, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15004(w_eco15004, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15005(w_eco15005, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15006(w_eco15006, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15007(w_eco15007, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15008(w_eco15008, Tgate[10], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15009(w_eco15009, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15010(w_eco15010, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15011(w_eco15011, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15012(w_eco15012, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_15013(w_eco15013, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15014(w_eco15014, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15015(w_eco15015, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15016(w_eco15016, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15017(w_eco15017, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15018(w_eco15018, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15019(w_eco15019, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15020(w_eco15020, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15021(w_eco15021, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15022(w_eco15022, Tgate[10], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15023(w_eco15023, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15024(w_eco15024, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15025(w_eco15025, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15026(w_eco15026, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15027(w_eco15027, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_15028(w_eco15028, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15029(w_eco15029, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15030(w_eco15030, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15031(w_eco15031, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15032(w_eco15032, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15033(w_eco15033, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15034(w_eco15034, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15035(w_eco15035, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15036(w_eco15036, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15037(w_eco15037, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15038(w_eco15038, Tgate[10], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15039(w_eco15039, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15040(w_eco15040, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15041(w_eco15041, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15042(w_eco15042, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15043(w_eco15043, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], prev_state[1]);
	and _ECO_15044(w_eco15044, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15045(w_eco15045, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15046(w_eco15046, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15047(w_eco15047, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15048(w_eco15048, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15049(w_eco15049, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15050(w_eco15050, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15051(w_eco15051, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15052(w_eco15052, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15053(w_eco15053, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15054(w_eco15054, Tgate[10], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15055(w_eco15055, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15056(w_eco15056, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15057(w_eco15057, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15058(w_eco15058, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15059(w_eco15059, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15060(w_eco15060, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15061(w_eco15061, Tgate[10], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15062(w_eco15062, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15063(w_eco15063, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15064(w_eco15064, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15065(w_eco15065, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15066(w_eco15066, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15067(w_eco15067, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15068(w_eco15068, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15069(w_eco15069, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15070(w_eco15070, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15071(w_eco15071, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15072(w_eco15072, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15073(w_eco15073, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15074(w_eco15074, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15075(w_eco15075, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15076(w_eco15076, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15077(w_eco15077, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15078(w_eco15078, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15079(w_eco15079, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15080(w_eco15080, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15081(w_eco15081, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15082(w_eco15082, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15083(w_eco15083, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15084(w_eco15084, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15085(w_eco15085, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15086(w_eco15086, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15087(w_eco15087, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15088(w_eco15088, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15089(w_eco15089, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15090(w_eco15090, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15091(w_eco15091, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15092(w_eco15092, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15093(w_eco15093, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15094(w_eco15094, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15095(w_eco15095, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15096(w_eco15096, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15097(w_eco15097, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15098(w_eco15098, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15099(w_eco15099, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15100(w_eco15100, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15101(w_eco15101, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15102(w_eco15102, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15103(w_eco15103, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15104(w_eco15104, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15105(w_eco15105, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15106(w_eco15106, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15107(w_eco15107, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15108(w_eco15108, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15109(w_eco15109, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15110(w_eco15110, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15111(w_eco15111, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15112(w_eco15112, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15113(w_eco15113, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15114(w_eco15114, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15115(w_eco15115, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15116(w_eco15116, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15117(w_eco15117, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15118(w_eco15118, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15119(w_eco15119, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15120(w_eco15120, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15121(w_eco15121, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15122(w_eco15122, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15123(w_eco15123, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15124(w_eco15124, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15125(w_eco15125, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15126(w_eco15126, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15127(w_eco15127, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15128(w_eco15128, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15129(w_eco15129, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15130(w_eco15130, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15131(w_eco15131, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15132(w_eco15132, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15133(w_eco15133, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15134(w_eco15134, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15135(w_eco15135, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15136(w_eco15136, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15137(w_eco15137, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15138(w_eco15138, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15139(w_eco15139, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15140(w_eco15140, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15141(w_eco15141, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15142(w_eco15142, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15143(w_eco15143, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15144(w_eco15144, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15145(w_eco15145, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15146(w_eco15146, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15147(w_eco15147, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15148(w_eco15148, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15149(w_eco15149, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15150(w_eco15150, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15151(w_eco15151, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15152(w_eco15152, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15153(w_eco15153, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15154(w_eco15154, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15155(w_eco15155, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_15156(w_eco15156, w_eco14848, w_eco14849, w_eco14850, w_eco14851, w_eco14852, w_eco14853, w_eco14854, w_eco14855, w_eco14856, w_eco14857, w_eco14858, w_eco14859, w_eco14860, w_eco14861, w_eco14862, w_eco14863, w_eco14864, w_eco14865, w_eco14866, w_eco14867, w_eco14868, w_eco14869, w_eco14870, w_eco14871, w_eco14872, w_eco14873, w_eco14874, w_eco14875, w_eco14876, w_eco14877, w_eco14878, w_eco14879, w_eco14880, w_eco14881, w_eco14882, w_eco14883, w_eco14884, w_eco14885, w_eco14886, w_eco14887, w_eco14888, w_eco14889, w_eco14890, w_eco14891, w_eco14892, w_eco14893, w_eco14894, w_eco14895, w_eco14896, w_eco14897, w_eco14898, w_eco14899, w_eco14900, w_eco14901, w_eco14902, w_eco14903, w_eco14904, w_eco14905, w_eco14906, w_eco14907, w_eco14908, w_eco14909, w_eco14910, w_eco14911, w_eco14912, w_eco14913, w_eco14914, w_eco14915, w_eco14916, w_eco14917, w_eco14918, w_eco14919, w_eco14920, w_eco14921, w_eco14922, w_eco14923, w_eco14924, w_eco14925, w_eco14926, w_eco14927, w_eco14928, w_eco14929, w_eco14930, w_eco14931, w_eco14932, w_eco14933, w_eco14934, w_eco14935, w_eco14936, w_eco14937, w_eco14938, w_eco14939, w_eco14940, w_eco14941, w_eco14942, w_eco14943, w_eco14944, w_eco14945, w_eco14946, w_eco14947, w_eco14948, w_eco14949, w_eco14950, w_eco14951, w_eco14952, w_eco14953, w_eco14954, w_eco14955, w_eco14956, w_eco14957, w_eco14958, w_eco14959, w_eco14960, w_eco14961, w_eco14962, w_eco14963, w_eco14964, w_eco14965, w_eco14966, w_eco14967, w_eco14968, w_eco14969, w_eco14970, w_eco14971, w_eco14972, w_eco14973, w_eco14974, w_eco14975, w_eco14976, w_eco14977, w_eco14978, w_eco14979, w_eco14980, w_eco14981, w_eco14982, w_eco14983, w_eco14984, w_eco14985, w_eco14986, w_eco14987, w_eco14988, w_eco14989, w_eco14990, w_eco14991, w_eco14992, w_eco14993, w_eco14994, w_eco14995, w_eco14996, w_eco14997, w_eco14998, w_eco14999, w_eco15000, w_eco15001, w_eco15002, w_eco15003, w_eco15004, w_eco15005, w_eco15006, w_eco15007, w_eco15008, w_eco15009, w_eco15010, w_eco15011, w_eco15012, w_eco15013, w_eco15014, w_eco15015, w_eco15016, w_eco15017, w_eco15018, w_eco15019, w_eco15020, w_eco15021, w_eco15022, w_eco15023, w_eco15024, w_eco15025, w_eco15026, w_eco15027, w_eco15028, w_eco15029, w_eco15030, w_eco15031, w_eco15032, w_eco15033, w_eco15034, w_eco15035, w_eco15036, w_eco15037, w_eco15038, w_eco15039, w_eco15040, w_eco15041, w_eco15042, w_eco15043, w_eco15044, w_eco15045, w_eco15046, w_eco15047, w_eco15048, w_eco15049, w_eco15050, w_eco15051, w_eco15052, w_eco15053, w_eco15054, w_eco15055, w_eco15056, w_eco15057, w_eco15058, w_eco15059, w_eco15060, w_eco15061, w_eco15062, w_eco15063, w_eco15064, w_eco15065, w_eco15066, w_eco15067, w_eco15068, w_eco15069, w_eco15070, w_eco15071, w_eco15072, w_eco15073, w_eco15074, w_eco15075, w_eco15076, w_eco15077, w_eco15078, w_eco15079, w_eco15080, w_eco15081, w_eco15082, w_eco15083, w_eco15084, w_eco15085, w_eco15086, w_eco15087, w_eco15088, w_eco15089, w_eco15090, w_eco15091, w_eco15092, w_eco15093, w_eco15094, w_eco15095, w_eco15096, w_eco15097, w_eco15098, w_eco15099, w_eco15100, w_eco15101, w_eco15102, w_eco15103, w_eco15104, w_eco15105, w_eco15106, w_eco15107, w_eco15108, w_eco15109, w_eco15110, w_eco15111, w_eco15112, w_eco15113, w_eco15114, w_eco15115, w_eco15116, w_eco15117, w_eco15118, w_eco15119, w_eco15120, w_eco15121, w_eco15122, w_eco15123, w_eco15124, w_eco15125, w_eco15126, w_eco15127, w_eco15128, w_eco15129, w_eco15130, w_eco15131, w_eco15132, w_eco15133, w_eco15134, w_eco15135, w_eco15136, w_eco15137, w_eco15138, w_eco15139, w_eco15140, w_eco15141, w_eco15142, w_eco15143, w_eco15144, w_eco15145, w_eco15146, w_eco15147, w_eco15148, w_eco15149, w_eco15150, w_eco15151, w_eco15152, w_eco15153, w_eco15154, w_eco15155);
	xor _ECO_out15(cnt[10], sub_wire15, w_eco15156);
	and _ECO_15157(w_eco15157, prev_cnt[9], rst);
	and _ECO_15158(w_eco15158, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15159(w_eco15159, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15160(w_eco15160, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15161(w_eco15161, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15162(w_eco15162, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15163(w_eco15163, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15164(w_eco15164, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15165(w_eco15165, prev_cnt[6], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_15166(w_eco15166, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15167(w_eco15167, prev_cnt[6], prev_cnt[9], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_15168(w_eco15168, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15169(w_eco15169, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15170(w_eco15170, prev_cnt[9], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15171(w_eco15171, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15172(w_eco15172, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15173(w_eco15173, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15174(w_eco15174, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15175(w_eco15175, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15176(w_eco15176, prev_cnt[8], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_15177(w_eco15177, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15178(w_eco15178, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15179(w_eco15179, prev_cnt[8], prev_cnt[9], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_15180(w_eco15180, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15181(w_eco15181, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15182(w_eco15182, prev_cnt[6], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15183(w_eco15183, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15184(w_eco15184, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15185(w_eco15185, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15186(w_eco15186, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15187(w_eco15187, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15188(w_eco15188, Tgate[9], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15189(w_eco15189, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15190(w_eco15190, Tgate[9], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15191(w_eco15191, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15192(w_eco15192, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15193(w_eco15193, prev_cnt[8], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15194(w_eco15194, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15195(w_eco15195, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15196(w_eco15196, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15197(w_eco15197, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15198(w_eco15198, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15199(w_eco15199, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15200(w_eco15200, Tgate[9], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15201(w_eco15201, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15202(w_eco15202, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15203(w_eco15203, Tgate[9], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15204(w_eco15204, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15205(w_eco15205, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15206(w_eco15206, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15207(w_eco15207, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15208(w_eco15208, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !ena, !rst);
	and _ECO_15209(w_eco15209, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15210(w_eco15210, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15211(w_eco15211, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15212(w_eco15212, Tgate[9], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15213(w_eco15213, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15214(w_eco15214, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15215(w_eco15215, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15216(w_eco15216, Tgate[9], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15217(w_eco15217, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15218(w_eco15218, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15219(w_eco15219, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15220(w_eco15220, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15221(w_eco15221, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15222(w_eco15222, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15223(w_eco15223, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !ena, !rst);
	and _ECO_15224(w_eco15224, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15225(w_eco15225, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15226(w_eco15226, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15227(w_eco15227, Tgate[9], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15228(w_eco15228, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15229(w_eco15229, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15230(w_eco15230, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15231(w_eco15231, Tgate[9], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15232(w_eco15232, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15233(w_eco15233, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15234(w_eco15234, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15235(w_eco15235, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_state[0]);
	and _ECO_15236(w_eco15236, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15237(w_eco15237, Tgate[9], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15238(w_eco15238, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15239(w_eco15239, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15240(w_eco15240, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15241(w_eco15241, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15242(w_eco15242, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15243(w_eco15243, Tgate[9], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15244(w_eco15244, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15245(w_eco15245, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15246(w_eco15246, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15247(w_eco15247, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15248(w_eco15248, Tgate[9], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15249(w_eco15249, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15250(w_eco15250, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15251(w_eco15251, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15252(w_eco15252, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15253(w_eco15253, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15254(w_eco15254, Tgate[9], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15255(w_eco15255, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15256(w_eco15256, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15257(w_eco15257, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15258(w_eco15258, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[0]);
	and _ECO_15259(w_eco15259, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_15260(w_eco15260, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15261(w_eco15261, Tgate[9], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15262(w_eco15262, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15263(w_eco15263, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15264(w_eco15264, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15265(w_eco15265, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_15266(w_eco15266, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15267(w_eco15267, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15268(w_eco15268, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15269(w_eco15269, Tgate[9], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15270(w_eco15270, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15271(w_eco15271, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15272(w_eco15272, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15273(w_eco15273, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15274(w_eco15274, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15275(w_eco15275, Tgate[9], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15276(w_eco15276, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15277(w_eco15277, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15278(w_eco15278, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15279(w_eco15279, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15280(w_eco15280, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15281(w_eco15281, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15282(w_eco15282, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15283(w_eco15283, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15284(w_eco15284, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15285(w_eco15285, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15286(w_eco15286, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15287(w_eco15287, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15288(w_eco15288, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15289(w_eco15289, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15290(w_eco15290, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15291(w_eco15291, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15292(w_eco15292, Tgate[9], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15293(w_eco15293, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[9], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15294(w_eco15294, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15295(w_eco15295, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15296(w_eco15296, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15297(w_eco15297, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15298(w_eco15298, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15299(w_eco15299, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15300(w_eco15300, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15301(w_eco15301, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15302(w_eco15302, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15303(w_eco15303, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15304(w_eco15304, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15305(w_eco15305, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15306(w_eco15306, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15307(w_eco15307, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15308(w_eco15308, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15309(w_eco15309, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15310(w_eco15310, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15311(w_eco15311, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15312(w_eco15312, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15313(w_eco15313, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15314(w_eco15314, Tgate[9], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15315(w_eco15315, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15316(w_eco15316, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15317(w_eco15317, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15318(w_eco15318, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15319(w_eco15319, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15320(w_eco15320, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15321(w_eco15321, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15322(w_eco15322, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15323(w_eco15323, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15324(w_eco15324, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15325(w_eco15325, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15326(w_eco15326, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15327(w_eco15327, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15328(w_eco15328, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15329(w_eco15329, Tgate[9], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15330(w_eco15330, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15331(w_eco15331, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15332(w_eco15332, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15333(w_eco15333, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15334(w_eco15334, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15335(w_eco15335, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15336(w_eco15336, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15337(w_eco15337, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15338(w_eco15338, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15339(w_eco15339, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15340(w_eco15340, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15341(w_eco15341, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15342(w_eco15342, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15343(w_eco15343, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15344(w_eco15344, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15345(w_eco15345, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15346(w_eco15346, Tgate[9], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15347(w_eco15347, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15348(w_eco15348, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15349(w_eco15349, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15350(w_eco15350, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15351(w_eco15351, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15352(w_eco15352, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15353(w_eco15353, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[9], prev_state[1]);
	and _ECO_15354(w_eco15354, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15355(w_eco15355, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15356(w_eco15356, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15357(w_eco15357, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15358(w_eco15358, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15359(w_eco15359, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15360(w_eco15360, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15361(w_eco15361, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15362(w_eco15362, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15363(w_eco15363, Tgate[9], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15364(w_eco15364, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15365(w_eco15365, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15366(w_eco15366, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15367(w_eco15367, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15368(w_eco15368, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15369(w_eco15369, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15370(w_eco15370, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15371(w_eco15371, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15372(w_eco15372, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15373(w_eco15373, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15374(w_eco15374, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15375(w_eco15375, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15376(w_eco15376, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15377(w_eco15377, Tgate[9], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1]);
	and _ECO_15378(w_eco15378, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15379(w_eco15379, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15380(w_eco15380, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15381(w_eco15381, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15382(w_eco15382, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15383(w_eco15383, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15384(w_eco15384, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15385(w_eco15385, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15386(w_eco15386, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15387(w_eco15387, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15388(w_eco15388, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15389(w_eco15389, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15390(w_eco15390, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15391(w_eco15391, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15392(w_eco15392, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15393(w_eco15393, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15394(w_eco15394, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15395(w_eco15395, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15396(w_eco15396, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15397(w_eco15397, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15398(w_eco15398, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15399(w_eco15399, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15400(w_eco15400, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15401(w_eco15401, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15402(w_eco15402, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15403(w_eco15403, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15404(w_eco15404, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15405(w_eco15405, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15406(w_eco15406, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15407(w_eco15407, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15408(w_eco15408, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15409(w_eco15409, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15410(w_eco15410, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15411(w_eco15411, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15412(w_eco15412, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15413(w_eco15413, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15414(w_eco15414, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15415(w_eco15415, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15416(w_eco15416, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15417(w_eco15417, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15418(w_eco15418, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15419(w_eco15419, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15420(w_eco15420, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15421(w_eco15421, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15422(w_eco15422, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15423(w_eco15423, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15424(w_eco15424, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15425(w_eco15425, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15426(w_eco15426, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15427(w_eco15427, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15428(w_eco15428, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15429(w_eco15429, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15430(w_eco15430, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15431(w_eco15431, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15432(w_eco15432, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15433(w_eco15433, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15434(w_eco15434, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15435(w_eco15435, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15436(w_eco15436, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15437(w_eco15437, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15438(w_eco15438, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15439(w_eco15439, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15440(w_eco15440, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15441(w_eco15441, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15442(w_eco15442, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15443(w_eco15443, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15444(w_eco15444, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15445(w_eco15445, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15446(w_eco15446, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15447(w_eco15447, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15448(w_eco15448, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15449(w_eco15449, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15450(w_eco15450, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15451(w_eco15451, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15452(w_eco15452, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15453(w_eco15453, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15454(w_eco15454, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15455(w_eco15455, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15456(w_eco15456, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15457(w_eco15457, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15458(w_eco15458, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15459(w_eco15459, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15460(w_eco15460, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15461(w_eco15461, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15462(w_eco15462, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15463(w_eco15463, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15464(w_eco15464, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15465(w_eco15465, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15466(w_eco15466, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15467(w_eco15467, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15468(w_eco15468, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15469(w_eco15469, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15470(w_eco15470, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15471(w_eco15471, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15472(w_eco15472, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15473(w_eco15473, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15474(w_eco15474, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15475(w_eco15475, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15476(w_eco15476, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15477(w_eco15477, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15478(w_eco15478, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15479(w_eco15479, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15480(w_eco15480, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15481(w_eco15481, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15482(w_eco15482, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_15483(w_eco15483, w_eco15157, w_eco15158, w_eco15159, w_eco15160, w_eco15161, w_eco15162, w_eco15163, w_eco15164, w_eco15165, w_eco15166, w_eco15167, w_eco15168, w_eco15169, w_eco15170, w_eco15171, w_eco15172, w_eco15173, w_eco15174, w_eco15175, w_eco15176, w_eco15177, w_eco15178, w_eco15179, w_eco15180, w_eco15181, w_eco15182, w_eco15183, w_eco15184, w_eco15185, w_eco15186, w_eco15187, w_eco15188, w_eco15189, w_eco15190, w_eco15191, w_eco15192, w_eco15193, w_eco15194, w_eco15195, w_eco15196, w_eco15197, w_eco15198, w_eco15199, w_eco15200, w_eco15201, w_eco15202, w_eco15203, w_eco15204, w_eco15205, w_eco15206, w_eco15207, w_eco15208, w_eco15209, w_eco15210, w_eco15211, w_eco15212, w_eco15213, w_eco15214, w_eco15215, w_eco15216, w_eco15217, w_eco15218, w_eco15219, w_eco15220, w_eco15221, w_eco15222, w_eco15223, w_eco15224, w_eco15225, w_eco15226, w_eco15227, w_eco15228, w_eco15229, w_eco15230, w_eco15231, w_eco15232, w_eco15233, w_eco15234, w_eco15235, w_eco15236, w_eco15237, w_eco15238, w_eco15239, w_eco15240, w_eco15241, w_eco15242, w_eco15243, w_eco15244, w_eco15245, w_eco15246, w_eco15247, w_eco15248, w_eco15249, w_eco15250, w_eco15251, w_eco15252, w_eco15253, w_eco15254, w_eco15255, w_eco15256, w_eco15257, w_eco15258, w_eco15259, w_eco15260, w_eco15261, w_eco15262, w_eco15263, w_eco15264, w_eco15265, w_eco15266, w_eco15267, w_eco15268, w_eco15269, w_eco15270, w_eco15271, w_eco15272, w_eco15273, w_eco15274, w_eco15275, w_eco15276, w_eco15277, w_eco15278, w_eco15279, w_eco15280, w_eco15281, w_eco15282, w_eco15283, w_eco15284, w_eco15285, w_eco15286, w_eco15287, w_eco15288, w_eco15289, w_eco15290, w_eco15291, w_eco15292, w_eco15293, w_eco15294, w_eco15295, w_eco15296, w_eco15297, w_eco15298, w_eco15299, w_eco15300, w_eco15301, w_eco15302, w_eco15303, w_eco15304, w_eco15305, w_eco15306, w_eco15307, w_eco15308, w_eco15309, w_eco15310, w_eco15311, w_eco15312, w_eco15313, w_eco15314, w_eco15315, w_eco15316, w_eco15317, w_eco15318, w_eco15319, w_eco15320, w_eco15321, w_eco15322, w_eco15323, w_eco15324, w_eco15325, w_eco15326, w_eco15327, w_eco15328, w_eco15329, w_eco15330, w_eco15331, w_eco15332, w_eco15333, w_eco15334, w_eco15335, w_eco15336, w_eco15337, w_eco15338, w_eco15339, w_eco15340, w_eco15341, w_eco15342, w_eco15343, w_eco15344, w_eco15345, w_eco15346, w_eco15347, w_eco15348, w_eco15349, w_eco15350, w_eco15351, w_eco15352, w_eco15353, w_eco15354, w_eco15355, w_eco15356, w_eco15357, w_eco15358, w_eco15359, w_eco15360, w_eco15361, w_eco15362, w_eco15363, w_eco15364, w_eco15365, w_eco15366, w_eco15367, w_eco15368, w_eco15369, w_eco15370, w_eco15371, w_eco15372, w_eco15373, w_eco15374, w_eco15375, w_eco15376, w_eco15377, w_eco15378, w_eco15379, w_eco15380, w_eco15381, w_eco15382, w_eco15383, w_eco15384, w_eco15385, w_eco15386, w_eco15387, w_eco15388, w_eco15389, w_eco15390, w_eco15391, w_eco15392, w_eco15393, w_eco15394, w_eco15395, w_eco15396, w_eco15397, w_eco15398, w_eco15399, w_eco15400, w_eco15401, w_eco15402, w_eco15403, w_eco15404, w_eco15405, w_eco15406, w_eco15407, w_eco15408, w_eco15409, w_eco15410, w_eco15411, w_eco15412, w_eco15413, w_eco15414, w_eco15415, w_eco15416, w_eco15417, w_eco15418, w_eco15419, w_eco15420, w_eco15421, w_eco15422, w_eco15423, w_eco15424, w_eco15425, w_eco15426, w_eco15427, w_eco15428, w_eco15429, w_eco15430, w_eco15431, w_eco15432, w_eco15433, w_eco15434, w_eco15435, w_eco15436, w_eco15437, w_eco15438, w_eco15439, w_eco15440, w_eco15441, w_eco15442, w_eco15443, w_eco15444, w_eco15445, w_eco15446, w_eco15447, w_eco15448, w_eco15449, w_eco15450, w_eco15451, w_eco15452, w_eco15453, w_eco15454, w_eco15455, w_eco15456, w_eco15457, w_eco15458, w_eco15459, w_eco15460, w_eco15461, w_eco15462, w_eco15463, w_eco15464, w_eco15465, w_eco15466, w_eco15467, w_eco15468, w_eco15469, w_eco15470, w_eco15471, w_eco15472, w_eco15473, w_eco15474, w_eco15475, w_eco15476, w_eco15477, w_eco15478, w_eco15479, w_eco15480, w_eco15481, w_eco15482);
	xor _ECO_out16(cnt[9], sub_wire16, w_eco15483);
	and _ECO_15484(w_eco15484, prev_cnt[8], rst);
	and _ECO_15485(w_eco15485, prev_cnt[1], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15486(w_eco15486, prev_cnt[1], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15487(w_eco15487, prev_cnt[1], !prev_cnt[6], !ena, !rst);
	and _ECO_15488(w_eco15488, prev_cnt[2], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15489(w_eco15489, prev_cnt[2], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15490(w_eco15490, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15491(w_eco15491, prev_cnt[2], !prev_cnt[6], !ena, !rst);
	and _ECO_15492(w_eco15492, prev_cnt[3], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15493(w_eco15493, prev_cnt[3], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15494(w_eco15494, prev_cnt[1], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15495(w_eco15495, prev_cnt[1], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15496(w_eco15496, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15497(w_eco15497, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15498(w_eco15498, prev_cnt[3], !prev_cnt[6], !ena, !rst);
	and _ECO_15499(w_eco15499, prev_cnt[6], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_15500(w_eco15500, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15501(w_eco15501, prev_cnt[0], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15502(w_eco15502, prev_cnt[6], prev_cnt[8], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_15503(w_eco15503, prev_cnt[0], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15504(w_eco15504, prev_cnt[2], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15505(w_eco15505, prev_cnt[8], ena, !prev_state[4], !prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15506(w_eco15506, prev_cnt[2], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15507(w_eco15507, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15508(w_eco15508, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15509(w_eco15509, prev_cnt[0], !prev_cnt[6], !ena, !rst);
	and _ECO_15510(w_eco15510, prev_cnt[3], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15511(w_eco15511, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15512(w_eco15512, Tgate[8], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15513(w_eco15513, prev_cnt[4], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15514(w_eco15514, Tgate[8], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15515(w_eco15515, prev_cnt[4], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15516(w_eco15516, prev_cnt[3], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15517(w_eco15517, prev_cnt[6], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15518(w_eco15518, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15519(w_eco15519, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15520(w_eco15520, prev_cnt[4], !prev_cnt[6], !ena, !rst);
	and _ECO_15521(w_eco15521, prev_cnt[0], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15522(w_eco15522, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15523(w_eco15523, Tgate[8], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15524(w_eco15524, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15525(w_eco15525, prev_cnt[5], !prev_cnt[6], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15526(w_eco15526, Tgate[8], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15527(w_eco15527, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15528(w_eco15528, prev_cnt[5], !prev_cnt[6], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15529(w_eco15529, prev_cnt[0], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15530(w_eco15530, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15531(w_eco15531, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15532(w_eco15532, prev_cnt[5], !prev_cnt[6], !ena, !rst);
	and _ECO_15533(w_eco15533, prev_cnt[4], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15534(w_eco15534, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15535(w_eco15535, Tgate[8], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15536(w_eco15536, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15537(w_eco15537, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15538(w_eco15538, !prev_cnt[6], prev_cnt[7], !rst, prev_state[4], !prev_state[2], prev_state[1]);
	and _ECO_15539(w_eco15539, Tgate[8], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15540(w_eco15540, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15541(w_eco15541, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15542(w_eco15542, !prev_cnt[6], prev_cnt[7], !rst, prev_state[3], !prev_state[2], prev_state[1]);
	and _ECO_15543(w_eco15543, prev_cnt[4], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15544(w_eco15544, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_state[0]);
	and _ECO_15545(w_eco15545, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15546(w_eco15546, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15547(w_eco15547, !prev_cnt[6], prev_cnt[7], !ena, !rst);
	and _ECO_15548(w_eco15548, prev_cnt[5], !prev_cnt[6], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15549(w_eco15549, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15550(w_eco15550, Tgate[8], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15551(w_eco15551, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15552(w_eco15552, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15553(w_eco15553, Tgate[8], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15554(w_eco15554, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15555(w_eco15555, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15556(w_eco15556, prev_cnt[5], !prev_cnt[6], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15557(w_eco15557, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_state[0]);
	and _ECO_15558(w_eco15558, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15559(w_eco15559, Tgate[8], prev_cnt[1], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15560(w_eco15560, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15561(w_eco15561, !prev_cnt[6], prev_cnt[7], !rst, !prev_state[3], prev_state[0]);
	and _ECO_15562(w_eco15562, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15563(w_eco15563, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15564(w_eco15564, Tgate[8], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15565(w_eco15565, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15566(w_eco15566, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15567(w_eco15567, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15568(w_eco15568, prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15569(w_eco15569, Tgate[8], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15570(w_eco15570, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15571(w_eco15571, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15572(w_eco15572, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15573(w_eco15573, !prev_cnt[6], prev_cnt[7], !rst, !prev_state[4], !prev_state[2], prev_state[0]);
	and _ECO_15574(w_eco15574, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[0]);
	and _ECO_15575(w_eco15575, Tgate[8], prev_cnt[2], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15576(w_eco15576, prev_cnt[1], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15577(w_eco15577, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15578(w_eco15578, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15579(w_eco15579, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[0]);
	and _ECO_15580(w_eco15580, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[3], prev_state[2], !prev_state[1]);
	and _ECO_15581(w_eco15581, Tgate[8], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15582(w_eco15582, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15583(w_eco15583, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15584(w_eco15584, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15585(w_eco15585, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15586(w_eco15586, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[3], !prev_state[1], prev_state[0]);
	and _ECO_15587(w_eco15587, prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15588(w_eco15588, Tgate[8], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15589(w_eco15589, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15590(w_eco15590, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15591(w_eco15591, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15592(w_eco15592, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15593(w_eco15593, Tgate[8], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[3], prev_state[2]);
	and _ECO_15594(w_eco15594, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15595(w_eco15595, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15596(w_eco15596, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15597(w_eco15597, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15598(w_eco15598, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15599(w_eco15599, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15600(w_eco15600, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15601(w_eco15601, prev_cnt[3], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15602(w_eco15602, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15603(w_eco15603, prev_cnt[1], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15604(w_eco15604, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15605(w_eco15605, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15606(w_eco15606, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15607(w_eco15607, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15608(w_eco15608, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[11], !rst, prev_state[3], prev_state[2]);
	and _ECO_15609(w_eco15609, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15610(w_eco15610, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15611(w_eco15611, Tgate[8], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !rst, prev_state[4], prev_state[2]);
	and _ECO_15612(w_eco15612, !prev_cnt[0], !prev_cnt[1], !prev_cnt[2], !prev_cnt[3], !prev_cnt[4], !prev_cnt[5], !prev_cnt[7], prev_cnt[8], ena, prev_state[4], prev_state[2], !prev_state[1], !prev_state[0]);
	and _ECO_15613(w_eco15613, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15614(w_eco15614, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15615(w_eco15615, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15616(w_eco15616, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15617(w_eco15617, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15618(w_eco15618, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15619(w_eco15619, prev_cnt[1], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15620(w_eco15620, prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15621(w_eco15621, prev_cnt[0], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15622(w_eco15622, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15623(w_eco15623, prev_cnt[2], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15624(w_eco15624, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15625(w_eco15625, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15626(w_eco15626, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15627(w_eco15627, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[15], !rst, prev_state[3], prev_state[2]);
	and _ECO_15628(w_eco15628, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15629(w_eco15629, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15630(w_eco15630, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15631(w_eco15631, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15632(w_eco15632, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15633(w_eco15633, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15634(w_eco15634, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15635(w_eco15635, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[11], !rst, prev_state[4], prev_state[2]);
	and _ECO_15636(w_eco15636, Tgate[8], prev_cnt[3], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15637(w_eco15637, prev_cnt[1], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15638(w_eco15638, prev_cnt[2], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15639(w_eco15639, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15640(w_eco15640, prev_cnt[2], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15641(w_eco15641, prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15642(w_eco15642, prev_cnt[4], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15643(w_eco15643, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15644(w_eco15644, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15645(w_eco15645, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15646(w_eco15646, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15647(w_eco15647, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15648(w_eco15648, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15649(w_eco15649, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15650(w_eco15650, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15651(w_eco15651, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15652(w_eco15652, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15653(w_eco15653, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[15], !rst, prev_state[4], prev_state[2]);
	and _ECO_15654(w_eco15654, Tgate[8], prev_cnt[0], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15655(w_eco15655, prev_cnt[2], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15656(w_eco15656, prev_cnt[3], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15657(w_eco15657, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15658(w_eco15658, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15659(w_eco15659, prev_cnt[3], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15660(w_eco15660, prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15661(w_eco15661, prev_cnt[5], !prev_cnt[6], prev_cnt[8], prev_state[1]);
	and _ECO_15662(w_eco15662, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15663(w_eco15663, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15664(w_eco15664, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15665(w_eco15665, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[9], !rst, prev_state[3], prev_state[2]);
	and _ECO_15666(w_eco15666, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15667(w_eco15667, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15668(w_eco15668, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15669(w_eco15669, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15670(w_eco15670, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15671(w_eco15671, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15672(w_eco15672, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15673(w_eco15673, Tgate[8], prev_cnt[4], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15674(w_eco15674, prev_cnt[1], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15675(w_eco15675, prev_cnt[3], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15676(w_eco15676, prev_cnt[0], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15677(w_eco15677, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15678(w_eco15678, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15679(w_eco15679, prev_cnt[0], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15680(w_eco15680, prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15681(w_eco15681, !prev_cnt[6], prev_cnt[7], prev_cnt[8], prev_state[1]);
	and _ECO_15682(w_eco15682, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15683(w_eco15683, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15684(w_eco15684, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[10], !rst, prev_state[3], prev_state[2]);
	and _ECO_15685(w_eco15685, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15686(w_eco15686, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15687(w_eco15687, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15688(w_eco15688, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15689(w_eco15689, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[9], !rst, prev_state[4], prev_state[2]);
	and _ECO_15690(w_eco15690, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15691(w_eco15691, Tgate[8], prev_cnt[5], !prev_cnt[6], !rst, prev_state[1]);
	and _ECO_15692(w_eco15692, prev_cnt[1], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15693(w_eco15693, prev_cnt[2], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15694(w_eco15694, prev_cnt[0], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15695(w_eco15695, prev_cnt[4], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15696(w_eco15696, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15697(w_eco15697, prev_cnt[4], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15698(w_eco15698, prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15699(w_eco15699, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15700(w_eco15700, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15701(w_eco15701, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[12], !rst, prev_state[3], prev_state[2]);
	and _ECO_15702(w_eco15702, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[2], !prev_state[1]);
	and _ECO_15703(w_eco15703, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15704(w_eco15704, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15705(w_eco15705, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[10], !rst, prev_state[4], prev_state[2]);
	and _ECO_15706(w_eco15706, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15707(w_eco15707, Tgate[8], !prev_cnt[6], prev_cnt[7], !rst, prev_state[1]);
	and _ECO_15708(w_eco15708, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15709(w_eco15709, prev_cnt[2], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15710(w_eco15710, prev_cnt[3], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15711(w_eco15711, prev_cnt[4], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15712(w_eco15712, prev_cnt[5], !prev_cnt[6], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15713(w_eco15713, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15714(w_eco15714, prev_cnt[5], !prev_cnt[6], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15715(w_eco15715, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15716(w_eco15716, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15717(w_eco15717, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15718(w_eco15718, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[13], !rst, prev_state[3], prev_state[2]);
	and _ECO_15719(w_eco15719, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15720(w_eco15720, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[12], !rst, prev_state[4], prev_state[2]);
	and _ECO_15721(w_eco15721, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15722(w_eco15722, !prev_cnt[14], prev_cnt[1], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15723(w_eco15723, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15724(w_eco15724, prev_cnt[3], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15725(w_eco15725, prev_cnt[0], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15726(w_eco15726, prev_cnt[5], !prev_cnt[6], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15727(w_eco15727, !prev_cnt[6], prev_cnt[7], prev_cnt[11], !rst, prev_state[1]);
	and _ECO_15728(w_eco15728, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15729(w_eco15729, !prev_cnt[6], prev_cnt[7], !prev_cnt[8], !prev_cnt[9], !prev_cnt[10], !prev_cnt[11], !prev_cnt[12], !prev_cnt[13], !prev_cnt[15], !rst, !prev_state[4], !prev_state[3], !prev_state[1]);
	and _ECO_15730(w_eco15730, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15731(w_eco15731, !prev_cnt[14], prev_cnt[2], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15732(w_eco15732, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15733(w_eco15733, prev_cnt[0], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15734(w_eco15734, prev_cnt[4], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15735(w_eco15735, !prev_cnt[6], prev_cnt[7], prev_cnt[15], !rst, prev_state[1]);
	and _ECO_15736(w_eco15736, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15737(w_eco15737, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15738(w_eco15738, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15739(w_eco15739, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15740(w_eco15740, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15741(w_eco15741, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15742(w_eco15742, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], !prev_cnt[8], prev_cnt[13], !rst, prev_state[4], prev_state[2]);
	and _ECO_15743(w_eco15743, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15744(w_eco15744, !prev_cnt[14], prev_cnt[3], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15745(w_eco15745, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15746(w_eco15746, prev_cnt[4], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15747(w_eco15747, prev_cnt[5], !prev_cnt[6], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15748(w_eco15748, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15749(w_eco15749, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15750(w_eco15750, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15751(w_eco15751, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15752(w_eco15752, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15753(w_eco15753, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15754(w_eco15754, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15755(w_eco15755, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15756(w_eco15756, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15757(w_eco15757, !prev_cnt[14], prev_cnt[0], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15758(w_eco15758, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15759(w_eco15759, prev_cnt[5], !prev_cnt[6], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15760(w_eco15760, !prev_cnt[6], prev_cnt[7], prev_cnt[9], !rst, prev_state[1]);
	and _ECO_15761(w_eco15761, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15762(w_eco15762, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15763(w_eco15763, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15764(w_eco15764, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15765(w_eco15765, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15766(w_eco15766, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15767(w_eco15767, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15768(w_eco15768, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15769(w_eco15769, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15770(w_eco15770, !prev_cnt[14], prev_cnt[4], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15771(w_eco15771, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15772(w_eco15772, !prev_cnt[6], prev_cnt[7], prev_cnt[10], !rst, prev_state[1]);
	and _ECO_15773(w_eco15773, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15774(w_eco15774, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15775(w_eco15775, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15776(w_eco15776, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15777(w_eco15777, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15778(w_eco15778, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15779(w_eco15779, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15780(w_eco15780, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15781(w_eco15781, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15782(w_eco15782, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15783(w_eco15783, !prev_cnt[14], prev_cnt[5], !prev_cnt[6], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15784(w_eco15784, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], prev_cnt[12], !rst, prev_state[1]);
	and _ECO_15785(w_eco15785, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15786(w_eco15786, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15787(w_eco15787, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15788(w_eco15788, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15789(w_eco15789, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15790(w_eco15790, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15791(w_eco15791, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15792(w_eco15792, prev_cnt[1], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15793(w_eco15793, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15794(w_eco15794, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15795(w_eco15795, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15796(w_eco15796, !prev_cnt[14], !prev_cnt[6], prev_cnt[7], prev_cnt[13], !rst, prev_state[1]);
	and _ECO_15797(w_eco15797, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15798(w_eco15798, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15799(w_eco15799, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15800(w_eco15800, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15801(w_eco15801, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15802(w_eco15802, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15803(w_eco15803, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15804(w_eco15804, prev_cnt[2], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15805(w_eco15805, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15806(w_eco15806, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15807(w_eco15807, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15808(w_eco15808, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15809(w_eco15809, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15810(w_eco15810, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15811(w_eco15811, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15812(w_eco15812, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15813(w_eco15813, prev_cnt[3], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15814(w_eco15814, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15815(w_eco15815, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15816(w_eco15816, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15817(w_eco15817, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15818(w_eco15818, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15819(w_eco15819, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15820(w_eco15820, prev_cnt[0], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15821(w_eco15821, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15822(w_eco15822, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15823(w_eco15823, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15824(w_eco15824, prev_cnt[4], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15825(w_eco15825, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15826(w_eco15826, prev_cnt[5], !prev_cnt[6], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15827(w_eco15827, !prev_cnt[6], prev_cnt[7], !rst, prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	or _ECO_15828(w_eco15828, w_eco15484, w_eco15485, w_eco15486, w_eco15487, w_eco15488, w_eco15489, w_eco15490, w_eco15491, w_eco15492, w_eco15493, w_eco15494, w_eco15495, w_eco15496, w_eco15497, w_eco15498, w_eco15499, w_eco15500, w_eco15501, w_eco15502, w_eco15503, w_eco15504, w_eco15505, w_eco15506, w_eco15507, w_eco15508, w_eco15509, w_eco15510, w_eco15511, w_eco15512, w_eco15513, w_eco15514, w_eco15515, w_eco15516, w_eco15517, w_eco15518, w_eco15519, w_eco15520, w_eco15521, w_eco15522, w_eco15523, w_eco15524, w_eco15525, w_eco15526, w_eco15527, w_eco15528, w_eco15529, w_eco15530, w_eco15531, w_eco15532, w_eco15533, w_eco15534, w_eco15535, w_eco15536, w_eco15537, w_eco15538, w_eco15539, w_eco15540, w_eco15541, w_eco15542, w_eco15543, w_eco15544, w_eco15545, w_eco15546, w_eco15547, w_eco15548, w_eco15549, w_eco15550, w_eco15551, w_eco15552, w_eco15553, w_eco15554, w_eco15555, w_eco15556, w_eco15557, w_eco15558, w_eco15559, w_eco15560, w_eco15561, w_eco15562, w_eco15563, w_eco15564, w_eco15565, w_eco15566, w_eco15567, w_eco15568, w_eco15569, w_eco15570, w_eco15571, w_eco15572, w_eco15573, w_eco15574, w_eco15575, w_eco15576, w_eco15577, w_eco15578, w_eco15579, w_eco15580, w_eco15581, w_eco15582, w_eco15583, w_eco15584, w_eco15585, w_eco15586, w_eco15587, w_eco15588, w_eco15589, w_eco15590, w_eco15591, w_eco15592, w_eco15593, w_eco15594, w_eco15595, w_eco15596, w_eco15597, w_eco15598, w_eco15599, w_eco15600, w_eco15601, w_eco15602, w_eco15603, w_eco15604, w_eco15605, w_eco15606, w_eco15607, w_eco15608, w_eco15609, w_eco15610, w_eco15611, w_eco15612, w_eco15613, w_eco15614, w_eco15615, w_eco15616, w_eco15617, w_eco15618, w_eco15619, w_eco15620, w_eco15621, w_eco15622, w_eco15623, w_eco15624, w_eco15625, w_eco15626, w_eco15627, w_eco15628, w_eco15629, w_eco15630, w_eco15631, w_eco15632, w_eco15633, w_eco15634, w_eco15635, w_eco15636, w_eco15637, w_eco15638, w_eco15639, w_eco15640, w_eco15641, w_eco15642, w_eco15643, w_eco15644, w_eco15645, w_eco15646, w_eco15647, w_eco15648, w_eco15649, w_eco15650, w_eco15651, w_eco15652, w_eco15653, w_eco15654, w_eco15655, w_eco15656, w_eco15657, w_eco15658, w_eco15659, w_eco15660, w_eco15661, w_eco15662, w_eco15663, w_eco15664, w_eco15665, w_eco15666, w_eco15667, w_eco15668, w_eco15669, w_eco15670, w_eco15671, w_eco15672, w_eco15673, w_eco15674, w_eco15675, w_eco15676, w_eco15677, w_eco15678, w_eco15679, w_eco15680, w_eco15681, w_eco15682, w_eco15683, w_eco15684, w_eco15685, w_eco15686, w_eco15687, w_eco15688, w_eco15689, w_eco15690, w_eco15691, w_eco15692, w_eco15693, w_eco15694, w_eco15695, w_eco15696, w_eco15697, w_eco15698, w_eco15699, w_eco15700, w_eco15701, w_eco15702, w_eco15703, w_eco15704, w_eco15705, w_eco15706, w_eco15707, w_eco15708, w_eco15709, w_eco15710, w_eco15711, w_eco15712, w_eco15713, w_eco15714, w_eco15715, w_eco15716, w_eco15717, w_eco15718, w_eco15719, w_eco15720, w_eco15721, w_eco15722, w_eco15723, w_eco15724, w_eco15725, w_eco15726, w_eco15727, w_eco15728, w_eco15729, w_eco15730, w_eco15731, w_eco15732, w_eco15733, w_eco15734, w_eco15735, w_eco15736, w_eco15737, w_eco15738, w_eco15739, w_eco15740, w_eco15741, w_eco15742, w_eco15743, w_eco15744, w_eco15745, w_eco15746, w_eco15747, w_eco15748, w_eco15749, w_eco15750, w_eco15751, w_eco15752, w_eco15753, w_eco15754, w_eco15755, w_eco15756, w_eco15757, w_eco15758, w_eco15759, w_eco15760, w_eco15761, w_eco15762, w_eco15763, w_eco15764, w_eco15765, w_eco15766, w_eco15767, w_eco15768, w_eco15769, w_eco15770, w_eco15771, w_eco15772, w_eco15773, w_eco15774, w_eco15775, w_eco15776, w_eco15777, w_eco15778, w_eco15779, w_eco15780, w_eco15781, w_eco15782, w_eco15783, w_eco15784, w_eco15785, w_eco15786, w_eco15787, w_eco15788, w_eco15789, w_eco15790, w_eco15791, w_eco15792, w_eco15793, w_eco15794, w_eco15795, w_eco15796, w_eco15797, w_eco15798, w_eco15799, w_eco15800, w_eco15801, w_eco15802, w_eco15803, w_eco15804, w_eco15805, w_eco15806, w_eco15807, w_eco15808, w_eco15809, w_eco15810, w_eco15811, w_eco15812, w_eco15813, w_eco15814, w_eco15815, w_eco15816, w_eco15817, w_eco15818, w_eco15819, w_eco15820, w_eco15821, w_eco15822, w_eco15823, w_eco15824, w_eco15825, w_eco15826, w_eco15827);
	xor _ECO_out17(cnt[8], sub_wire17, w_eco15828);
	and _ECO_15829(w_eco15829, prev_cnt[15], rst);
	and _ECO_15830(w_eco15830, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[0]);
	and _ECO_15831(w_eco15831, prev_cnt[15], prev_state[1], prev_cnt_len[0]);
	and _ECO_15832(w_eco15832, prev_cnt[15], !ena, prev_cnt_len[0]);
	and _ECO_15833(w_eco15833, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[0]);
	and _ECO_15834(w_eco15834, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15835(w_eco15835, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15836(w_eco15836, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15837(w_eco15837, prev_cnt[15], prev_state[1], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15838(w_eco15838, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15839(w_eco15839, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15840(w_eco15840, prev_cnt[15], prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15841(w_eco15841, !prev_cnt[15], !ena, !rst, prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15842(w_eco15842, prev_cnt[15], !ena, prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15843(w_eco15843, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15844(w_eco15844, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15845(w_eco15845, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15846(w_eco15846, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15847(w_eco15847, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15848(w_eco15848, prev_cnt[15], prev_state[1], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15849(w_eco15849, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15850(w_eco15850, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15851(w_eco15851, prev_cnt[15], prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15852(w_eco15852, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[9], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15853(w_eco15853, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[3], !prev_cnt_len[1]);
	and _ECO_15854(w_eco15854, prev_cnt[15], !ena, prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15855(w_eco15855, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15856(w_eco15856, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15857(w_eco15857, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15858(w_eco15858, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15859(w_eco15859, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15860(w_eco15860, prev_cnt[15], prev_state[1], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15861(w_eco15861, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15862(w_eco15862, prev_cnt[15], prev_state[1], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15863(w_eco15863, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15864(w_eco15864, prev_cnt[15], !ena, prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15865(w_eco15865, !prev_cnt[15], !ena, !rst, prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15866(w_eco15866, !prev_cnt[15], !ena, !rst, prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15867(w_eco15867, prev_cnt[15], !ena, prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15868(w_eco15868, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15869(w_eco15869, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15870(w_eco15870, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15871(w_eco15871, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15872(w_eco15872, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15873(w_eco15873, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15874(w_eco15874, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15875(w_eco15875, prev_cnt[15], prev_state[1], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15876(w_eco15876, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15877(w_eco15877, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15878(w_eco15878, prev_cnt[15], prev_state[1], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15879(w_eco15879, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[2], !prev_cnt_len[1]);
	and _ECO_15880(w_eco15880, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15881(w_eco15881, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15882(w_eco15882, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15883(w_eco15883, prev_cnt[15], !ena, prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15884(w_eco15884, !prev_cnt[15], !ena, !rst, prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15885(w_eco15885, prev_cnt[15], !ena, prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15886(w_eco15886, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15887(w_eco15887, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15888(w_eco15888, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15889(w_eco15889, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15890(w_eco15890, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15891(w_eco15891, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15892(w_eco15892, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15893(w_eco15893, prev_cnt[15], prev_state[1], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15894(w_eco15894, prev_cnt[15], prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15895(w_eco15895, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15896(w_eco15896, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15897(w_eco15897, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[13], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15898(w_eco15898, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15899(w_eco15899, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[5], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15900(w_eco15900, prev_cnt[15], !ena, prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15901(w_eco15901, !prev_cnt[15], !ena, !rst, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15902(w_eco15902, !prev_cnt[15], !ena, !rst, prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15903(w_eco15903, prev_cnt[15], !ena, prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15904(w_eco15904, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15905(w_eco15905, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15906(w_eco15906, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15907(w_eco15907, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15908(w_eco15908, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15909(w_eco15909, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15910(w_eco15910, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15911(w_eco15911, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15912(w_eco15912, prev_cnt[15], prev_state[1], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15913(w_eco15913, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15914(w_eco15914, prev_cnt[15], prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15915(w_eco15915, !prev_cnt[15], !rst, prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15916(w_eco15916, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[7], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15917(w_eco15917, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15918(w_eco15918, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[11], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15919(w_eco15919, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[4], !prev_cnt_len[6], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15920(w_eco15920, prev_cnt[15], !ena, prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15921(w_eco15921, prev_cnt[15], !ena, prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15922(w_eco15922, !prev_cnt[15], !ena, !rst, prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15923(w_eco15923, !prev_cnt[15], !ena, !rst, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15924(w_eco15924, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15925(w_eco15925, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15926(w_eco15926, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15927(w_eco15927, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15928(w_eco15928, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15929(w_eco15929, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15930(w_eco15930, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15931(w_eco15931, prev_cnt[15], prev_state[1], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15932(w_eco15932, !prev_cnt[15], !rst, prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15933(w_eco15933, !prev_cnt[15], !rst, prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15934(w_eco15934, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15935(w_eco15935, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15936(w_eco15936, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[10], !prev_cnt_len[8], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15937(w_eco15937, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15938(w_eco15938, prev_cnt[15], !ena, prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15939(w_eco15939, !prev_cnt[15], !ena, !rst, prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15940(w_eco15940, prev_cnt[15], !ena, prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15941(w_eco15941, !prev_cnt[15], !ena, !rst, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15942(w_eco15942, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15943(w_eco15943, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15944(w_eco15944, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15945(w_eco15945, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15946(w_eco15946, prev_cnt[15], !prev_state[4], !prev_state[2], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15947(w_eco15947, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15948(w_eco15948, prev_cnt[15], prev_state[1], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15949(w_eco15949, !prev_cnt[15], !rst, prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15950(w_eco15950, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15951(w_eco15951, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15952(w_eco15952, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], prev_cnt_len[8], !prev_cnt_len[9]);
	and _ECO_15953(w_eco15953, !prev_cnt[15], !rst, prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15954(w_eco15954, prev_cnt[15], !ena, prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15955(w_eco15955, !prev_cnt[15], !ena, !rst, prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15956(w_eco15956, !prev_cnt[15], !ena, !rst, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15957(w_eco15957, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15958(w_eco15958, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15959(w_eco15959, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15960(w_eco15960, !prev_cnt[15], !rst, !prev_state[4], !prev_state[2], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15961(w_eco15961, !prev_cnt[15], !rst, prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15962(w_eco15962, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[15], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15963(w_eco15963, !prev_cnt[15], !rst, prev_state[0], prev_cnt_len[12], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15964(w_eco15964, !prev_cnt[15], !rst, prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[0]);
	and _ECO_15965(w_eco15965, prev_cnt[15], !ena, prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15966(w_eco15966, !prev_cnt[15], !ena, !rst, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15967(w_eco15967, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15968(w_eco15968, ena, !rst, prev_state[4], prev_state[3], !prev_state[2], !prev_state[1], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15969(w_eco15969, prev_cnt[15], !prev_state[3], prev_state[0], prev_cnt_len[14], !prev_cnt_len[12], !prev_cnt_len[10], !prev_cnt_len[11], !prev_cnt_len[9]);
	and _ECO_15970(w_eco15970, !prev_cnt[15], !rst, prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], prev_cnt_len[6], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15971(w_eco15971, !prev_cnt[15], !ena, !rst, !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15972(w_eco15972, ena, !rst, prev_state[3], prev_state[2], !prev_state[1], prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	and _ECO_15973(w_eco15973, !prev_cnt[15], !rst, prev_state[0], !prev_cnt_len[14], !prev_cnt_len[15], !prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[5], !prev_cnt_len[7], !prev_cnt_len[3], !prev_cnt_len[2], !prev_cnt_len[0]);
	or _ECO_15974(w_eco15974, w_eco15829, w_eco15830, w_eco15831, w_eco15832, w_eco15833, w_eco15834, w_eco15835, w_eco15836, w_eco15837, w_eco15838, w_eco15839, w_eco15840, w_eco15841, w_eco15842, w_eco15843, w_eco15844, w_eco15845, w_eco15846, w_eco15847, w_eco15848, w_eco15849, w_eco15850, w_eco15851, w_eco15852, w_eco15853, w_eco15854, w_eco15855, w_eco15856, w_eco15857, w_eco15858, w_eco15859, w_eco15860, w_eco15861, w_eco15862, w_eco15863, w_eco15864, w_eco15865, w_eco15866, w_eco15867, w_eco15868, w_eco15869, w_eco15870, w_eco15871, w_eco15872, w_eco15873, w_eco15874, w_eco15875, w_eco15876, w_eco15877, w_eco15878, w_eco15879, w_eco15880, w_eco15881, w_eco15882, w_eco15883, w_eco15884, w_eco15885, w_eco15886, w_eco15887, w_eco15888, w_eco15889, w_eco15890, w_eco15891, w_eco15892, w_eco15893, w_eco15894, w_eco15895, w_eco15896, w_eco15897, w_eco15898, w_eco15899, w_eco15900, w_eco15901, w_eco15902, w_eco15903, w_eco15904, w_eco15905, w_eco15906, w_eco15907, w_eco15908, w_eco15909, w_eco15910, w_eco15911, w_eco15912, w_eco15913, w_eco15914, w_eco15915, w_eco15916, w_eco15917, w_eco15918, w_eco15919, w_eco15920, w_eco15921, w_eco15922, w_eco15923, w_eco15924, w_eco15925, w_eco15926, w_eco15927, w_eco15928, w_eco15929, w_eco15930, w_eco15931, w_eco15932, w_eco15933, w_eco15934, w_eco15935, w_eco15936, w_eco15937, w_eco15938, w_eco15939, w_eco15940, w_eco15941, w_eco15942, w_eco15943, w_eco15944, w_eco15945, w_eco15946, w_eco15947, w_eco15948, w_eco15949, w_eco15950, w_eco15951, w_eco15952, w_eco15953, w_eco15954, w_eco15955, w_eco15956, w_eco15957, w_eco15958, w_eco15959, w_eco15960, w_eco15961, w_eco15962, w_eco15963, w_eco15964, w_eco15965, w_eco15966, w_eco15967, w_eco15968, w_eco15969, w_eco15970, w_eco15971, w_eco15972, w_eco15973);
	xor _ECO_out18(Done, sub_wire18, w_eco15974);

endmodule