module top(parity,overflow,greater,is_eq,less,y,a,b,op);
	input [7:0]a, b;
	input [1:0]op;
	output parity, overflow, greater, is_eq, less;
	output [7:0]y;
	wire \mux_44_12_g156/w_0, \mux_44_12_g156/w_1, \mux_44_12_g156/w_2, \mux_temp_y_21_12_g792/w_0, \mux_temp_y_21_12_g792/w_1, \mux_temp_y_21_12_g19/w_0, \mux_temp_y_21_12_g19/w_1, \mux_temp_y_21_12_g19/w_2, \mux_temp_y_21_12_g19/w_3, \mux_temp_y_21_12_g18/w_0, \mux_temp_y_21_12_g18/w_1, \mux_temp_y_21_12_g18/w_2, \mux_temp_y_21_12_g18/w_3, \mux_temp_y_21_12_g17/w_0, \mux_temp_y_21_12_g17/w_1, \mux_temp_y_21_12_g17/w_2, \mux_temp_y_21_12_g17/w_3, \mux_temp_y_21_12_g16/w_0, \mux_temp_y_21_12_g16/w_1, \mux_temp_y_21_12_g16/w_2, \mux_temp_y_21_12_g16/w_3, \mux_temp_y_21_12_g15/w_0, \mux_temp_y_21_12_g15/w_1, \mux_temp_y_21_12_g15/w_2, \mux_temp_y_21_12_g15/w_3, \mux_temp_y_21_12_g10/w_0, \mux_temp_y_21_12_g10/w_1, \mux_temp_y_21_12_g10/w_2, \mux_temp_y_21_12_g10/w_3, sub_29_29_n_1105, sub_29_29_n_1103, sub_29_29_n_320, sub_29_29_n_69, sub_29_29_n_66, sub_29_29_n_63, sub_29_29_n_59, sub_29_29_n_54, sub_29_29_n_37, sub_29_29_n_32, n_1123, n_1114, n_1113, n_1112, n_1111, n_1106, n_1104, n_1102, n_1101, n_1099, n_1098, n_1097, n_1096, n_1095, n_988, n_987, n_986, n_985, n_984, n_983, n_982, n_981, n_980, n_979, n_978, n_977, n_976, n_975, n_974, n_973, n_972, n_971, n_970, n_969, n_968, n_967, n_966, n_965, n_964, n_963, n_962, n_961, n_960, n_959, n_958, n_957, n_956, n_955, n_954, n_953, n_952, n_951, n_950, n_949, n_948, n_947, n_946, n_945, n_944, n_943, n_942, n_940, n_939, n_938, n_937, n_936, n_935, n_934, n_933, n_932, n_931, n_930, n_929, n_928, n_927, n_926, n_925, n_924, n_923, n_922, n_921, n_920, n_919, n_918, n_917, n_916, n_915, n_914, n_913, n_912, n_911, n_910, n_909, n_908, n_907, n_906, n_905, n_904, n_903, n_902, n_901, n_900, n_898, n_897, n_895, n_894, n_892, n_891, n_890, n_889, n_888, n_887, n_886, n_885, n_884, n_883, n_882, n_881, n_880, n_878, n_877, n_876, n_875, n_874, n_873, n_872, n_871, n_870, n_869, n_867, n_866, n_865, n_864, n_863, n_862, n_861, n_860, n_859, n_858, n_857, n_856, n_840, n_827, n_806, n_805, n_620, n_619, n_618, n_617, n_616, n_615, n_437, n_436, n_435, n_431, n_429, n_428, n_419, n_416, n_415, n_397, n_395, n_379, n_367, n_323, n_318, n_308, n_301, n_300, n_298, n_136, n_135, n_133, n_132, n_131, n_130, n_129, n_77, n_76, n_75, n_74, n_73, n_43, n_41, n_39, n_38, n_37, n_35, n_34, n_33, n_31, n_30, n_29, n_26, n_25, n_23, n_22, n_21, n_19, n_18, n_17, n_16, gt_39_12_n_57, gt_39_12_n_52, gt_39_12_n_46, gt_25_24_n_35, add_24_29_n_1115, add_24_29_n_57, add_24_29_n_55, add_24_29_n_53, add_24_29_n_51, add_24_29_n_50, add_24_29_n_49, add_24_29_n_48, add_24_29_n_47, add_24_29_n_43, add_24_29_n_39, add_24_29_n_37, add_24_29_n_33, add_24_29_n_27, less, is_eq, greater, overflow, parity, oe, clk, \mux_44_12_g156/data0;
	wire [7:0]y;
	wire [1:0]op;
	wire [7:0]b, a;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, sub_wire1, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, sub_wire2, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, sub_wire3, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, sub_wire4, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634, w_eco1635, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833, w_eco1834, sub_wire5, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914, w_eco1915, w_eco1916, w_eco1917, w_eco1918, w_eco1919, w_eco1920, w_eco1921, w_eco1922, w_eco1923, w_eco1924, w_eco1925, w_eco1926, w_eco1927, w_eco1928, w_eco1929, w_eco1930, w_eco1931, w_eco1932, w_eco1933, w_eco1934, w_eco1935, w_eco1936, w_eco1937, w_eco1938, w_eco1939, w_eco1940, w_eco1941, w_eco1942, w_eco1943, w_eco1944, w_eco1945, w_eco1946, w_eco1947, w_eco1948, w_eco1949, w_eco1950, w_eco1951, w_eco1952, w_eco1953, w_eco1954, w_eco1955, w_eco1956, w_eco1957, w_eco1958, w_eco1959, w_eco1960, w_eco1961, w_eco1962, w_eco1963, w_eco1964, w_eco1965, w_eco1966, w_eco1967, w_eco1968, w_eco1969, w_eco1970, w_eco1971, w_eco1972, w_eco1973, w_eco1974, w_eco1975, w_eco1976, w_eco1977, w_eco1978, w_eco1979, w_eco1980, w_eco1981, w_eco1982, w_eco1983, w_eco1984, w_eco1985, w_eco1986, w_eco1987, w_eco1988, w_eco1989, w_eco1990, w_eco1991, w_eco1992, w_eco1993, w_eco1994, w_eco1995, w_eco1996, w_eco1997, w_eco1998, w_eco1999, w_eco2000, w_eco2001, w_eco2002, w_eco2003, w_eco2004, w_eco2005, w_eco2006, w_eco2007, w_eco2008, w_eco2009, w_eco2010, w_eco2011, w_eco2012, w_eco2013, w_eco2014, w_eco2015, w_eco2016, w_eco2017, w_eco2018, w_eco2019, w_eco2020, w_eco2021, w_eco2022, w_eco2023, w_eco2024, w_eco2025, w_eco2026, w_eco2027, w_eco2028, w_eco2029, w_eco2030, w_eco2031, w_eco2032, w_eco2033, w_eco2034, w_eco2035, w_eco2036, w_eco2037, w_eco2038, w_eco2039, w_eco2040, w_eco2041, w_eco2042, w_eco2043, w_eco2044, w_eco2045, w_eco2046, w_eco2047, w_eco2048, w_eco2049, w_eco2050, w_eco2051, w_eco2052, w_eco2053, w_eco2054, w_eco2055, w_eco2056, w_eco2057, w_eco2058, w_eco2059, w_eco2060, w_eco2061, w_eco2062, w_eco2063, w_eco2064, w_eco2065, w_eco2066, w_eco2067, w_eco2068, w_eco2069, w_eco2070, w_eco2071, w_eco2072, w_eco2073, w_eco2074, w_eco2075, w_eco2076, w_eco2077, w_eco2078, w_eco2079, w_eco2080, w_eco2081, w_eco2082, w_eco2083, w_eco2084, w_eco2085, w_eco2086, w_eco2087, w_eco2088, w_eco2089, w_eco2090, w_eco2091, w_eco2092, w_eco2093, w_eco2094, w_eco2095, w_eco2096, w_eco2097, w_eco2098, w_eco2099, w_eco2100, w_eco2101, w_eco2102, w_eco2103, w_eco2104, w_eco2105, w_eco2106, w_eco2107, w_eco2108, w_eco2109, w_eco2110, w_eco2111, w_eco2112, w_eco2113, w_eco2114, w_eco2115, w_eco2116, w_eco2117, w_eco2118, w_eco2119, w_eco2120, w_eco2121, w_eco2122, w_eco2123, w_eco2124, w_eco2125, w_eco2126, w_eco2127, w_eco2128, w_eco2129, w_eco2130, w_eco2131, w_eco2132, w_eco2133, w_eco2134, w_eco2135, w_eco2136, w_eco2137, w_eco2138, w_eco2139, w_eco2140, w_eco2141, w_eco2142, w_eco2143, w_eco2144, w_eco2145, w_eco2146, w_eco2147, w_eco2148, w_eco2149, w_eco2150, w_eco2151, w_eco2152, w_eco2153, w_eco2154, w_eco2155, w_eco2156, w_eco2157, w_eco2158, w_eco2159, w_eco2160, w_eco2161, w_eco2162, w_eco2163, w_eco2164, w_eco2165, w_eco2166, w_eco2167, w_eco2168, w_eco2169, w_eco2170, w_eco2171, w_eco2172, w_eco2173, w_eco2174, w_eco2175, w_eco2176, w_eco2177, w_eco2178, w_eco2179, w_eco2180, w_eco2181, w_eco2182, w_eco2183, w_eco2184, w_eco2185, w_eco2186, w_eco2187, w_eco2188, w_eco2189, w_eco2190, w_eco2191, w_eco2192, w_eco2193, w_eco2194, w_eco2195, w_eco2196, w_eco2197, w_eco2198, w_eco2199, w_eco2200, w_eco2201, w_eco2202, w_eco2203, w_eco2204, w_eco2205, w_eco2206, w_eco2207, w_eco2208, w_eco2209, w_eco2210, w_eco2211, w_eco2212, w_eco2213, w_eco2214, w_eco2215, w_eco2216, w_eco2217, w_eco2218, w_eco2219, w_eco2220, w_eco2221, w_eco2222, w_eco2223, w_eco2224, w_eco2225, w_eco2226, w_eco2227, w_eco2228, w_eco2229, w_eco2230, w_eco2231, w_eco2232, w_eco2233, w_eco2234, w_eco2235, w_eco2236, w_eco2237, w_eco2238, w_eco2239, w_eco2240, w_eco2241, w_eco2242, w_eco2243, w_eco2244, w_eco2245, w_eco2246, w_eco2247, w_eco2248, w_eco2249, w_eco2250, w_eco2251, w_eco2252, w_eco2253, w_eco2254, w_eco2255, w_eco2256, w_eco2257, w_eco2258, w_eco2259, w_eco2260, w_eco2261, w_eco2262, w_eco2263, w_eco2264, w_eco2265, w_eco2266, w_eco2267, w_eco2268, w_eco2269, w_eco2270, w_eco2271, w_eco2272, w_eco2273, w_eco2274, w_eco2275, w_eco2276, w_eco2277, w_eco2278, w_eco2279, w_eco2280, w_eco2281, w_eco2282, w_eco2283, w_eco2284, w_eco2285, w_eco2286, w_eco2287, w_eco2288, w_eco2289, w_eco2290, w_eco2291, w_eco2292, w_eco2293, w_eco2294, w_eco2295, w_eco2296, w_eco2297, w_eco2298, w_eco2299, w_eco2300, w_eco2301, w_eco2302, w_eco2303, w_eco2304, w_eco2305, w_eco2306, w_eco2307, w_eco2308, w_eco2309, w_eco2310, w_eco2311, w_eco2312, w_eco2313, w_eco2314, w_eco2315, w_eco2316, w_eco2317, w_eco2318, w_eco2319, w_eco2320, w_eco2321, w_eco2322, w_eco2323, w_eco2324, w_eco2325, w_eco2326, w_eco2327, w_eco2328, w_eco2329, w_eco2330, w_eco2331, w_eco2332, w_eco2333, w_eco2334, w_eco2335, w_eco2336, w_eco2337, w_eco2338, w_eco2339, w_eco2340, w_eco2341, w_eco2342, w_eco2343, w_eco2344, w_eco2345, w_eco2346, w_eco2347, w_eco2348, w_eco2349, w_eco2350, w_eco2351, w_eco2352, w_eco2353, w_eco2354, w_eco2355, w_eco2356, w_eco2357, w_eco2358, w_eco2359, w_eco2360, w_eco2361, w_eco2362, w_eco2363, w_eco2364, w_eco2365, w_eco2366, w_eco2367, w_eco2368, w_eco2369, w_eco2370, w_eco2371, w_eco2372, w_eco2373, w_eco2374, w_eco2375, w_eco2376, w_eco2377, w_eco2378, w_eco2379, w_eco2380, w_eco2381, w_eco2382, w_eco2383, w_eco2384, w_eco2385, w_eco2386, w_eco2387, w_eco2388, w_eco2389, w_eco2390, w_eco2391, w_eco2392, w_eco2393, w_eco2394, w_eco2395, w_eco2396, w_eco2397, w_eco2398, w_eco2399, w_eco2400, w_eco2401, w_eco2402, w_eco2403, w_eco2404, w_eco2405, w_eco2406, w_eco2407, w_eco2408, w_eco2409, w_eco2410, w_eco2411, w_eco2412, w_eco2413, w_eco2414, w_eco2415, w_eco2416, w_eco2417, w_eco2418, w_eco2419, w_eco2420, w_eco2421, w_eco2422, w_eco2423, w_eco2424, w_eco2425, w_eco2426, w_eco2427, w_eco2428, w_eco2429, w_eco2430, w_eco2431, w_eco2432, w_eco2433, w_eco2434, w_eco2435, w_eco2436, w_eco2437, w_eco2438, w_eco2439, w_eco2440, w_eco2441, w_eco2442, w_eco2443, w_eco2444, w_eco2445, w_eco2446, w_eco2447, w_eco2448, w_eco2449, w_eco2450, w_eco2451, w_eco2452, w_eco2453, w_eco2454, w_eco2455, w_eco2456, w_eco2457, w_eco2458, w_eco2459, w_eco2460, w_eco2461, w_eco2462, w_eco2463, w_eco2464, w_eco2465, w_eco2466, w_eco2467, w_eco2468, w_eco2469, w_eco2470, w_eco2471, w_eco2472, w_eco2473, w_eco2474, w_eco2475, w_eco2476, w_eco2477, w_eco2478, w_eco2479, w_eco2480, w_eco2481, w_eco2482, w_eco2483, w_eco2484, w_eco2485, w_eco2486, w_eco2487, sub_wire6, w_eco2488, w_eco2489, w_eco2490, w_eco2491, w_eco2492, w_eco2493, w_eco2494, w_eco2495, w_eco2496, w_eco2497, w_eco2498, w_eco2499, w_eco2500, w_eco2501, w_eco2502, w_eco2503, w_eco2504, w_eco2505, w_eco2506, w_eco2507, w_eco2508, w_eco2509, w_eco2510, w_eco2511, w_eco2512, w_eco2513, w_eco2514, w_eco2515, w_eco2516, w_eco2517, w_eco2518, w_eco2519, w_eco2520, w_eco2521, w_eco2522, w_eco2523, w_eco2524, w_eco2525, w_eco2526, w_eco2527, w_eco2528, w_eco2529, w_eco2530, w_eco2531, w_eco2532, w_eco2533, w_eco2534, w_eco2535, w_eco2536, w_eco2537, w_eco2538, w_eco2539, w_eco2540, w_eco2541, w_eco2542, w_eco2543, w_eco2544, w_eco2545, w_eco2546, w_eco2547, w_eco2548, w_eco2549, w_eco2550, w_eco2551, w_eco2552, w_eco2553, w_eco2554, w_eco2555, w_eco2556, w_eco2557, w_eco2558, w_eco2559, w_eco2560, w_eco2561, w_eco2562, w_eco2563, w_eco2564, w_eco2565, w_eco2566, w_eco2567, w_eco2568, w_eco2569, w_eco2570, w_eco2571, w_eco2572, w_eco2573, w_eco2574, w_eco2575, w_eco2576, w_eco2577, w_eco2578, w_eco2579, w_eco2580, w_eco2581, w_eco2582, w_eco2583, w_eco2584, w_eco2585, w_eco2586, w_eco2587, w_eco2588, w_eco2589, w_eco2590, w_eco2591, w_eco2592, w_eco2593, w_eco2594, w_eco2595, w_eco2596, w_eco2597, w_eco2598, w_eco2599, w_eco2600, w_eco2601, w_eco2602, w_eco2603, w_eco2604, w_eco2605, w_eco2606, w_eco2607, w_eco2608, w_eco2609, w_eco2610, w_eco2611, w_eco2612, w_eco2613, w_eco2614, w_eco2615, w_eco2616, w_eco2617, w_eco2618, w_eco2619, w_eco2620, w_eco2621, w_eco2622, w_eco2623, w_eco2624, w_eco2625, w_eco2626, w_eco2627, w_eco2628, w_eco2629, w_eco2630, w_eco2631, w_eco2632, w_eco2633, w_eco2634, w_eco2635, w_eco2636, w_eco2637, w_eco2638, w_eco2639, w_eco2640, w_eco2641, w_eco2642, w_eco2643, w_eco2644, w_eco2645, w_eco2646, w_eco2647, w_eco2648, w_eco2649, w_eco2650, w_eco2651, w_eco2652, w_eco2653, w_eco2654, w_eco2655, w_eco2656, w_eco2657, w_eco2658, w_eco2659, w_eco2660, w_eco2661, w_eco2662, w_eco2663, w_eco2664, w_eco2665, w_eco2666, w_eco2667, w_eco2668, w_eco2669, w_eco2670, w_eco2671, w_eco2672, w_eco2673, w_eco2674, w_eco2675, w_eco2676, w_eco2677, w_eco2678, w_eco2679, w_eco2680, w_eco2681, w_eco2682, w_eco2683, w_eco2684, w_eco2685, w_eco2686, w_eco2687, w_eco2688, w_eco2689, w_eco2690, w_eco2691, w_eco2692, w_eco2693, w_eco2694, w_eco2695, w_eco2696, w_eco2697, w_eco2698, w_eco2699, w_eco2700, w_eco2701, w_eco2702, w_eco2703, w_eco2704, w_eco2705, w_eco2706, w_eco2707, w_eco2708, w_eco2709, w_eco2710, w_eco2711, w_eco2712, w_eco2713, w_eco2714, w_eco2715, w_eco2716, w_eco2717, w_eco2718, w_eco2719, w_eco2720, w_eco2721, w_eco2722, w_eco2723, w_eco2724, w_eco2725, w_eco2726, w_eco2727, w_eco2728, w_eco2729, w_eco2730, w_eco2731, w_eco2732, w_eco2733, w_eco2734, w_eco2735, w_eco2736, w_eco2737, w_eco2738, w_eco2739, w_eco2740, w_eco2741, w_eco2742, w_eco2743, w_eco2744, w_eco2745, w_eco2746, w_eco2747, w_eco2748, w_eco2749, w_eco2750, w_eco2751, w_eco2752, w_eco2753, w_eco2754, w_eco2755, w_eco2756, w_eco2757, w_eco2758, w_eco2759, w_eco2760, w_eco2761, w_eco2762, w_eco2763, w_eco2764, w_eco2765, w_eco2766, w_eco2767, w_eco2768, w_eco2769, w_eco2770, w_eco2771, w_eco2772, w_eco2773, w_eco2774, w_eco2775, w_eco2776, w_eco2777, w_eco2778, w_eco2779, w_eco2780, w_eco2781, w_eco2782, w_eco2783, w_eco2784, w_eco2785, w_eco2786, w_eco2787, w_eco2788, w_eco2789, w_eco2790, w_eco2791, w_eco2792, w_eco2793, w_eco2794, w_eco2795, w_eco2796, w_eco2797, w_eco2798, w_eco2799, w_eco2800, w_eco2801, w_eco2802, w_eco2803, w_eco2804, w_eco2805, w_eco2806, w_eco2807, w_eco2808, w_eco2809, w_eco2810, w_eco2811, w_eco2812, w_eco2813, w_eco2814, w_eco2815, w_eco2816, w_eco2817, w_eco2818, w_eco2819, w_eco2820, w_eco2821, w_eco2822, w_eco2823, w_eco2824, w_eco2825, w_eco2826, w_eco2827, w_eco2828, w_eco2829, w_eco2830, w_eco2831, w_eco2832, w_eco2833, w_eco2834, w_eco2835, w_eco2836, w_eco2837, w_eco2838, w_eco2839, w_eco2840, w_eco2841, w_eco2842, w_eco2843, w_eco2844, w_eco2845, w_eco2846, w_eco2847, w_eco2848, w_eco2849, w_eco2850, w_eco2851, w_eco2852, w_eco2853, w_eco2854, w_eco2855, w_eco2856, w_eco2857, w_eco2858, w_eco2859, w_eco2860, w_eco2861, w_eco2862, w_eco2863, w_eco2864, w_eco2865, w_eco2866, w_eco2867, w_eco2868, w_eco2869, w_eco2870, w_eco2871, w_eco2872, w_eco2873, w_eco2874, w_eco2875, w_eco2876, w_eco2877, w_eco2878, w_eco2879, w_eco2880, w_eco2881, w_eco2882, w_eco2883, w_eco2884, w_eco2885, w_eco2886, w_eco2887, w_eco2888, w_eco2889, w_eco2890, w_eco2891, w_eco2892, w_eco2893, w_eco2894, w_eco2895, w_eco2896, w_eco2897, w_eco2898, w_eco2899, w_eco2900, w_eco2901, w_eco2902, w_eco2903, w_eco2904, w_eco2905, w_eco2906, w_eco2907, w_eco2908, w_eco2909, w_eco2910, w_eco2911, w_eco2912, w_eco2913, w_eco2914, w_eco2915, w_eco2916, w_eco2917, w_eco2918, w_eco2919, w_eco2920, w_eco2921, w_eco2922, w_eco2923, w_eco2924, w_eco2925, w_eco2926, w_eco2927, w_eco2928, w_eco2929, w_eco2930, w_eco2931, w_eco2932, w_eco2933, w_eco2934, w_eco2935, w_eco2936, w_eco2937, w_eco2938, w_eco2939, w_eco2940, w_eco2941, w_eco2942, w_eco2943, w_eco2944, w_eco2945, w_eco2946, w_eco2947, w_eco2948, w_eco2949, w_eco2950, w_eco2951, w_eco2952, w_eco2953, w_eco2954, w_eco2955, w_eco2956, w_eco2957, w_eco2958, w_eco2959, w_eco2960, w_eco2961, w_eco2962, w_eco2963, w_eco2964, w_eco2965, w_eco2966, w_eco2967, w_eco2968, w_eco2969, w_eco2970, w_eco2971, w_eco2972, w_eco2973, w_eco2974, w_eco2975, w_eco2976, w_eco2977, w_eco2978, w_eco2979, w_eco2980, w_eco2981, w_eco2982, w_eco2983, w_eco2984, w_eco2985, w_eco2986, w_eco2987, w_eco2988, w_eco2989, w_eco2990, w_eco2991, w_eco2992, w_eco2993, w_eco2994, w_eco2995, w_eco2996, w_eco2997, w_eco2998, w_eco2999, w_eco3000, w_eco3001, w_eco3002, w_eco3003, w_eco3004, w_eco3005, w_eco3006, w_eco3007, w_eco3008, w_eco3009, w_eco3010, w_eco3011, w_eco3012, w_eco3013, w_eco3014, w_eco3015, w_eco3016, w_eco3017, w_eco3018, w_eco3019, w_eco3020, w_eco3021, w_eco3022, w_eco3023, w_eco3024, w_eco3025, w_eco3026, w_eco3027, w_eco3028, w_eco3029, w_eco3030, w_eco3031, w_eco3032, w_eco3033, w_eco3034, w_eco3035, w_eco3036, w_eco3037, w_eco3038, w_eco3039, w_eco3040, w_eco3041, w_eco3042, w_eco3043, w_eco3044, w_eco3045, w_eco3046, w_eco3047, w_eco3048, w_eco3049, w_eco3050, w_eco3051, w_eco3052, w_eco3053, w_eco3054, w_eco3055, w_eco3056, w_eco3057, w_eco3058, w_eco3059, w_eco3060, w_eco3061, w_eco3062, w_eco3063, w_eco3064, w_eco3065, w_eco3066, w_eco3067, w_eco3068, w_eco3069, w_eco3070, w_eco3071, w_eco3072, w_eco3073, w_eco3074, w_eco3075, w_eco3076, w_eco3077, w_eco3078, w_eco3079, w_eco3080, w_eco3081, w_eco3082, w_eco3083, w_eco3084, w_eco3085, w_eco3086, w_eco3087, w_eco3088, w_eco3089, w_eco3090, w_eco3091, w_eco3092, w_eco3093, w_eco3094, w_eco3095, w_eco3096, w_eco3097, w_eco3098, w_eco3099, w_eco3100, w_eco3101, w_eco3102, w_eco3103, w_eco3104, w_eco3105, w_eco3106, w_eco3107, w_eco3108, w_eco3109, w_eco3110, w_eco3111, w_eco3112, w_eco3113, w_eco3114, w_eco3115, w_eco3116, w_eco3117, w_eco3118, w_eco3119, w_eco3120, w_eco3121, w_eco3122, w_eco3123, w_eco3124, w_eco3125, w_eco3126, w_eco3127, w_eco3128, w_eco3129, w_eco3130, w_eco3131, w_eco3132, w_eco3133, w_eco3134, w_eco3135, w_eco3136, w_eco3137, w_eco3138, w_eco3139, w_eco3140, w_eco3141, w_eco3142, w_eco3143, w_eco3144, w_eco3145, w_eco3146, w_eco3147, w_eco3148, w_eco3149, w_eco3150, w_eco3151, w_eco3152, w_eco3153, w_eco3154, w_eco3155, w_eco3156, w_eco3157, w_eco3158, w_eco3159, w_eco3160, w_eco3161, w_eco3162, w_eco3163, w_eco3164, w_eco3165, w_eco3166, w_eco3167, w_eco3168, w_eco3169, w_eco3170, w_eco3171, w_eco3172, w_eco3173, w_eco3174, w_eco3175, w_eco3176, w_eco3177, w_eco3178, w_eco3179, w_eco3180, w_eco3181, w_eco3182, w_eco3183, w_eco3184, w_eco3185, w_eco3186, w_eco3187, w_eco3188, w_eco3189, w_eco3190, w_eco3191, w_eco3192, w_eco3193, w_eco3194, w_eco3195, w_eco3196, w_eco3197, w_eco3198, w_eco3199, w_eco3200, w_eco3201, w_eco3202, w_eco3203, w_eco3204, w_eco3205, w_eco3206, w_eco3207, w_eco3208, w_eco3209, w_eco3210, w_eco3211, w_eco3212, w_eco3213, w_eco3214, w_eco3215, w_eco3216, w_eco3217, w_eco3218, w_eco3219, w_eco3220, w_eco3221, w_eco3222, w_eco3223, w_eco3224, w_eco3225, w_eco3226, w_eco3227, w_eco3228, w_eco3229, w_eco3230, w_eco3231, w_eco3232, w_eco3233, w_eco3234, w_eco3235, w_eco3236, w_eco3237, w_eco3238, w_eco3239, w_eco3240, w_eco3241, w_eco3242, w_eco3243, w_eco3244, w_eco3245, w_eco3246, w_eco3247, w_eco3248, w_eco3249, w_eco3250, w_eco3251, w_eco3252, w_eco3253, w_eco3254, w_eco3255, w_eco3256, w_eco3257, w_eco3258, w_eco3259, w_eco3260, w_eco3261, w_eco3262, w_eco3263, w_eco3264, w_eco3265, w_eco3266, w_eco3267, w_eco3268, w_eco3269, w_eco3270, w_eco3271, w_eco3272, w_eco3273, w_eco3274, w_eco3275, w_eco3276, w_eco3277, w_eco3278, w_eco3279, w_eco3280, w_eco3281, w_eco3282, w_eco3283, w_eco3284, w_eco3285, w_eco3286, w_eco3287, w_eco3288, w_eco3289, w_eco3290, w_eco3291, w_eco3292, w_eco3293, w_eco3294, w_eco3295, w_eco3296, w_eco3297, w_eco3298, w_eco3299, w_eco3300, w_eco3301, w_eco3302, w_eco3303, w_eco3304, w_eco3305, w_eco3306, w_eco3307, w_eco3308, w_eco3309, w_eco3310, w_eco3311, w_eco3312, w_eco3313, w_eco3314, w_eco3315, w_eco3316, w_eco3317, w_eco3318, w_eco3319, w_eco3320, w_eco3321, w_eco3322, w_eco3323, w_eco3324, w_eco3325, w_eco3326, w_eco3327, w_eco3328, w_eco3329, w_eco3330, w_eco3331, w_eco3332, w_eco3333, w_eco3334, w_eco3335, w_eco3336, w_eco3337, w_eco3338, sub_wire7, w_eco3339, w_eco3340, w_eco3341, w_eco3342, w_eco3343, w_eco3344, w_eco3345, w_eco3346, w_eco3347, w_eco3348, w_eco3349, w_eco3350, w_eco3351, w_eco3352, w_eco3353, w_eco3354, w_eco3355, w_eco3356, w_eco3357, w_eco3358, w_eco3359, w_eco3360, w_eco3361, w_eco3362, w_eco3363, w_eco3364, w_eco3365, w_eco3366, w_eco3367, w_eco3368, w_eco3369, w_eco3370, w_eco3371, w_eco3372, w_eco3373, w_eco3374, w_eco3375, w_eco3376, w_eco3377, w_eco3378, w_eco3379, w_eco3380, w_eco3381, w_eco3382, w_eco3383, w_eco3384, w_eco3385, w_eco3386, w_eco3387, w_eco3388, w_eco3389, w_eco3390, w_eco3391, w_eco3392, w_eco3393, w_eco3394, w_eco3395, w_eco3396, w_eco3397, w_eco3398, w_eco3399, w_eco3400, w_eco3401, w_eco3402, w_eco3403, w_eco3404, w_eco3405, w_eco3406, w_eco3407, w_eco3408, w_eco3409, w_eco3410, w_eco3411, w_eco3412, w_eco3413, w_eco3414, w_eco3415, w_eco3416, w_eco3417, w_eco3418, w_eco3419, w_eco3420, w_eco3421, w_eco3422, w_eco3423, w_eco3424, w_eco3425, w_eco3426, w_eco3427, w_eco3428, w_eco3429, w_eco3430, w_eco3431, w_eco3432, w_eco3433, w_eco3434, w_eco3435, w_eco3436, w_eco3437, w_eco3438, w_eco3439, w_eco3440, w_eco3441, w_eco3442, w_eco3443, w_eco3444, w_eco3445, w_eco3446, w_eco3447, w_eco3448, w_eco3449, w_eco3450, w_eco3451, w_eco3452, w_eco3453, w_eco3454, w_eco3455, w_eco3456, w_eco3457, w_eco3458, w_eco3459, w_eco3460, w_eco3461, w_eco3462, w_eco3463, w_eco3464, w_eco3465, w_eco3466, w_eco3467, w_eco3468, w_eco3469, w_eco3470, w_eco3471, w_eco3472, w_eco3473, w_eco3474, w_eco3475, w_eco3476, w_eco3477, w_eco3478, w_eco3479, w_eco3480, w_eco3481, w_eco3482, w_eco3483, w_eco3484, w_eco3485, w_eco3486, w_eco3487, w_eco3488, w_eco3489, w_eco3490, w_eco3491, w_eco3492, w_eco3493, w_eco3494, w_eco3495, w_eco3496, w_eco3497, w_eco3498, w_eco3499, w_eco3500, w_eco3501, w_eco3502, w_eco3503, w_eco3504, w_eco3505, w_eco3506, w_eco3507, w_eco3508, w_eco3509, w_eco3510, w_eco3511, w_eco3512, w_eco3513, w_eco3514, w_eco3515, w_eco3516, w_eco3517, w_eco3518, w_eco3519, w_eco3520, w_eco3521, w_eco3522, w_eco3523, w_eco3524, w_eco3525, w_eco3526, w_eco3527, w_eco3528, w_eco3529, w_eco3530, w_eco3531, w_eco3532, w_eco3533, w_eco3534, w_eco3535, w_eco3536, w_eco3537, w_eco3538, w_eco3539, w_eco3540, w_eco3541, w_eco3542, w_eco3543, w_eco3544, w_eco3545, w_eco3546, w_eco3547, w_eco3548, w_eco3549, w_eco3550, w_eco3551, w_eco3552, w_eco3553, w_eco3554, w_eco3555, w_eco3556, w_eco3557, w_eco3558, w_eco3559, w_eco3560, w_eco3561, w_eco3562, w_eco3563, w_eco3564, w_eco3565, w_eco3566, w_eco3567, w_eco3568, w_eco3569, w_eco3570, w_eco3571, w_eco3572, w_eco3573, w_eco3574, w_eco3575, w_eco3576, w_eco3577, w_eco3578, w_eco3579, w_eco3580, w_eco3581, w_eco3582, w_eco3583, w_eco3584, w_eco3585, w_eco3586, w_eco3587, w_eco3588, w_eco3589, w_eco3590, w_eco3591, w_eco3592, w_eco3593, w_eco3594, w_eco3595, w_eco3596, w_eco3597, w_eco3598, w_eco3599, w_eco3600, w_eco3601, w_eco3602, w_eco3603, w_eco3604, w_eco3605, w_eco3606, w_eco3607, w_eco3608, w_eco3609, w_eco3610, w_eco3611, w_eco3612, w_eco3613, w_eco3614, w_eco3615, w_eco3616, w_eco3617, w_eco3618, w_eco3619, w_eco3620, w_eco3621, w_eco3622, w_eco3623, w_eco3624, w_eco3625, w_eco3626, w_eco3627, w_eco3628, w_eco3629, w_eco3630, w_eco3631, w_eco3632, w_eco3633, w_eco3634, w_eco3635, w_eco3636, w_eco3637, w_eco3638, w_eco3639, w_eco3640, w_eco3641, w_eco3642, w_eco3643, w_eco3644, w_eco3645, w_eco3646, w_eco3647, w_eco3648, w_eco3649, w_eco3650, w_eco3651, w_eco3652, w_eco3653, w_eco3654, w_eco3655, w_eco3656, w_eco3657, w_eco3658, w_eco3659, w_eco3660, w_eco3661, w_eco3662, w_eco3663, w_eco3664, w_eco3665, w_eco3666, w_eco3667, w_eco3668, w_eco3669, w_eco3670, w_eco3671, w_eco3672, w_eco3673, w_eco3674, w_eco3675, w_eco3676, w_eco3677, w_eco3678, w_eco3679, w_eco3680, w_eco3681, w_eco3682, w_eco3683, w_eco3684, w_eco3685, w_eco3686, w_eco3687, w_eco3688, w_eco3689, w_eco3690, w_eco3691, w_eco3692, w_eco3693, w_eco3694, w_eco3695, w_eco3696, w_eco3697, w_eco3698, w_eco3699, w_eco3700, w_eco3701, w_eco3702, w_eco3703, w_eco3704, w_eco3705, w_eco3706, w_eco3707, w_eco3708, w_eco3709, w_eco3710, w_eco3711, w_eco3712, w_eco3713, w_eco3714, w_eco3715, w_eco3716, w_eco3717, w_eco3718, w_eco3719, w_eco3720, w_eco3721, w_eco3722, w_eco3723, w_eco3724, w_eco3725, w_eco3726, w_eco3727, w_eco3728, w_eco3729, w_eco3730, w_eco3731, w_eco3732, w_eco3733, w_eco3734, w_eco3735, w_eco3736, w_eco3737, w_eco3738, w_eco3739, w_eco3740, w_eco3741, w_eco3742, w_eco3743, w_eco3744, w_eco3745, w_eco3746, w_eco3747, w_eco3748, w_eco3749, w_eco3750, w_eco3751, w_eco3752, w_eco3753, w_eco3754, w_eco3755, w_eco3756, w_eco3757, w_eco3758, w_eco3759, w_eco3760, w_eco3761, w_eco3762, w_eco3763, w_eco3764, w_eco3765, w_eco3766, w_eco3767, w_eco3768, w_eco3769, w_eco3770, w_eco3771, w_eco3772, w_eco3773, w_eco3774, w_eco3775, w_eco3776, w_eco3777, w_eco3778, w_eco3779, w_eco3780, w_eco3781, w_eco3782, w_eco3783, w_eco3784, w_eco3785, w_eco3786, w_eco3787, w_eco3788, w_eco3789, w_eco3790, w_eco3791, w_eco3792, w_eco3793, w_eco3794, w_eco3795, w_eco3796, w_eco3797, w_eco3798, w_eco3799, w_eco3800, w_eco3801, w_eco3802, w_eco3803, w_eco3804, w_eco3805, w_eco3806, w_eco3807, w_eco3808, w_eco3809, w_eco3810, w_eco3811, w_eco3812, w_eco3813, w_eco3814, w_eco3815, w_eco3816, w_eco3817, w_eco3818, w_eco3819, w_eco3820, w_eco3821, w_eco3822, w_eco3823, w_eco3824, w_eco3825, w_eco3826, w_eco3827, w_eco3828, w_eco3829, w_eco3830, w_eco3831, w_eco3832, w_eco3833, w_eco3834, w_eco3835, w_eco3836, w_eco3837, w_eco3838, w_eco3839, w_eco3840, w_eco3841, w_eco3842, w_eco3843, w_eco3844, w_eco3845, w_eco3846, w_eco3847, w_eco3848, w_eco3849, w_eco3850, w_eco3851, w_eco3852, w_eco3853, w_eco3854, w_eco3855, w_eco3856, w_eco3857, w_eco3858, w_eco3859, w_eco3860, w_eco3861, w_eco3862, w_eco3863, w_eco3864, w_eco3865, w_eco3866, w_eco3867, w_eco3868, w_eco3869, w_eco3870, w_eco3871, w_eco3872, w_eco3873, w_eco3874, w_eco3875, w_eco3876, w_eco3877, w_eco3878, w_eco3879, w_eco3880, w_eco3881, w_eco3882, w_eco3883, w_eco3884, w_eco3885, w_eco3886, w_eco3887, w_eco3888, w_eco3889, w_eco3890, w_eco3891, w_eco3892, w_eco3893, w_eco3894, w_eco3895, w_eco3896, w_eco3897, w_eco3898, w_eco3899, w_eco3900, w_eco3901, w_eco3902, w_eco3903, w_eco3904, w_eco3905, w_eco3906, w_eco3907, w_eco3908, w_eco3909, w_eco3910, w_eco3911, w_eco3912, w_eco3913, w_eco3914, w_eco3915, w_eco3916, w_eco3917, w_eco3918, w_eco3919, w_eco3920, w_eco3921, w_eco3922, w_eco3923, w_eco3924, w_eco3925, w_eco3926, w_eco3927, w_eco3928, w_eco3929, w_eco3930, w_eco3931, w_eco3932, w_eco3933, w_eco3934, w_eco3935, w_eco3936, w_eco3937, w_eco3938, w_eco3939, w_eco3940, w_eco3941, w_eco3942, w_eco3943, w_eco3944, w_eco3945, w_eco3946, w_eco3947, w_eco3948, w_eco3949, w_eco3950, w_eco3951, w_eco3952, w_eco3953, w_eco3954, w_eco3955, w_eco3956, w_eco3957, w_eco3958, w_eco3959, w_eco3960, w_eco3961, w_eco3962, w_eco3963, w_eco3964, w_eco3965, w_eco3966, w_eco3967, w_eco3968, w_eco3969, w_eco3970, w_eco3971, w_eco3972, w_eco3973, w_eco3974, w_eco3975, w_eco3976, w_eco3977, w_eco3978, w_eco3979, w_eco3980, w_eco3981, w_eco3982, w_eco3983, w_eco3984, w_eco3985, w_eco3986, w_eco3987, w_eco3988, w_eco3989, w_eco3990, w_eco3991, w_eco3992, w_eco3993, w_eco3994, w_eco3995, w_eco3996, w_eco3997, w_eco3998, w_eco3999, w_eco4000, w_eco4001, w_eco4002, w_eco4003, w_eco4004, w_eco4005, w_eco4006, w_eco4007, w_eco4008, w_eco4009, w_eco4010, w_eco4011, w_eco4012, w_eco4013, w_eco4014, w_eco4015, w_eco4016, w_eco4017, w_eco4018, w_eco4019, w_eco4020, w_eco4021, w_eco4022, w_eco4023, w_eco4024, w_eco4025, w_eco4026, w_eco4027, w_eco4028, w_eco4029, w_eco4030, w_eco4031, w_eco4032, w_eco4033, w_eco4034, w_eco4035, w_eco4036, w_eco4037, w_eco4038, w_eco4039, w_eco4040, w_eco4041, w_eco4042, w_eco4043, w_eco4044, w_eco4045, w_eco4046, w_eco4047, w_eco4048, w_eco4049, w_eco4050, w_eco4051, w_eco4052, w_eco4053, w_eco4054, w_eco4055, w_eco4056, w_eco4057, w_eco4058, w_eco4059, w_eco4060, w_eco4061, w_eco4062, w_eco4063, w_eco4064, w_eco4065, w_eco4066, w_eco4067, w_eco4068, w_eco4069, w_eco4070, w_eco4071, w_eco4072, w_eco4073, w_eco4074, w_eco4075, w_eco4076, w_eco4077, w_eco4078, w_eco4079, w_eco4080, w_eco4081, w_eco4082, w_eco4083, w_eco4084, w_eco4085, w_eco4086, w_eco4087, w_eco4088, w_eco4089, w_eco4090, w_eco4091, w_eco4092, w_eco4093, w_eco4094, w_eco4095, w_eco4096, w_eco4097, w_eco4098, w_eco4099, w_eco4100, w_eco4101, w_eco4102, w_eco4103, w_eco4104, w_eco4105, w_eco4106, w_eco4107, w_eco4108, w_eco4109, w_eco4110, w_eco4111, w_eco4112, w_eco4113, w_eco4114, w_eco4115, w_eco4116, w_eco4117, w_eco4118, w_eco4119, w_eco4120, w_eco4121, w_eco4122, w_eco4123, w_eco4124, w_eco4125, w_eco4126, w_eco4127, w_eco4128, w_eco4129, w_eco4130, w_eco4131, w_eco4132, w_eco4133, w_eco4134, w_eco4135, w_eco4136, w_eco4137, w_eco4138, w_eco4139, w_eco4140, w_eco4141, w_eco4142, w_eco4143, w_eco4144, w_eco4145, w_eco4146, w_eco4147, w_eco4148, w_eco4149, w_eco4150, w_eco4151, w_eco4152, w_eco4153, w_eco4154, w_eco4155, w_eco4156, w_eco4157, w_eco4158, w_eco4159, w_eco4160, w_eco4161, w_eco4162, w_eco4163, w_eco4164, w_eco4165, w_eco4166, w_eco4167, w_eco4168, w_eco4169, w_eco4170, w_eco4171, w_eco4172, w_eco4173, w_eco4174, w_eco4175, w_eco4176, w_eco4177, w_eco4178, w_eco4179, w_eco4180, w_eco4181, w_eco4182, w_eco4183, w_eco4184, w_eco4185, w_eco4186, w_eco4187, w_eco4188, w_eco4189, w_eco4190, w_eco4191, w_eco4192, w_eco4193, w_eco4194, w_eco4195, w_eco4196, w_eco4197, w_eco4198, w_eco4199, w_eco4200, w_eco4201, w_eco4202, w_eco4203, w_eco4204, w_eco4205, w_eco4206, w_eco4207, w_eco4208, w_eco4209, w_eco4210, w_eco4211, w_eco4212, w_eco4213, w_eco4214, w_eco4215, w_eco4216, w_eco4217, w_eco4218, w_eco4219, w_eco4220, w_eco4221, w_eco4222, w_eco4223, w_eco4224, w_eco4225, w_eco4226, w_eco4227, w_eco4228, w_eco4229, w_eco4230, w_eco4231, w_eco4232, w_eco4233, w_eco4234, w_eco4235, w_eco4236, w_eco4237, w_eco4238, w_eco4239, w_eco4240, w_eco4241, w_eco4242, w_eco4243, w_eco4244, w_eco4245, w_eco4246, w_eco4247, w_eco4248, w_eco4249, w_eco4250, w_eco4251, w_eco4252, w_eco4253, w_eco4254, w_eco4255, w_eco4256, w_eco4257, w_eco4258, w_eco4259, w_eco4260, w_eco4261, w_eco4262, w_eco4263, w_eco4264, w_eco4265, w_eco4266, w_eco4267, w_eco4268, w_eco4269, w_eco4270, w_eco4271, w_eco4272, w_eco4273, w_eco4274, w_eco4275, w_eco4276, w_eco4277, w_eco4278, w_eco4279, w_eco4280, w_eco4281, w_eco4282, w_eco4283, w_eco4284, w_eco4285, sub_wire8, w_eco4286, w_eco4287, w_eco4288, w_eco4289, w_eco4290, w_eco4291, w_eco4292, w_eco4293, w_eco4294, w_eco4295, w_eco4296, w_eco4297, w_eco4298, w_eco4299, w_eco4300, w_eco4301, w_eco4302, w_eco4303, w_eco4304, w_eco4305, w_eco4306, w_eco4307, w_eco4308, w_eco4309, w_eco4310, w_eco4311, w_eco4312, w_eco4313, w_eco4314, w_eco4315, w_eco4316, w_eco4317, w_eco4318, w_eco4319, w_eco4320, w_eco4321, w_eco4322, w_eco4323, w_eco4324, w_eco4325, w_eco4326, w_eco4327, w_eco4328, w_eco4329, w_eco4330, w_eco4331, w_eco4332, w_eco4333, w_eco4334, w_eco4335, w_eco4336, w_eco4337, w_eco4338, w_eco4339, w_eco4340, w_eco4341, w_eco4342, w_eco4343, w_eco4344, w_eco4345, w_eco4346, w_eco4347, w_eco4348, w_eco4349, w_eco4350, w_eco4351, w_eco4352, w_eco4353, w_eco4354, w_eco4355, w_eco4356, w_eco4357, w_eco4358, w_eco4359, w_eco4360, w_eco4361, w_eco4362, w_eco4363, w_eco4364, w_eco4365, w_eco4366, w_eco4367, w_eco4368, w_eco4369, w_eco4370, w_eco4371, w_eco4372, w_eco4373, w_eco4374, w_eco4375, w_eco4376, w_eco4377, w_eco4378, w_eco4379, w_eco4380, w_eco4381, w_eco4382, w_eco4383, w_eco4384, w_eco4385, w_eco4386, w_eco4387, w_eco4388, w_eco4389, w_eco4390, w_eco4391, w_eco4392, w_eco4393, w_eco4394, w_eco4395, w_eco4396, w_eco4397, w_eco4398, w_eco4399, w_eco4400, w_eco4401, w_eco4402, w_eco4403, w_eco4404, w_eco4405, w_eco4406, w_eco4407, w_eco4408, w_eco4409, w_eco4410, w_eco4411, w_eco4412, w_eco4413, w_eco4414, w_eco4415, w_eco4416, w_eco4417, w_eco4418, w_eco4419, w_eco4420, w_eco4421, w_eco4422, w_eco4423, w_eco4424, w_eco4425, w_eco4426, w_eco4427, w_eco4428, w_eco4429, w_eco4430, w_eco4431, w_eco4432, w_eco4433, w_eco4434, w_eco4435, w_eco4436, w_eco4437, w_eco4438, w_eco4439, w_eco4440, w_eco4441, w_eco4442, w_eco4443, w_eco4444, w_eco4445, w_eco4446, w_eco4447, w_eco4448, w_eco4449, w_eco4450, w_eco4451, w_eco4452, w_eco4453, w_eco4454, w_eco4455, w_eco4456, w_eco4457, w_eco4458, w_eco4459, w_eco4460, w_eco4461, w_eco4462, w_eco4463, w_eco4464, w_eco4465, w_eco4466, w_eco4467, w_eco4468, w_eco4469, w_eco4470, w_eco4471, w_eco4472, w_eco4473, w_eco4474, w_eco4475, w_eco4476, w_eco4477, w_eco4478, w_eco4479, w_eco4480, w_eco4481, w_eco4482, w_eco4483, w_eco4484, w_eco4485, w_eco4486, w_eco4487, w_eco4488, w_eco4489, w_eco4490, w_eco4491, w_eco4492, w_eco4493, w_eco4494, w_eco4495, w_eco4496, w_eco4497, w_eco4498, w_eco4499, w_eco4500, w_eco4501, w_eco4502, w_eco4503, w_eco4504, w_eco4505, w_eco4506, w_eco4507, w_eco4508, w_eco4509, w_eco4510, w_eco4511, w_eco4512, w_eco4513, w_eco4514, w_eco4515, w_eco4516, w_eco4517, w_eco4518, w_eco4519, w_eco4520, w_eco4521, w_eco4522, w_eco4523, w_eco4524, w_eco4525, w_eco4526, w_eco4527, w_eco4528, w_eco4529, w_eco4530, w_eco4531, w_eco4532, w_eco4533, w_eco4534, w_eco4535, w_eco4536, w_eco4537, w_eco4538, w_eco4539, w_eco4540, w_eco4541, w_eco4542, w_eco4543, w_eco4544, w_eco4545, w_eco4546, w_eco4547, w_eco4548, w_eco4549, w_eco4550, w_eco4551, w_eco4552, w_eco4553, w_eco4554, w_eco4555, w_eco4556, w_eco4557, w_eco4558, w_eco4559, w_eco4560, w_eco4561, w_eco4562, w_eco4563, w_eco4564, w_eco4565, w_eco4566, w_eco4567, w_eco4568, w_eco4569, w_eco4570, w_eco4571, w_eco4572, w_eco4573, w_eco4574, w_eco4575, w_eco4576, w_eco4577, w_eco4578, w_eco4579, w_eco4580, w_eco4581, w_eco4582, w_eco4583, w_eco4584, w_eco4585, w_eco4586, w_eco4587, w_eco4588, w_eco4589, w_eco4590, w_eco4591, w_eco4592, w_eco4593, w_eco4594, w_eco4595, w_eco4596, w_eco4597, w_eco4598, w_eco4599, w_eco4600, w_eco4601, w_eco4602, w_eco4603, w_eco4604, w_eco4605, w_eco4606, w_eco4607, w_eco4608, w_eco4609, w_eco4610, w_eco4611, w_eco4612, w_eco4613, w_eco4614, w_eco4615, w_eco4616, w_eco4617, w_eco4618, w_eco4619, w_eco4620, w_eco4621, w_eco4622, w_eco4623, w_eco4624, w_eco4625, w_eco4626, w_eco4627, w_eco4628, w_eco4629, w_eco4630, w_eco4631, w_eco4632, w_eco4633, w_eco4634, w_eco4635, w_eco4636, w_eco4637, w_eco4638, w_eco4639, w_eco4640, w_eco4641, w_eco4642, w_eco4643, w_eco4644, w_eco4645, w_eco4646, w_eco4647, w_eco4648, w_eco4649, w_eco4650, w_eco4651, w_eco4652, w_eco4653, w_eco4654, w_eco4655, w_eco4656, w_eco4657, w_eco4658, w_eco4659, w_eco4660, w_eco4661, w_eco4662, w_eco4663, w_eco4664, w_eco4665, w_eco4666, w_eco4667, w_eco4668, w_eco4669, w_eco4670, w_eco4671, w_eco4672, w_eco4673, w_eco4674, w_eco4675, w_eco4676, w_eco4677, w_eco4678, w_eco4679, w_eco4680, w_eco4681, w_eco4682, w_eco4683, w_eco4684, w_eco4685, w_eco4686, w_eco4687, w_eco4688, w_eco4689, w_eco4690, w_eco4691, w_eco4692, w_eco4693, w_eco4694, w_eco4695, w_eco4696, w_eco4697, w_eco4698, w_eco4699, w_eco4700, w_eco4701, w_eco4702, w_eco4703, w_eco4704, w_eco4705, w_eco4706, w_eco4707, w_eco4708, w_eco4709, w_eco4710, w_eco4711, w_eco4712, w_eco4713, w_eco4714, w_eco4715, w_eco4716, w_eco4717, w_eco4718, w_eco4719, w_eco4720, w_eco4721, w_eco4722, w_eco4723, w_eco4724, w_eco4725, w_eco4726, w_eco4727, w_eco4728, w_eco4729, w_eco4730, w_eco4731, w_eco4732, w_eco4733, w_eco4734, w_eco4735, w_eco4736, w_eco4737, w_eco4738, w_eco4739, w_eco4740, w_eco4741, w_eco4742, w_eco4743, w_eco4744, w_eco4745, w_eco4746, w_eco4747, w_eco4748, w_eco4749, w_eco4750, w_eco4751, w_eco4752, w_eco4753, w_eco4754, w_eco4755, w_eco4756, w_eco4757, w_eco4758, w_eco4759, w_eco4760, w_eco4761, w_eco4762, w_eco4763, w_eco4764, w_eco4765, w_eco4766, w_eco4767, w_eco4768, w_eco4769, w_eco4770, w_eco4771, w_eco4772, w_eco4773, w_eco4774, w_eco4775, w_eco4776, w_eco4777, w_eco4778, w_eco4779, w_eco4780, w_eco4781, w_eco4782, w_eco4783, w_eco4784, w_eco4785, w_eco4786, w_eco4787, w_eco4788, w_eco4789, w_eco4790, w_eco4791, w_eco4792, w_eco4793, w_eco4794, w_eco4795, w_eco4796, w_eco4797, w_eco4798, w_eco4799, w_eco4800, w_eco4801, w_eco4802, w_eco4803, w_eco4804, w_eco4805, w_eco4806, w_eco4807, w_eco4808, w_eco4809, w_eco4810, w_eco4811, w_eco4812, w_eco4813, w_eco4814, w_eco4815, w_eco4816, w_eco4817, w_eco4818, w_eco4819, w_eco4820, w_eco4821, w_eco4822, w_eco4823, w_eco4824, w_eco4825, w_eco4826, w_eco4827, w_eco4828, w_eco4829, w_eco4830, w_eco4831, w_eco4832, w_eco4833, w_eco4834, w_eco4835, w_eco4836, w_eco4837, w_eco4838, w_eco4839, w_eco4840, w_eco4841, w_eco4842, w_eco4843, w_eco4844, w_eco4845, w_eco4846, w_eco4847, w_eco4848, w_eco4849, w_eco4850, w_eco4851, w_eco4852, w_eco4853, w_eco4854, w_eco4855, w_eco4856, w_eco4857, w_eco4858, w_eco4859, w_eco4860, w_eco4861, w_eco4862, w_eco4863, w_eco4864, w_eco4865, w_eco4866, w_eco4867, w_eco4868, w_eco4869, w_eco4870, w_eco4871, w_eco4872, w_eco4873, w_eco4874, w_eco4875, w_eco4876, w_eco4877, w_eco4878, w_eco4879, w_eco4880, w_eco4881, w_eco4882, w_eco4883, w_eco4884, w_eco4885, w_eco4886, w_eco4887, w_eco4888, w_eco4889, w_eco4890, w_eco4891, w_eco4892, w_eco4893, w_eco4894, w_eco4895, w_eco4896, w_eco4897, w_eco4898, w_eco4899, w_eco4900, w_eco4901, w_eco4902, w_eco4903, w_eco4904, w_eco4905, w_eco4906, w_eco4907, w_eco4908, w_eco4909, w_eco4910, w_eco4911, w_eco4912, w_eco4913, w_eco4914, w_eco4915, w_eco4916, w_eco4917, w_eco4918, w_eco4919, w_eco4920, w_eco4921, w_eco4922, w_eco4923, w_eco4924, w_eco4925, w_eco4926, w_eco4927, w_eco4928, w_eco4929, w_eco4930, w_eco4931, w_eco4932, w_eco4933, w_eco4934, w_eco4935, w_eco4936, w_eco4937, w_eco4938, w_eco4939, w_eco4940, w_eco4941, w_eco4942, w_eco4943, w_eco4944, w_eco4945, w_eco4946, w_eco4947, w_eco4948, w_eco4949, w_eco4950, w_eco4951, w_eco4952, w_eco4953, w_eco4954, w_eco4955, w_eco4956, w_eco4957, w_eco4958, w_eco4959, w_eco4960, w_eco4961, w_eco4962, w_eco4963, w_eco4964, w_eco4965, w_eco4966, w_eco4967, w_eco4968, w_eco4969, w_eco4970, w_eco4971, w_eco4972, w_eco4973, w_eco4974, w_eco4975, w_eco4976, w_eco4977, w_eco4978, w_eco4979, w_eco4980, w_eco4981, w_eco4982, w_eco4983, w_eco4984, w_eco4985, w_eco4986, w_eco4987, w_eco4988, w_eco4989, w_eco4990, w_eco4991, w_eco4992, w_eco4993, w_eco4994, w_eco4995, w_eco4996, w_eco4997, w_eco4998, w_eco4999, w_eco5000, w_eco5001, w_eco5002, w_eco5003, w_eco5004, w_eco5005, w_eco5006, w_eco5007, w_eco5008, w_eco5009, w_eco5010, w_eco5011, w_eco5012, w_eco5013, w_eco5014, w_eco5015, w_eco5016, w_eco5017, w_eco5018, w_eco5019, w_eco5020, w_eco5021, w_eco5022, w_eco5023, w_eco5024, w_eco5025, w_eco5026, w_eco5027, w_eco5028, w_eco5029, w_eco5030, w_eco5031, w_eco5032, w_eco5033, w_eco5034, w_eco5035, w_eco5036, w_eco5037, w_eco5038, w_eco5039, w_eco5040, w_eco5041, w_eco5042, w_eco5043, w_eco5044, w_eco5045, w_eco5046, w_eco5047, w_eco5048, w_eco5049, w_eco5050, w_eco5051, w_eco5052, w_eco5053, w_eco5054, w_eco5055, w_eco5056, w_eco5057, w_eco5058, w_eco5059, w_eco5060, w_eco5061, w_eco5062, w_eco5063, w_eco5064, w_eco5065, w_eco5066, w_eco5067, w_eco5068, w_eco5069, w_eco5070, w_eco5071, w_eco5072, w_eco5073, w_eco5074, w_eco5075, w_eco5076, w_eco5077, w_eco5078, w_eco5079, w_eco5080, w_eco5081, w_eco5082, sub_wire9, w_eco5083, w_eco5084, w_eco5085, w_eco5086, w_eco5087, w_eco5088, w_eco5089, w_eco5090, w_eco5091, w_eco5092, w_eco5093, w_eco5094, w_eco5095, w_eco5096, w_eco5097, w_eco5098, w_eco5099, w_eco5100, w_eco5101, w_eco5102, w_eco5103, w_eco5104, w_eco5105, w_eco5106, w_eco5107, w_eco5108, w_eco5109, w_eco5110, w_eco5111, w_eco5112, w_eco5113, w_eco5114, w_eco5115, w_eco5116, w_eco5117, w_eco5118, w_eco5119, w_eco5120, w_eco5121, w_eco5122, w_eco5123, w_eco5124, w_eco5125, w_eco5126, w_eco5127, w_eco5128, w_eco5129, w_eco5130, w_eco5131, w_eco5132, w_eco5133, w_eco5134, w_eco5135, w_eco5136, w_eco5137, w_eco5138, w_eco5139, w_eco5140, w_eco5141, w_eco5142, w_eco5143, w_eco5144, w_eco5145, w_eco5146, w_eco5147, w_eco5148, w_eco5149, w_eco5150, w_eco5151, w_eco5152, w_eco5153, w_eco5154, w_eco5155, w_eco5156, w_eco5157, w_eco5158, w_eco5159, w_eco5160, w_eco5161, w_eco5162, w_eco5163, w_eco5164, w_eco5165, w_eco5166, w_eco5167, w_eco5168, w_eco5169, w_eco5170, w_eco5171, w_eco5172, w_eco5173, w_eco5174, w_eco5175, w_eco5176, w_eco5177, w_eco5178, w_eco5179, w_eco5180, w_eco5181, w_eco5182, w_eco5183, w_eco5184, w_eco5185, w_eco5186, w_eco5187, w_eco5188, w_eco5189, w_eco5190, w_eco5191, w_eco5192, w_eco5193, w_eco5194, w_eco5195, w_eco5196, w_eco5197, w_eco5198, w_eco5199, w_eco5200, w_eco5201, w_eco5202, w_eco5203, w_eco5204, w_eco5205, w_eco5206, w_eco5207, w_eco5208, w_eco5209, w_eco5210, w_eco5211, w_eco5212, w_eco5213, w_eco5214, w_eco5215, w_eco5216, w_eco5217, w_eco5218, w_eco5219, w_eco5220, w_eco5221, w_eco5222, w_eco5223, w_eco5224, w_eco5225, w_eco5226, w_eco5227, w_eco5228, w_eco5229, w_eco5230, w_eco5231, w_eco5232, w_eco5233, w_eco5234, w_eco5235, w_eco5236, w_eco5237, w_eco5238, w_eco5239, w_eco5240, w_eco5241, w_eco5242, w_eco5243, w_eco5244, w_eco5245, w_eco5246, w_eco5247, w_eco5248, w_eco5249, w_eco5250, w_eco5251, w_eco5252, w_eco5253, w_eco5254, w_eco5255, w_eco5256, w_eco5257, w_eco5258, w_eco5259, w_eco5260, w_eco5261, w_eco5262, w_eco5263, w_eco5264, w_eco5265, w_eco5266, w_eco5267, w_eco5268, w_eco5269, w_eco5270, w_eco5271, w_eco5272, w_eco5273, w_eco5274, w_eco5275, w_eco5276, w_eco5277, w_eco5278, w_eco5279, w_eco5280, w_eco5281, w_eco5282, w_eco5283, w_eco5284, w_eco5285, w_eco5286, w_eco5287, w_eco5288, w_eco5289, w_eco5290, w_eco5291, w_eco5292, w_eco5293, w_eco5294, w_eco5295, w_eco5296, w_eco5297, w_eco5298, w_eco5299, w_eco5300, w_eco5301, w_eco5302, w_eco5303, w_eco5304, w_eco5305, w_eco5306, w_eco5307, w_eco5308, w_eco5309, w_eco5310, w_eco5311, w_eco5312, w_eco5313, w_eco5314, w_eco5315, w_eco5316, w_eco5317, w_eco5318, w_eco5319, w_eco5320, w_eco5321, w_eco5322, w_eco5323, w_eco5324, w_eco5325, w_eco5326, w_eco5327, w_eco5328, w_eco5329, w_eco5330, w_eco5331, w_eco5332, w_eco5333, w_eco5334, w_eco5335, w_eco5336, w_eco5337, w_eco5338, w_eco5339, w_eco5340, w_eco5341, w_eco5342, w_eco5343, w_eco5344, w_eco5345, w_eco5346, w_eco5347, w_eco5348, w_eco5349, w_eco5350, w_eco5351, w_eco5352, w_eco5353, w_eco5354, w_eco5355, w_eco5356, w_eco5357, w_eco5358, w_eco5359, w_eco5360, w_eco5361, w_eco5362, w_eco5363, w_eco5364, w_eco5365, w_eco5366, w_eco5367, w_eco5368, w_eco5369, w_eco5370, w_eco5371, w_eco5372, w_eco5373, w_eco5374, w_eco5375, w_eco5376, w_eco5377, w_eco5378, w_eco5379, w_eco5380, w_eco5381, w_eco5382, w_eco5383, w_eco5384, w_eco5385, w_eco5386, w_eco5387, w_eco5388, w_eco5389, w_eco5390, w_eco5391, w_eco5392, w_eco5393, w_eco5394, w_eco5395, w_eco5396, w_eco5397, w_eco5398, w_eco5399, w_eco5400, w_eco5401, w_eco5402, w_eco5403, w_eco5404, w_eco5405, w_eco5406, w_eco5407, w_eco5408, w_eco5409, w_eco5410, w_eco5411, w_eco5412, w_eco5413, w_eco5414, w_eco5415, w_eco5416, w_eco5417, w_eco5418, w_eco5419, w_eco5420, w_eco5421, w_eco5422, w_eco5423, w_eco5424, w_eco5425, w_eco5426, w_eco5427, w_eco5428, w_eco5429, w_eco5430, w_eco5431, w_eco5432, w_eco5433, w_eco5434, w_eco5435, w_eco5436, w_eco5437, w_eco5438, w_eco5439, w_eco5440, w_eco5441, w_eco5442, w_eco5443, w_eco5444, w_eco5445, w_eco5446, w_eco5447, w_eco5448, w_eco5449, w_eco5450, w_eco5451, w_eco5452, w_eco5453, w_eco5454, w_eco5455, w_eco5456, w_eco5457, w_eco5458, w_eco5459, w_eco5460, w_eco5461, w_eco5462, w_eco5463, w_eco5464, w_eco5465, w_eco5466, w_eco5467, w_eco5468, w_eco5469, w_eco5470, w_eco5471, w_eco5472, w_eco5473, w_eco5474, w_eco5475, w_eco5476, w_eco5477, w_eco5478, w_eco5479, w_eco5480, w_eco5481, w_eco5482, w_eco5483, w_eco5484, w_eco5485, w_eco5486, w_eco5487, w_eco5488, w_eco5489, w_eco5490, w_eco5491, w_eco5492, w_eco5493, w_eco5494, w_eco5495, w_eco5496, w_eco5497, w_eco5498, w_eco5499, w_eco5500, w_eco5501, w_eco5502, w_eco5503, w_eco5504, w_eco5505, w_eco5506, w_eco5507, w_eco5508, w_eco5509, w_eco5510, w_eco5511, w_eco5512, w_eco5513, w_eco5514, w_eco5515, w_eco5516, w_eco5517, w_eco5518, w_eco5519, w_eco5520, w_eco5521, w_eco5522, w_eco5523, w_eco5524, w_eco5525, w_eco5526, w_eco5527, w_eco5528, w_eco5529, w_eco5530, w_eco5531, w_eco5532, w_eco5533, w_eco5534, w_eco5535, w_eco5536, w_eco5537, w_eco5538, w_eco5539, w_eco5540, w_eco5541, w_eco5542, w_eco5543, w_eco5544, w_eco5545, w_eco5546, w_eco5547, w_eco5548, w_eco5549, w_eco5550, w_eco5551, w_eco5552, w_eco5553, w_eco5554, w_eco5555, w_eco5556, w_eco5557, w_eco5558, w_eco5559, w_eco5560, w_eco5561, w_eco5562, w_eco5563, w_eco5564, w_eco5565, w_eco5566, w_eco5567, w_eco5568, w_eco5569, w_eco5570, w_eco5571, w_eco5572, w_eco5573, w_eco5574, w_eco5575, w_eco5576, w_eco5577, w_eco5578, w_eco5579, w_eco5580, w_eco5581, w_eco5582, w_eco5583, w_eco5584, w_eco5585, w_eco5586, w_eco5587, w_eco5588, w_eco5589, w_eco5590, w_eco5591, w_eco5592, w_eco5593, w_eco5594, w_eco5595, w_eco5596, w_eco5597, w_eco5598, w_eco5599, w_eco5600, w_eco5601, w_eco5602, w_eco5603, w_eco5604, w_eco5605, w_eco5606, w_eco5607, w_eco5608, w_eco5609, w_eco5610, w_eco5611, w_eco5612, w_eco5613, w_eco5614, w_eco5615, w_eco5616, w_eco5617, w_eco5618, w_eco5619, w_eco5620, w_eco5621, w_eco5622;

	//input clk(oe, 	assign \mux_44_12_g156/data0 = 0;
	or \mux_44_12_g156/org(sub_wire0, \mux_44_12_g156/w_0, \mux_44_12_g156/w_1, \mux_44_12_g156/w_2);
	and \mux_44_12_g156/a_2(\mux_44_12_g156/w_2, n_988, n_43);
	and \mux_44_12_g156/a_1(\mux_44_12_g156/w_1, n_987, n_41);
	and \mux_44_12_g156/a_0(\mux_44_12_g156/w_0, n_986, \mux_44_12_g156/data0);
	or \mux_temp_y_21_12_g792/org(n_129, \mux_temp_y_21_12_g792/w_0, \mux_temp_y_21_12_g792/w_1);
	and \mux_temp_y_21_12_g792/a_1(\mux_temp_y_21_12_g792/w_1, n_805, n_16);
	and \mux_temp_y_21_12_g792/a_0(\mux_temp_y_21_12_g792/w_0, n_318, n_1114);
	or \mux_temp_y_21_12_g19/org(n_136, \mux_temp_y_21_12_g19/w_0, \mux_temp_y_21_12_g19/w_1, \mux_temp_y_21_12_g19/w_2, \mux_temp_y_21_12_g19/w_3);
	and \mux_temp_y_21_12_g19/a_3(\mux_temp_y_21_12_g19/w_3, n_301, n_616);
	and \mux_temp_y_21_12_g19/a_2(\mux_temp_y_21_12_g19/w_2, n_318, n_35);
	and \mux_temp_y_21_12_g19/a_1(\mux_temp_y_21_12_g19/w_1, n_1095, n_34);
	and \mux_temp_y_21_12_g19/a_0(\mux_temp_y_21_12_g19/w_0, n_1111, n_33);
	or \mux_temp_y_21_12_g18/org(n_135, \mux_temp_y_21_12_g18/w_0, \mux_temp_y_21_12_g18/w_1, \mux_temp_y_21_12_g18/w_2, \mux_temp_y_21_12_g18/w_3);
	and \mux_temp_y_21_12_g18/a_3(\mux_temp_y_21_12_g18/w_3, n_301, n_615);
	and \mux_temp_y_21_12_g18/a_2(\mux_temp_y_21_12_g18/w_2, n_318, n_39);
	and \mux_temp_y_21_12_g18/a_1(\mux_temp_y_21_12_g18/w_1, n_1095, n_38);
	and \mux_temp_y_21_12_g18/a_0(\mux_temp_y_21_12_g18/w_0, n_1111, n_37);
	or \mux_temp_y_21_12_g17/org(n_133, \mux_temp_y_21_12_g17/w_0, \mux_temp_y_21_12_g17/w_1, \mux_temp_y_21_12_g17/w_2, \mux_temp_y_21_12_g17/w_3);
	and \mux_temp_y_21_12_g17/a_3(\mux_temp_y_21_12_g17/w_3, n_301, n_620);
	and \mux_temp_y_21_12_g17/a_2(\mux_temp_y_21_12_g17/w_2, n_318, n_1113);
	and \mux_temp_y_21_12_g17/a_1(\mux_temp_y_21_12_g17/w_1, n_1095, n_26);
	and \mux_temp_y_21_12_g17/a_0(\mux_temp_y_21_12_g17/w_0, n_1111, n_25);
	or \mux_temp_y_21_12_g16/org(n_132, \mux_temp_y_21_12_g16/w_0, \mux_temp_y_21_12_g16/w_1, \mux_temp_y_21_12_g16/w_2, \mux_temp_y_21_12_g16/w_3);
	and \mux_temp_y_21_12_g16/a_3(\mux_temp_y_21_12_g16/w_3, n_301, n_619);
	and \mux_temp_y_21_12_g16/a_2(\mux_temp_y_21_12_g16/w_2, n_318, n_31);
	and \mux_temp_y_21_12_g16/a_1(\mux_temp_y_21_12_g16/w_1, n_1095, n_30);
	and \mux_temp_y_21_12_g16/a_0(\mux_temp_y_21_12_g16/w_0, n_1111, n_29);
	or \mux_temp_y_21_12_g15/org(n_131, \mux_temp_y_21_12_g15/w_0, \mux_temp_y_21_12_g15/w_1, \mux_temp_y_21_12_g15/w_2, \mux_temp_y_21_12_g15/w_3);
	and \mux_temp_y_21_12_g15/a_3(\mux_temp_y_21_12_g15/w_3, n_301, n_618);
	and \mux_temp_y_21_12_g15/a_2(\mux_temp_y_21_12_g15/w_2, n_318, n_23);
	and \mux_temp_y_21_12_g15/a_1(\mux_temp_y_21_12_g15/w_1, n_1095, n_22);
	and \mux_temp_y_21_12_g15/a_0(\mux_temp_y_21_12_g15/w_0, n_1111, n_21);
	or \mux_temp_y_21_12_g10/org(n_130, \mux_temp_y_21_12_g10/w_0, \mux_temp_y_21_12_g10/w_1, \mux_temp_y_21_12_g10/w_2, \mux_temp_y_21_12_g10/w_3);
	and \mux_temp_y_21_12_g10/a_3(\mux_temp_y_21_12_g10/w_3, n_301, n_617);
	and \mux_temp_y_21_12_g10/a_2(\mux_temp_y_21_12_g10/w_2, n_318, n_19);
	and \mux_temp_y_21_12_g10/a_1(\mux_temp_y_21_12_g10/w_1, n_1095, n_18);
	and \mux_temp_y_21_12_g10/a_0(\mux_temp_y_21_12_g10/w_0, n_1111, n_17);
	nor add_24_29_g10(add_24_29_n_33, a[3], b[3]);
	nor add_24_29_g12(add_24_29_n_43, a[4], b[4]);
	nor add_24_29_g14(add_24_29_n_39, a[5], b[5]);
	nor add_24_29_g16(add_24_29_n_50, a[6], b[6]);
	nor add_24_29_g23(add_24_29_n_48, n_880, n_1113);
	nor add_24_29_g24(add_24_29_n_47, add_24_29_n_37, add_24_29_n_33);
	nor add_24_29_g27(add_24_29_n_51, n_884, n_35);
	nor add_24_29_g28(add_24_29_n_55, add_24_29_n_43, add_24_29_n_39);
	nand add_24_29_g32(add_24_29_n_49, add_24_29_n_47, add_24_29_n_1115);
	nand add_24_29_g33(add_24_29_n_57, add_24_29_n_48, add_24_29_n_49);
	nor add_24_29_g34(add_24_29_n_53, add_24_29_n_50, add_24_29_n_51);
	xnor add_24_29_g48(n_17, n_1114, n_965);
	xnor add_24_29_g50(n_21, add_24_29_n_1115, n_966);
	xnor add_24_29_g53(n_25, n_972, n_970);
	xnor add_24_29_g55(n_29, add_24_29_n_57, n_969);
	xnor add_24_29_g58(n_33, n_979, n_968);
	nor add_24_29_g6(add_24_29_n_27, a[1], b[1]);
	xnor add_24_29_g60(n_37, n_978, n_967);
	nor add_24_29_g8(add_24_29_n_37, a[2], b[2]);
	xor g15(n_16, a[0], b[0]);
	xor g21(n_74, n_129, n_135);
	xor g22(n_75, n_136, n_130);
	xor g23(n_76, n_131, n_73);
	xor g24(n_77, n_74, n_75);
	xor g25(parity, n_76, n_77);
	xor g3(n_73, n_132, n_133);
	not gt_39_12_g10(greater, n_840);
	nand sub_29_29_g38(sub_29_29_n_54, sub_29_29_n_320, n_1104);
	nand sub_29_29_g46(sub_29_29_n_69, sub_29_29_n_63, n_300);
	xnor sub_29_29_g56(n_18, sub_29_29_n_37, n_617);
	xnor sub_29_29_g58(n_22, sub_29_29_n_320, n_618);
	xnor sub_29_29_g61(n_26, n_977, n_620);
	xnor sub_29_29_g63(n_30, sub_29_29_n_1105, n_619);
	xnor sub_29_29_g66(n_34, n_985, n_616);
	xnor sub_29_29_g68(n_38, n_984, n_615);
	not sub_29_29_g9(n_43, sub_29_29_n_32);
	nor g251(n_395, n_916, n_1096, gt_39_12_n_57);
	nor g287(n_419, n_1102, a[0]);
	nor g298(n_429, n_1096, gt_39_12_n_57, n_397);
	nor g299(n_428, gt_39_12_n_57, n_323, n_397);
	nor g303(n_431, n_1104, gt_39_12_n_46);
	not g793(n_805, n_318);
	not g904(n_872, a[7]);
	not g907(n_875, add_24_29_n_33);
	not g915(n_881, n_1113);
	not g916(n_882, add_24_29_n_37);
	not g931(n_891, gt_39_12_n_52);
	not g933(n_892, n_308);
	nor g936(gt_39_12_n_57, n_872, b[7]);
	not g937(n_894, gt_39_12_n_57);
	nand g938(n_895, n_891, n_892, n_1097, n_894);
	not g942(n_897, n_431);
	not g949(n_901, n_419);
	nor g952(n_903, n_1102, n_871);
	not g953(n_904, n_903);
	nand g954(n_905, n_901, sub_29_29_n_1103, n_904);
	nand g955(n_906, n_1098, n_1101, n_905);
	nand g956(n_907, n_897, n_1099, n_906);
	not g957(n_908, n_907);
	nor g958(n_909, n_895, n_908);
	not g959(n_910, n_909);
	not g965(n_913, sub_29_29_n_63);
	nor g966(n_914, n_891, n_911);
	not g967(n_915, n_914);
	nand g968(n_916, n_913, n_915);
	nand g971(n_323, n_872, b[7]);
	not g972(n_918, n_323);
	nor g973(n_919, n_395, n_917, n_918);
	not g974(n_920, n_919);
	nor g975(n_921, n_395, n_894, n_918);
	not g976(n_922, n_921);
	nand g977(n_923, n_920, n_922);
	nand g978(n_840, n_910, n_923);
	not g985(n_928, sub_29_29_n_69);
	nor g992(n_397, n_918, n_932);
	not g993(n_933, n_429);
	not g994(n_934, n_428);
	nand g995(n_367, n_933, n_934);
	not g996(n_935, n_367);
	nor g997(n_936, greater, n_367);
	not g998(n_937, n_936);
	nand g1004(n_379, n_928, n_323, sub_29_29_n_1105);
	not g1005(n_942, n_379);
	nor g1006(n_943, greater, n_379);
	not g1007(n_944, n_943);
	nand g1008(is_eq, n_937, n_944);
	nor g1009(sub_wire1, greater, n_935, n_942);
	nor g1036(n_318, n_1123, op[0]);
	nor g1037(n_301, n_1123, n_869);
	nand g1038(n_965, n_888, n_887);
	nand g1039(n_966, n_882, n_1112);
	nand g1041(n_615, n_300, n_1097);
	nand g1043(n_616, n_891, n_298);
	nand g1044(n_617, n_900, sub_29_29_n_1103);
	nand g1045(n_618, n_1101, n_1104);
	nand g1047(n_619, n_892, sub_29_29_n_66);
	nand g1048(n_970, n_875, n_881);
	nand g1049(n_620, n_1098, n_1099);
	nand g1050(n_971, n_882, add_24_29_n_1115);
	nand g1051(n_972, n_1112, n_971);
	nand g1056(n_977, sub_29_29_n_54, n_1101);
	nor g1059(n_980, n_913, n_1106);
	not g1060(n_981, n_980);
	nor g1061(n_982, n_912, n_1106);
	not g1062(n_983, n_982);
	nand g1063(n_984, sub_29_29_n_59, n_981);
	nand g1064(n_985, n_892, n_983);
	not g901(n_869, op[0]);
	nor g1029(n_1095, op[1], n_869);
	not g1030(n_960, n_1095);
	not g895(n_863, a[6]);
	nor g934(n_1096, n_863, b[6]);
	not g935(n_1097, n_1096);
	nand g969(n_300, n_863, b[6]);
	not g970(n_917, n_300);
	not g893(n_861, a[5]);
	nor g930(gt_39_12_n_52, n_861, b[5]);
	nand g960(n_298, n_861, b[5]);
	nor g282(n_416, gt_39_12_n_52, n_298);
	not g987(n_930, n_416);
	not g891(n_859, a[4]);
	nor g932(n_308, n_859, b[4]);
	nor g283(n_415, gt_39_12_n_52, n_308);
	not g988(n_931, n_415);
	nand g989(sub_29_29_n_59, n_930, n_931);
	nor g990(n_827, n_917, sub_29_29_n_59);
	not g991(n_932, n_827);
	not g961(n_911, n_298);
	nand g962(sub_29_29_n_66, n_859, b[4]);
	not g963(n_912, sub_29_29_n_66);
	nor g964(sub_29_29_n_63, n_911, n_912);
	not g889(n_857, a[3]);
	nor g940(gt_39_12_n_46, n_857, b[3]);
	not g941(n_1098, gt_39_12_n_46);
	nand g943(n_1099, n_857, b[3]);
	not g944(n_898, n_1099);
	not g899(n_867, a[2]);
	nor g945(n_806, n_867, b[2]);
	not g946(n_1101, n_806);
	nor g999(n_938, n_898, n_1101);
	not g1000(n_939, n_938);
	not g897(n_865, a[1]);
	nor g947(n_1102, n_865, b[1]);
	not g948(n_900, n_1102);
	nand g950(sub_29_29_n_1103, n_865, b[1]);
	not g951(n_902, sub_29_29_n_1103);
	not g902(n_870, a[0]);
	nand g979(sub_29_29_n_37, n_870, b[0]);
	not g980(n_924, sub_29_29_n_37);
	nor g981(n_925, n_902, n_924);
	not g982(n_926, n_925);
	nand g983(sub_29_29_n_320, n_900, n_926);
	nand g939(n_1104, n_867, b[2]);
	not g984(n_927, sub_29_29_n_54);
	nand g1001(n_940, n_927, n_1099);
	nand g1002(sub_29_29_n_1105, n_1098, n_939, n_940);
	not g1003(n_1106, sub_29_29_n_1105);
	nor g1010(n_945, sub_29_29_n_69, n_1106);
	not g1011(n_946, n_945);
	nand g1012(sub_29_29_n_32, n_1097, n_932, n_946);
	nor g1031(n_961, n_960, sub_29_29_n_32);
	not g1032(n_962, n_961);
	nor g108(n_1111, op[0], op[1]);
	not g986(n_929, n_1111);
	not g890(n_858, b[4]);
	nor g917(n_31, n_859, n_858);
	not g918(n_883, n_31);
	nor g919(n_884, add_24_29_n_39, n_883);
	not g892(n_860, b[5]);
	nor g920(n_35, n_861, n_860);
	not g922(n_886, add_24_29_n_55);
	not g898(n_866, b[2]);
	nor g911(n_23, n_867, n_866);
	not g912(n_1112, n_23);
	nor g913(n_880, add_24_29_n_33, n_1112);
	not g888(n_856, b[3]);
	nor g914(n_1113, n_857, n_856);
	not g896(n_864, b[1]);
	nor g923(n_19, n_865, n_864);
	not g924(n_887, n_19);
	not g925(n_888, add_24_29_n_27);
	not g903(n_871, b[0]);
	nor g926(n_1114, n_870, n_871);
	nand g927(n_889, n_888, n_1114);
	nand g928(add_24_29_n_1115, n_887, n_889);
	not g1013(n_947, add_24_29_n_57);
	nor g1052(n_973, n_886, n_947);
	not g1053(n_974, n_973);
	nand g1057(n_978, add_24_29_n_51, n_974);
	not g910(n_878, add_24_29_n_50);
	not g894(n_862, b[6]);
	nor g1014(n_39, n_863, n_862);
	not g1015(n_948, n_39);
	nand g1040(n_967, n_878, n_948);
	not g905(n_873, n_37);
	not g908(n_876, add_24_29_n_43);
	nand g1046(n_969, n_876, n_883);
	not g929(n_890, add_24_29_n_53);
	nand g1016(n_949, n_878, add_24_29_n_55);
	nor g1017(n_950, n_947, n_949);
	not g1018(n_951, n_950);
	nand g1019(n_41, n_890, n_948, n_951);
	nor g307(n_436, n_29, n_41);
	not g1021(n_953, n_436);
	nor g1054(n_975, add_24_29_n_43, n_947);
	not g1055(n_976, n_975);
	nand g1058(n_979, n_883, n_976);
	not g909(n_877, add_24_29_n_39);
	not g921(n_885, n_35);
	nand g1042(n_968, n_877, n_885);
	nor g308(n_435, n_33, n_41);
	not g1022(n_954, n_435);
	nand g1023(n_437, n_953, n_954);
	nor g1024(n_955, n_873, n_437);
	not g1025(n_956, n_955);
	not g1020(n_952, n_41);
	nor g1026(n_957, n_952, n_437);
	not g1027(n_958, n_957);
	nand g1028(n_959, n_956, n_958);
	nand g498(gt_25_24_n_35, n_959, n_41);
	nor g1033(n_963, n_929, gt_25_24_n_35);
	not g1034(n_964, n_963);
	nand g1035(sub_wire2, n_962, n_964);
	not g900(n_1123, op[1]);
	nand g1065(n_986, overflow, n_1123);
	not g906(n_874, overflow);
	nor g1066(n_987, n_874, n_929);
	nor g1067(n_988, n_874, n_960);
	and g1068(sub_wire3, overflow, n_135);
	and g1069(sub_wire4, overflow, n_136);
	and g1070(sub_wire5, overflow, n_132);
	and g1071(sub_wire6, overflow, n_133);
	and g1072(sub_wire7, overflow, n_131);
	and g1073(sub_wire8, overflow, n_130);
	and g1074(sub_wire9, overflow, n_129);
	and _ECO_0(w_eco0, a[7], !b[7], !op[1]);
	and _ECO_1(w_eco1, !a[7], b[7], !op[1]);
	or _ECO_2(w_eco2, w_eco0, w_eco1);
	xor _ECO_out0(y[7], sub_wire0, w_eco2);
	and _ECO_3(w_eco3, !b[4], !b[5], !b[6], a[7]);
	and _ECO_4(w_eco4, !b[4], a[5], !b[6], a[7]);
	and _ECO_5(w_eco5, a[4], !b[5], !b[6], a[7]);
	and _ECO_6(w_eco6, !b[4], !b[5], a[6], a[7]);
	and _ECO_7(w_eco7, !b[4], !b[5], !b[6], !b[7]);
	and _ECO_8(w_eco8, a[4], a[5], !b[6], a[7]);
	and _ECO_9(w_eco9, !b[4], a[5], a[6], a[7]);
	and _ECO_10(w_eco10, !b[4], a[5], !b[6], !b[7]);
	and _ECO_11(w_eco11, a[3], !b[3], b[1], !a[0], b[0]);
	and _ECO_12(w_eco12, a[3], !b[3], !a[1], b[1]);
	and _ECO_13(w_eco13, a[3], !b[3], !a[2], b[2]);
	and _ECO_14(w_eco14, a[4], !b[5], a[6], a[7]);
	and _ECO_15(w_eco15, a[4], !b[5], !b[6], !b[7]);
	and _ECO_16(w_eco16, !b[4], !b[5], a[6], !b[7]);
	and _ECO_17(w_eco17, a[4], a[5], a[6], a[7]);
	and _ECO_18(w_eco18, a[4], a[5], !b[6], !b[7]);
	and _ECO_19(w_eco19, !b[4], a[5], a[6], !b[7]);
	and _ECO_20(w_eco20, a[3], b[1], a[2], !b[2], !a[0], b[0]);
	and _ECO_21(w_eco21, a[3], !a[1], b[1], a[2], !b[2]);
	and _ECO_22(w_eco22, a[3], !b[3], !a[1], !a[0], b[0]);
	and _ECO_23(w_eco23, !b[3], b[1], a[2], !b[2], !a[0], b[0]);
	and _ECO_24(w_eco24, !b[3], !a[1], b[1], a[2], !b[2]);
	and _ECO_25(w_eco25, a[4], !b[5], a[6], !b[7]);
	and _ECO_26(w_eco26, a[4], a[5], a[6], !b[7]);
	and _ECO_27(w_eco27, a[3], !a[1], a[2], !b[2], !a[0], b[0]);
	and _ECO_28(w_eco28, !b[3], !a[1], a[2], !b[2], !a[0], b[0]);
	or _ECO_29(w_eco29, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28);
	xor _ECO_out1(less, sub_wire1, w_eco29);
	and _ECO_30(w_eco30, a[4], b[4], a[5], b[5], a[6], b[6], op[0], !op[1]);
	and _ECO_31(w_eco31, a[4], b[4], a[5], b[5], !a[6], !b[6], op[0], !op[1]);
	and _ECO_32(w_eco32, !a[4], !b[4], a[5], b[5], a[6], b[6], op[0], !op[1]);
	and _ECO_33(w_eco33, !a[4], !b[4], a[5], b[5], !a[6], !b[6], op[0], !op[1]);
	and _ECO_34(w_eco34, a[4], b[4], !a[5], !b[5], a[6], b[6], op[0], !op[1]);
	and _ECO_35(w_eco35, a[4], b[4], !a[5], !b[5], !a[6], !b[6], op[0], !op[1]);
	and _ECO_36(w_eco36, !a[4], !b[4], !a[5], !b[5], a[6], b[6], op[0], !op[1]);
	and _ECO_37(w_eco37, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], op[0], !op[1]);
	and _ECO_38(w_eco38, !a[4], !b[4], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_39(w_eco39, !a[4], !b[4], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_40(w_eco40, !a[4], !b[4], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_41(w_eco41, !a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_42(w_eco42, !a[3], a[4], b[4], a[5], b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_43(w_eco43, b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_44(w_eco44, b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_45(w_eco45, !a[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_46(w_eco46, !a[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_47(w_eco47, !a[4], !b[4], a[6], b[6], a[7], !b[7], !op[1]);
	and _ECO_48(w_eco48, !a[4], !b[4], a[5], b[5], b[6], a[7], !b[7], !op[1]);
	and _ECO_49(w_eco49, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_50(w_eco50, !a[4], !b[4], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_51(w_eco51, !a[5], !b[5], a[6], b[6], a[7], !b[7], !op[1]);
	and _ECO_52(w_eco52, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_53(w_eco53, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_54(w_eco54, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], op[0], !op[1]);
	and _ECO_55(w_eco55, b[3], a[4], b[4], a[5], b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_56(w_eco56, !a[3], !b[3], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_57(w_eco57, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], op[0], !op[1]);
	and _ECO_58(w_eco58, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_59(w_eco59, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_60(w_eco60, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], op[0], !op[1]);
	and _ECO_61(w_eco61, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_62(w_eco62, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], op[0], !op[1]);
	and _ECO_63(w_eco63, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], op[0], !op[1]);
	and _ECO_64(w_eco64, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_65(w_eco65, !a[3], !b[3], a[5], b[5], b[6], a[7], !b[7], !op[1]);
	and _ECO_66(w_eco66, !a[3], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_67(w_eco67, !a[3], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_68(w_eco68, !a[3], !b[3], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_69(w_eco69, !a[3], !b[3], a[4], b[4], b[5], b[6], a[7], !b[7], !op[1]);
	and _ECO_70(w_eco70, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_71(w_eco71, !a[3], !b[3], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_72(w_eco72, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_73(w_eco73, b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_74(w_eco74, a[4], b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_75(w_eco75, !a[3], !b[3], a[4], b[4], a[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_76(w_eco76, !b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_77(w_eco77, !a[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_78(w_eco78, !a[3], b[3], a[7], !b[7], op[0], !op[1]);
	and _ECO_79(w_eco79, !a[3], b[3], !a[7], b[7], op[0], !op[1]);
	and _ECO_80(w_eco80, b[3], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_81(w_eco81, b[3], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_82(w_eco82, !a[3], !b[3], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_83(w_eco83, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_84(w_eco84, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_85(w_eco85, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_86(w_eco86, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_87(w_eco87, !a[3], !b[3], a[4], b[4], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_88(w_eco88, !a[3], !b[3], a[6], b[6], a[7], !b[7], !op[1]);
	and _ECO_89(w_eco89, !a[3], !b[3], a[4], b[4], a[5], b[6], a[7], !b[7], !op[1]);
	and _ECO_90(w_eco90, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_91(w_eco91, a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_92(w_eco92, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_93(w_eco93, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_94(w_eco94, b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_95(w_eco95, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_96(w_eco96, a[4], b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_97(w_eco97, a[4], b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_98(w_eco98, a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_99(w_eco99, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_100(w_eco100, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_101(w_eco101, !b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_102(w_eco102, !a[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_103(w_eco103, !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_104(w_eco104, !b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_105(w_eco105, !b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_106(w_eco106, !a[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_107(w_eco107, !a[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_108(w_eco108, !a[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_109(w_eco109, !b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_110(w_eco110, !a[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_111(w_eco111, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_112(w_eco112, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_113(w_eco113, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_114(w_eco114, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_115(w_eco115, !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_116(w_eco116, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_117(w_eco117, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_118(w_eco118, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_119(w_eco119, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[1]);
	and _ECO_120(w_eco120, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_121(w_eco121, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_122(w_eco122, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_123(w_eco123, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_124(w_eco124, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_125(w_eco125, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_126(w_eco126, !b[3], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_127(w_eco127, !a[3], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_128(w_eco128, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_129(w_eco129, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_130(w_eco130, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_131(w_eco131, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_132(w_eco132, a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_133(w_eco133, a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_134(w_eco134, a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_135(w_eco135, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_136(w_eco136, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_137(w_eco137, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_138(w_eco138, !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_139(w_eco139, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_140(w_eco140, b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[0], op[0], !op[1]);
	and _ECO_141(w_eco141, b[3], a[4], b[4], a[5], b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_142(w_eco142, a[4], b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_143(w_eco143, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_144(w_eco144, !a[3], a[4], b[4], a[5], b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_145(w_eco145, a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_146(w_eco146, a[4], b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_147(w_eco147, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_148(w_eco148, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_149(w_eco149, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_150(w_eco150, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_151(w_eco151, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_152(w_eco152, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_153(w_eco153, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_154(w_eco154, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_155(w_eco155, a[3], !b[3], !a[4], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_156(w_eco156, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_157(w_eco157, a[3], !b[3], !a[4], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_158(w_eco158, !b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_159(w_eco159, !b[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_160(w_eco160, !b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_161(w_eco161, !a[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_162(w_eco162, !a[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_163(w_eco163, !a[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_164(w_eco164, !b[3], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_165(w_eco165, !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_166(w_eco166, !b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_167(w_eco167, !a[3], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_168(w_eco168, !a[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_169(w_eco169, !a[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_170(w_eco170, b[3], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_171(w_eco171, b[3], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_172(w_eco172, !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_173(w_eco173, !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_174(w_eco174, !b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_175(w_eco175, !a[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_176(w_eco176, !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_177(w_eco177, !b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_178(w_eco178, !b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_179(w_eco179, !a[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_180(w_eco180, !a[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_181(w_eco181, !a[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_182(w_eco182, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[0], op[0], !op[1]);
	and _ECO_183(w_eco183, b[3], !a[4], !b[4], a[5], b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_184(w_eco184, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_185(w_eco185, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_186(w_eco186, !a[3], !a[4], !b[4], a[5], b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_187(w_eco187, !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_188(w_eco188, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_189(w_eco189, a[3], !b[3], b[4], !a[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_190(w_eco190, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_191(w_eco191, a[3], !b[3], b[4], !a[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_192(w_eco192, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_193(w_eco193, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_194(w_eco194, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_195(w_eco195, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_196(w_eco196, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_197(w_eco197, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_198(w_eco198, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_199(w_eco199, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_200(w_eco200, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_201(w_eco201, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_202(w_eco202, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_203(w_eco203, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_204(w_eco204, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_205(w_eco205, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_206(w_eco206, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_207(w_eco207, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_208(w_eco208, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_209(w_eco209, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_210(w_eco210, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_211(w_eco211, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_212(w_eco212, !b[3], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_213(w_eco213, !a[3], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_214(w_eco214, !b[3], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_215(w_eco215, !b[3], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_216(w_eco216, !b[3], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_217(w_eco217, !a[3], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_218(w_eco218, !a[3], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_219(w_eco219, !a[3], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_220(w_eco220, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_221(w_eco221, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_222(w_eco222, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_223(w_eco223, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_224(w_eco224, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_225(w_eco225, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_226(w_eco226, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_227(w_eco227, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_228(w_eco228, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[0], op[0], !op[1]);
	and _ECO_229(w_eco229, b[3], a[4], b[4], !a[5], !b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_230(w_eco230, a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_231(w_eco231, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_232(w_eco232, !a[3], a[4], b[4], !a[5], !b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_233(w_eco233, a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_234(w_eco234, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_235(w_eco235, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[0], op[0], !op[1]);
	and _ECO_236(w_eco236, b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_237(w_eco237, !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_238(w_eco238, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_239(w_eco239, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], op[0], !op[1]);
	and _ECO_240(w_eco240, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_241(w_eco241, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_242(w_eco242, a[3], !b[3], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_243(w_eco243, a[3], !b[3], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_244(w_eco244, a[3], !b[3], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_245(w_eco245, a[4], b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_246(w_eco246, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_247(w_eco247, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_248(w_eco248, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_249(w_eco249, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_250(w_eco250, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_251(w_eco251, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_252(w_eco252, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_253(w_eco253, !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_254(w_eco254, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_255(w_eco255, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_256(w_eco256, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_257(w_eco257, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_258(w_eco258, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_259(w_eco259, a[3], !a[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_260(w_eco260, a[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_261(w_eco261, a[3], !b[3], !a[4], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_262(w_eco262, !b[3], !a[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_263(w_eco263, !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_264(w_eco264, !b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_265(w_eco265, !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_266(w_eco266, !b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_267(w_eco267, !b[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_268(w_eco268, !a[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_269(w_eco269, !a[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_270(w_eco270, !a[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_271(w_eco271, !a[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_272(w_eco272, !b[3], a[5], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_273(w_eco273, !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_274(w_eco274, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_275(w_eco275, !a[3], a[5], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_276(w_eco276, !a[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_277(w_eco277, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_278(w_eco278, b[3], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_279(w_eco279, b[3], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_280(w_eco280, b[3], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_281(w_eco281, b[3], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_282(w_eco282, !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_283(w_eco283, !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_284(w_eco284, a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_285(w_eco285, a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_286(w_eco286, !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_287(w_eco287, !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_288(w_eco288, !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_289(w_eco289, !b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_290(w_eco290, !b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_291(w_eco291, !a[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_292(w_eco292, !a[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_293(w_eco293, !a[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_294(w_eco294, !b[3], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_295(w_eco295, !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_296(w_eco296, !b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_297(w_eco297, !a[3], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_298(w_eco298, !a[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_299(w_eco299, !a[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_300(w_eco300, a[3], !b[3], !a[4], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_301(w_eco301, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_302(w_eco302, a[3], !b[3], !a[4], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_303(w_eco303, a[4], !b[4], a[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_304(w_eco304, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_305(w_eco305, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_306(w_eco306, a[3], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_307(w_eco307, a[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_308(w_eco308, a[3], !b[3], b[4], !a[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_309(w_eco309, !b[3], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_310(w_eco310, !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_311(w_eco311, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[1]);
	and _ECO_312(w_eco312, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_313(w_eco313, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_314(w_eco314, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_315(w_eco315, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_316(w_eco316, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_317(w_eco317, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_318(w_eco318, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_319(w_eco319, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_320(w_eco320, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[1]);
	and _ECO_321(w_eco321, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_322(w_eco322, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_323(w_eco323, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_324(w_eco324, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_325(w_eco325, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_326(w_eco326, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_327(w_eco327, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_328(w_eco328, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_329(w_eco329, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_330(w_eco330, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_331(w_eco331, !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_332(w_eco332, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_333(w_eco333, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_334(w_eco334, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_335(w_eco335, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_336(w_eco336, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_337(w_eco337, a[3], !b[3], b[4], !a[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_338(w_eco338, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_339(w_eco339, a[3], !b[3], b[4], !a[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_340(w_eco340, !b[3], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_341(w_eco341, !b[3], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_342(w_eco342, !b[3], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_343(w_eco343, !a[3], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_344(w_eco344, !a[3], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_345(w_eco345, !a[3], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_346(w_eco346, !b[3], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_347(w_eco347, !b[3], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_348(w_eco348, !b[3], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_349(w_eco349, !a[3], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_350(w_eco350, !a[3], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_351(w_eco351, !a[3], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_352(w_eco352, a[3], !b[3], !a[5], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_353(w_eco353, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_354(w_eco354, a[3], !b[3], !a[5], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_355(w_eco355, a[3], !b[3], !a[5], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_356(w_eco356, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_357(w_eco357, a[3], !b[3], !a[5], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_358(w_eco358, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_359(w_eco359, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_360(w_eco360, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_361(w_eco361, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_362(w_eco362, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_363(w_eco363, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_364(w_eco364, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_365(w_eco365, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_366(w_eco366, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_367(w_eco367, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_368(w_eco368, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_369(w_eco369, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_370(w_eco370, a[5], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_371(w_eco371, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_372(w_eco372, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_373(w_eco373, a[4], !b[4], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_374(w_eco374, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_375(w_eco375, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_376(w_eco376, a[3], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_377(w_eco377, a[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_378(w_eco378, a[3], !b[3], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_379(w_eco379, !b[3], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_380(w_eco380, !b[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_381(w_eco381, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_382(w_eco382, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_383(w_eco383, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_384(w_eco384, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_385(w_eco385, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_386(w_eco386, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_387(w_eco387, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_388(w_eco388, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_389(w_eco389, !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_390(w_eco390, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_391(w_eco391, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_392(w_eco392, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_393(w_eco393, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_394(w_eco394, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_395(w_eco395, a[3], !a[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_396(w_eco396, !b[3], !a[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_397(w_eco397, !b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_398(w_eco398, !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_399(w_eco399, !a[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_400(w_eco400, !a[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_401(w_eco401, !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_402(w_eco402, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_403(w_eco403, !a[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_404(w_eco404, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_405(w_eco405, b[3], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_406(w_eco406, b[3], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_407(w_eco407, b[3], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_408(w_eco408, b[3], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_409(w_eco409, a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_410(w_eco410, a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_411(w_eco411, a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_412(w_eco412, a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_413(w_eco413, !a[3], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_414(w_eco414, !a[3], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_415(w_eco415, !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_416(w_eco416, !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_417(w_eco417, a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_418(w_eco418, a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_419(w_eco419, !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_420(w_eco420, !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_421(w_eco421, !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_422(w_eco422, !b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_423(w_eco423, !a[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_424(w_eco424, !a[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_425(w_eco425, !a[3], b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_426(w_eco426, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_427(w_eco427, !b[3], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_428(w_eco428, !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_429(w_eco429, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_430(w_eco430, !a[3], a[5], b[5], a[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_431(w_eco431, !a[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_432(w_eco432, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_433(w_eco433, a[3], !a[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_434(w_eco434, a[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_435(w_eco435, a[3], !b[3], !a[4], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_436(w_eco436, !b[3], !a[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_437(w_eco437, !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_438(w_eco438, a[3], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_439(w_eco439, !b[3], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_440(w_eco440, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_441(w_eco441, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_442(w_eco442, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_443(w_eco443, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_444(w_eco444, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_445(w_eco445, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_446(w_eco446, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_447(w_eco447, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_448(w_eco448, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_449(w_eco449, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_450(w_eco450, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_451(w_eco451, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_452(w_eco452, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_453(w_eco453, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_454(w_eco454, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_455(w_eco455, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_456(w_eco456, !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_457(w_eco457, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_458(w_eco458, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_459(w_eco459, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_460(w_eco460, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_461(w_eco461, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_462(w_eco462, a[3], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_463(w_eco463, a[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_464(w_eco464, a[3], !b[3], b[4], !a[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_465(w_eco465, !b[3], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_466(w_eco466, !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_467(w_eco467, !b[3], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_468(w_eco468, !b[3], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_469(w_eco469, !b[3], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_470(w_eco470, !b[3], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_471(w_eco471, !a[3], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_472(w_eco472, !a[3], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_473(w_eco473, !a[3], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_474(w_eco474, !a[3], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_475(w_eco475, !b[3], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_476(w_eco476, !b[3], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_477(w_eco477, !b[3], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_478(w_eco478, !a[3], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_479(w_eco479, !a[3], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_480(w_eco480, !a[3], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_481(w_eco481, a[3], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_482(w_eco482, a[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_483(w_eco483, a[3], !b[3], !a[5], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_484(w_eco484, !b[3], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_485(w_eco485, !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_486(w_eco486, a[3], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_487(w_eco487, a[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_488(w_eco488, a[3], !b[3], !a[5], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_489(w_eco489, !b[3], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_490(w_eco490, !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_491(w_eco491, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_492(w_eco492, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_493(w_eco493, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_494(w_eco494, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_495(w_eco495, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_496(w_eco496, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_497(w_eco497, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_498(w_eco498, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_499(w_eco499, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_500(w_eco500, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_501(w_eco501, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_502(w_eco502, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_503(w_eco503, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_504(w_eco504, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_505(w_eco505, a[3], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_506(w_eco506, !b[3], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_507(w_eco507, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_508(w_eco508, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_509(w_eco509, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_510(w_eco510, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_511(w_eco511, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_512(w_eco512, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_513(w_eco513, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_514(w_eco514, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_515(w_eco515, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_516(w_eco516, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_517(w_eco517, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_518(w_eco518, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_519(w_eco519, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_520(w_eco520, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_521(w_eco521, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_522(w_eco522, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_523(w_eco523, a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_524(w_eco524, a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_525(w_eco525, a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_526(w_eco526, a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_527(w_eco527, !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_528(w_eco528, !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_529(w_eco529, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_530(w_eco530, !a[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_531(w_eco531, !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_532(w_eco532, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_533(w_eco533, !a[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_534(w_eco534, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_535(w_eco535, a[3], !a[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_536(w_eco536, !b[3], !a[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_537(w_eco537, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_538(w_eco538, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_539(w_eco539, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_540(w_eco540, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_541(w_eco541, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_542(w_eco542, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_543(w_eco543, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_544(w_eco544, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_545(w_eco545, a[3], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_546(w_eco546, !b[3], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_547(w_eco547, !b[3], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_548(w_eco548, !b[3], a[6], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_549(w_eco549, !a[3], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_550(w_eco550, !a[3], a[6], b[6], !a[1], !b[1], !b[2], a[7], !b[7], !op[1]);
	and _ECO_551(w_eco551, !b[3], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_552(w_eco552, !b[3], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_553(w_eco553, !a[3], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_554(w_eco554, !a[3], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_555(w_eco555, a[3], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_556(w_eco556, !b[3], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_557(w_eco557, a[3], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_558(w_eco558, !b[3], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	or _ECO_559(w_eco559, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558);
	xor _ECO_out2(overflow, sub_wire2, w_eco559);
	and _ECO_560(w_eco560, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_561(w_eco561, !a[3], a[4], b[4], a[5], b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_562(w_eco562, !a[4], !b[4], a[5], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_563(w_eco563, !a[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_564(w_eco564, !a[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_565(w_eco565, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_566(w_eco566, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !b[6], op[0], !op[1]);
	and _ECO_567(w_eco567, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_568(w_eco568, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], op[0], !op[1]);
	and _ECO_569(w_eco569, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_570(w_eco570, !a[5], b[5], a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_571(w_eco571, !a[5], b[5], a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_572(w_eco572, !a[5], b[5], !a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_573(w_eco573, !a[5], b[5], !a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_574(w_eco574, !a[3], !b[4], a[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_575(w_eco575, !a[3], !b[4], a[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_576(w_eco576, !a[3], !b[4], a[5], a[6], !b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_577(w_eco577, !a[3], !b[4], a[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_578(w_eco578, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], op[0], !op[1]);
	and _ECO_579(w_eco579, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_580(w_eco580, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], op[0], !op[1]);
	and _ECO_581(w_eco581, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !a[2], op[0], !op[1]);
	and _ECO_582(w_eco582, !a[3], !b[3], a[4], b[4], a[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_583(w_eco583, !a[3], a[4], a[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_584(w_eco584, !a[3], a[4], a[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_585(w_eco585, !a[4], b[4], b[5], a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_586(w_eco586, !a[4], b[4], b[5], a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_587(w_eco587, !a[3], !b[3], a[5], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_588(w_eco588, !a[4], b[4], b[5], !a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_589(w_eco589, !a[4], b[4], b[5], !a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_590(w_eco590, !a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_591(w_eco591, !a[3], a[4], a[5], a[6], !b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_592(w_eco592, !a[3], a[4], a[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_593(w_eco593, a[5], !b[5], !a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_594(w_eco594, a[5], !b[5], !a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_595(w_eco595, a[5], !b[5], a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_596(w_eco596, !a[3], a[5], !b[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_597(w_eco597, !a[3], b[3], !b[4], a[5], a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_598(w_eco598, b[3], !b[4], a[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_599(w_eco599, !a[3], a[4], !b[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_600(w_eco600, !a[3], a[4], !b[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_601(w_eco601, !a[4], b[4], !a[5], a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_602(w_eco602, !a[4], b[4], !a[5], a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_603(w_eco603, !a[4], b[4], !a[5], !a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_604(w_eco604, !a[4], b[4], !a[5], !a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_605(w_eco605, !a[3], a[4], !b[5], a[6], !b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_606(w_eco606, !a[3], a[4], !b[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_607(w_eco607, !a[3], !b[4], !b[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_608(w_eco608, !a[3], !b[4], !b[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_609(w_eco609, !a[3], !b[3], a[4], b[4], a[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_610(w_eco610, !a[3], b[3], a[4], a[5], !a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_611(w_eco611, !a[3], b[3], a[4], a[5], !a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_612(w_eco612, b[3], a[4], a[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_613(w_eco613, b[3], a[4], a[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_614(w_eco614, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_615(w_eco615, a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_616(w_eco616, !a[3], !b[3], a[5], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_617(w_eco617, !a[3], b[3], a[4], a[5], a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_618(w_eco618, b[3], a[4], a[5], a[6], !b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_619(w_eco619, !a[3], b[3], !b[4], a[5], !a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_620(w_eco620, !a[3], b[3], !b[4], a[5], !a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_621(w_eco621, b[3], !b[4], a[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_622(w_eco622, b[3], !b[4], a[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_623(w_eco623, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_624(w_eco624, !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_625(w_eco625, !a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_626(w_eco626, !a[3], b[3], a[4], a[5], a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_627(w_eco627, b[3], a[4], a[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_628(w_eco628, !a[3], b[3], a[5], !b[5], a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_629(w_eco629, b[3], a[5], !b[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_630(w_eco630, !a[3], b[3], a[4], !b[5], !a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_631(w_eco631, !a[3], b[3], a[4], !b[5], !a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_632(w_eco632, b[3], a[4], !b[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_633(w_eco633, b[3], a[4], !b[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_634(w_eco634, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_635(w_eco635, a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_636(w_eco636, !a[3], b[3], a[4], !b[5], a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_637(w_eco637, !a[3], b[3], a[4], !b[5], a[6], !b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_638(w_eco638, b[3], a[4], !b[5], a[6], !b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_639(w_eco639, b[3], a[4], !b[5], a[6], !b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_640(w_eco640, !a[3], b[3], !b[4], !b[5], !a[6], b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_641(w_eco641, !a[3], b[3], !b[4], !b[5], !a[6], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_642(w_eco642, b[3], !b[4], !b[5], !a[6], b[6], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_643(w_eco643, b[3], !b[4], !b[5], !a[6], b[6], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_644(w_eco644, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[0], op[0], !op[1]);
	and _ECO_645(w_eco645, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_646(w_eco646, a[3], !b[3], b[4], b[5], a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_647(w_eco647, a[3], !b[3], b[4], b[5], a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_648(w_eco648, a[3], !b[3], b[4], b[5], a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_649(w_eco649, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_650(w_eco650, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_651(w_eco651, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_652(w_eco652, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_653(w_eco653, a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_654(w_eco654, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_655(w_eco655, a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_656(w_eco656, a[3], !b[3], b[4], b[5], !a[6], !b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_657(w_eco657, a[3], !b[3], b[4], b[5], !a[6], !b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_658(w_eco658, a[3], !b[3], b[4], b[5], !a[6], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_659(w_eco659, !b[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_660(w_eco660, !a[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_661(w_eco661, a[3], !b[3], a[4], !b[4], a[5], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_662(w_eco662, a[3], !b[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_663(w_eco663, a[3], !b[3], a[4], !b[4], a[5], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_664(w_eco664, a[3], !b[3], !a[4], b[5], a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_665(w_eco665, a[3], !b[3], !a[4], b[5], a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_666(w_eco666, a[3], !b[3], !a[4], b[5], a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_667(w_eco667, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_668(w_eco668, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_669(w_eco669, !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_670(w_eco670, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_671(w_eco671, !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_672(w_eco672, a[3], !b[3], !a[4], b[5], !a[6], !b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_673(w_eco673, a[3], !b[3], !a[4], b[5], !a[6], !b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_674(w_eco674, a[3], !b[3], !a[4], b[5], !a[6], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_675(w_eco675, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_676(w_eco676, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_677(w_eco677, a[3], !b[3], b[4], !a[5], a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_678(w_eco678, a[3], !b[3], b[4], !a[5], a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_679(w_eco679, a[3], !b[3], b[4], !a[5], a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_680(w_eco680, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_681(w_eco681, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_682(w_eco682, a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_683(w_eco683, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_684(w_eco684, a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_685(w_eco685, a[3], !b[3], b[4], !a[5], !a[6], !b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_686(w_eco686, a[3], !b[3], b[4], !a[5], !a[6], !b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_687(w_eco687, a[3], !b[3], b[4], !a[5], !a[6], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_688(w_eco688, a[3], !b[3], a[4], !b[4], !b[5], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_689(w_eco689, a[3], !b[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_690(w_eco690, a[3], !b[3], a[4], !b[4], !b[5], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_691(w_eco691, a[3], !b[3], !a[4], !a[5], a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_692(w_eco692, a[3], !b[3], !a[4], !a[5], a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_693(w_eco693, a[3], !b[3], !a[4], !a[5], a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_694(w_eco694, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[0], op[0], !op[1]);
	and _ECO_695(w_eco695, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[0], op[0], !op[1]);
	and _ECO_696(w_eco696, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_697(w_eco697, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_698(w_eco698, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_699(w_eco699, a[3], !b[3], !a[4], !a[5], !a[6], !b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_700(w_eco700, a[3], !b[3], !a[4], !a[5], !a[6], !b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_701(w_eco701, a[3], !b[3], !a[4], !a[5], !a[6], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_702(w_eco702, a[3], b[4], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_703(w_eco703, a[3], b[4], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_704(w_eco704, a[3], !b[3], b[4], b[5], a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_705(w_eco705, !b[3], b[4], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_706(w_eco706, !b[3], b[4], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_707(w_eco707, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_708(w_eco708, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_709(w_eco709, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_710(w_eco710, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_711(w_eco711, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_712(w_eco712, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_713(w_eco713, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_714(w_eco714, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_715(w_eco715, b[3], a[4], a[5], !a[6], b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_716(w_eco716, b[3], a[4], a[5], !a[6], b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_717(w_eco717, a[4], a[5], !a[6], b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_718(w_eco718, a[4], a[5], !a[6], b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_719(w_eco719, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], a[1], a[0], op[0], !op[1]);
	and _ECO_720(w_eco720, b[3], a[4], b[4], a[5], b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_721(w_eco721, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_722(w_eco722, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_723(w_eco723, !a[3], a[4], b[4], a[5], b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_724(w_eco724, a[4], b[4], a[5], b[5], a[6], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_725(w_eco725, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_726(w_eco726, a[3], b[4], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_727(w_eco727, a[3], b[4], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_728(w_eco728, a[3], !b[3], b[4], b[5], !a[6], !b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_729(w_eco729, !b[3], b[4], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_730(w_eco730, !b[3], b[4], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_731(w_eco731, !b[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_732(w_eco732, !a[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_733(w_eco733, !b[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_734(w_eco734, !b[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_735(w_eco735, !b[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_736(w_eco736, !a[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_737(w_eco737, !a[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_738(w_eco738, !a[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_739(w_eco739, a[3], a[4], !b[4], a[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_740(w_eco740, a[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_741(w_eco741, a[3], !b[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_742(w_eco742, !b[3], a[4], !b[4], a[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_743(w_eco743, !b[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_744(w_eco744, b[3], a[4], a[5], a[6], !b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_745(w_eco745, b[3], a[4], a[5], a[6], !b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_746(w_eco746, a[4], a[5], a[6], !b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_747(w_eco747, a[4], a[5], a[6], !b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_748(w_eco748, a[3], !a[4], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_749(w_eco749, a[3], !a[4], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_750(w_eco750, a[3], !b[3], !a[4], b[5], a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_751(w_eco751, !b[3], !a[4], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_752(w_eco752, !b[3], !a[4], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_753(w_eco753, b[3], !b[4], a[5], !a[6], b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_754(w_eco754, b[3], !b[4], a[5], !a[6], b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_755(w_eco755, !b[4], a[5], !a[6], b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_756(w_eco756, !b[4], a[5], !a[6], b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_757(w_eco757, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], a[0], op[0], !op[1]);
	and _ECO_758(w_eco758, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_759(w_eco759, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_760(w_eco760, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_761(w_eco761, !a[3], !a[4], !b[4], a[5], b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_762(w_eco762, !a[4], !b[4], a[5], b[5], a[6], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_763(w_eco763, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_764(w_eco764, a[3], !a[4], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_765(w_eco765, a[3], !a[4], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_766(w_eco766, a[3], !b[3], !a[4], b[5], !a[6], !b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_767(w_eco767, !b[3], !a[4], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_768(w_eco768, !b[3], !a[4], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_769(w_eco769, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_770(w_eco770, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_771(w_eco771, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_772(w_eco772, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[1]);
	and _ECO_773(w_eco773, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_774(w_eco774, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_775(w_eco775, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_776(w_eco776, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_777(w_eco777, b[3], a[5], !b[5], a[6], !b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_778(w_eco778, a[5], !b[5], a[6], !b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_779(w_eco779, a[3], b[4], !a[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_780(w_eco780, a[3], b[4], !a[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_781(w_eco781, a[3], !b[3], b[4], !a[5], a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_782(w_eco782, !b[3], b[4], !a[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_783(w_eco783, !b[3], b[4], !a[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_784(w_eco784, b[3], a[4], !b[5], !a[6], b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_785(w_eco785, b[3], a[4], !b[5], !a[6], b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_786(w_eco786, a[4], !b[5], !a[6], b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_787(w_eco787, a[4], !b[5], !a[6], b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_788(w_eco788, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], a[0], op[0], !op[1]);
	and _ECO_789(w_eco789, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_790(w_eco790, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_791(w_eco791, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_792(w_eco792, !a[3], a[4], b[4], !a[5], !b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_793(w_eco793, a[4], b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_794(w_eco794, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_795(w_eco795, a[3], b[4], !a[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_796(w_eco796, a[3], b[4], !a[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_797(w_eco797, a[3], !b[3], b[4], !a[5], !a[6], !b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_798(w_eco798, !b[3], b[4], !a[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_799(w_eco799, !b[3], b[4], !a[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_800(w_eco800, a[3], a[4], !b[4], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_801(w_eco801, a[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_802(w_eco802, a[3], !b[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_803(w_eco803, !b[3], a[4], !b[4], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_804(w_eco804, !b[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_805(w_eco805, b[3], a[4], !b[5], a[6], !b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_806(w_eco806, b[3], a[4], !b[5], a[6], !b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_807(w_eco807, a[4], !b[5], a[6], !b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_808(w_eco808, a[4], !b[5], a[6], !b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_809(w_eco809, a[3], !a[4], !a[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_810(w_eco810, a[3], !a[4], !a[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_811(w_eco811, a[3], !b[3], !a[4], !a[5], a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_812(w_eco812, !b[3], !a[4], !a[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_813(w_eco813, !b[3], !a[4], !a[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_814(w_eco814, b[3], !b[4], !b[5], !a[6], b[6], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_815(w_eco815, b[3], !b[4], !b[5], !a[6], b[6], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_816(w_eco816, !b[4], !b[5], !a[6], b[6], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_817(w_eco817, !b[4], !b[5], !a[6], b[6], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_818(w_eco818, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], a[0], op[0], !op[1]);
	and _ECO_819(w_eco819, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_820(w_eco820, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_821(w_eco821, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_822(w_eco822, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[6], b[2], op[0], !op[1]);
	and _ECO_823(w_eco823, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_824(w_eco824, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_825(w_eco825, a[3], !a[4], !a[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_826(w_eco826, a[3], !a[4], !a[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_827(w_eco827, a[3], !b[3], !a[4], !a[5], !a[6], !b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_828(w_eco828, !b[3], !a[4], !a[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_829(w_eco829, !b[3], !a[4], !a[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_830(w_eco830, a[3], b[4], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_831(w_eco831, !b[3], b[4], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_832(w_eco832, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_833(w_eco833, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_834(w_eco834, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_835(w_eco835, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_836(w_eco836, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_837(w_eco837, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_838(w_eco838, !b[3], a[4], b[4], a[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_839(w_eco839, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_840(w_eco840, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_841(w_eco841, !a[3], a[4], b[4], a[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_842(w_eco842, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_843(w_eco843, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_844(w_eco844, b[3], a[4], a[5], !a[6], b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_845(w_eco845, b[3], a[4], a[5], !a[6], b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_846(w_eco846, b[3], a[4], a[5], !a[6], b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_847(w_eco847, b[3], a[4], a[5], !a[6], b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_848(w_eco848, a[4], a[5], !a[6], b[6], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_849(w_eco849, a[4], a[5], !a[6], b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_850(w_eco850, a[4], a[5], !a[6], b[6], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_851(w_eco851, a[4], a[5], !a[6], b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_852(w_eco852, a[4], a[5], !a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_853(w_eco853, a[4], a[5], !a[6], b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_854(w_eco854, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_855(w_eco855, a[4], b[4], a[5], b[5], a[6], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_856(w_eco856, a[3], b[4], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_857(w_eco857, !b[3], b[4], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_858(w_eco858, !b[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_859(w_eco859, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_860(w_eco860, !b[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_861(w_eco861, !a[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_862(w_eco862, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_863(w_eco863, !a[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_864(w_eco864, !b[3], a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_865(w_eco865, !b[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_866(w_eco866, !b[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_867(w_eco867, !a[3], a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_868(w_eco868, !a[3], a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_869(w_eco869, !a[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_870(w_eco870, a[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_871(w_eco871, !b[3], a[4], !b[4], a[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_872(w_eco872, b[3], a[4], a[5], a[6], !b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_873(w_eco873, b[3], a[4], a[5], a[6], !b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_874(w_eco874, b[3], a[4], a[5], a[6], !b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_875(w_eco875, b[3], a[4], a[5], a[6], !b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_876(w_eco876, a[4], !b[4], a[5], a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_877(w_eco877, a[4], a[5], a[6], !b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_878(w_eco878, a[4], a[5], a[6], !b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_879(w_eco879, a[4], a[5], a[6], !b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_880(w_eco880, a[3], !a[4], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_881(w_eco881, !b[3], !a[4], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_882(w_eco882, b[3], !b[4], a[5], !a[6], b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_883(w_eco883, b[3], !b[4], a[5], !a[6], b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_884(w_eco884, b[3], !b[4], a[5], !a[6], b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_885(w_eco885, b[3], !b[4], a[5], !a[6], b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_886(w_eco886, !b[4], a[5], !a[6], b[6], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_887(w_eco887, !b[4], a[5], !a[6], b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_888(w_eco888, !b[4], a[5], !a[6], b[6], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_889(w_eco889, !b[4], a[5], !a[6], b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_890(w_eco890, !b[4], a[5], !a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_891(w_eco891, !b[4], a[5], !a[6], b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_892(w_eco892, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_893(w_eco893, !a[4], !b[4], a[5], b[5], a[6], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_894(w_eco894, a[3], !a[4], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_895(w_eco895, !b[3], !a[4], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_896(w_eco896, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_897(w_eco897, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_898(w_eco898, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_899(w_eco899, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_900(w_eco900, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_901(w_eco901, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_902(w_eco902, !b[3], a[4], b[4], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_903(w_eco903, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_904(w_eco904, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !a[2], !b[0], !b[7], !op[1]);
	and _ECO_905(w_eco905, !a[3], a[4], b[4], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_906(w_eco906, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_907(w_eco907, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_908(w_eco908, a[3], !b[3], !a[5], b[5], a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_909(w_eco909, a[3], !b[3], !a[5], b[5], a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_910(w_eco910, a[3], !b[3], !a[5], b[5], a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_911(w_eco911, a[3], !b[3], !a[5], b[5], !a[6], !b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_912(w_eco912, a[3], !b[3], !a[5], b[5], !a[6], !b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_913(w_eco913, a[3], !b[3], !a[5], b[5], !a[6], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_914(w_eco914, a[3], !b[3], a[5], !b[5], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_915(w_eco915, a[3], !b[3], a[5], !b[5], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_916(w_eco916, a[3], !b[3], a[5], !b[5], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_917(w_eco917, b[3], a[5], !b[5], a[6], !b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_918(w_eco918, b[3], a[5], !b[5], a[6], !b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_919(w_eco919, a[5], !b[5], a[6], !b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_920(w_eco920, a[5], !b[5], a[6], !b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_921(w_eco921, a[5], !b[5], a[6], !b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_922(w_eco922, a[3], b[4], !a[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_923(w_eco923, !b[3], b[4], !a[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_924(w_eco924, b[3], a[4], !b[5], !a[6], b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_925(w_eco925, b[3], a[4], !b[5], !a[6], b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_926(w_eco926, b[3], a[4], !b[5], !a[6], b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_927(w_eco927, b[3], a[4], !b[5], !a[6], b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_928(w_eco928, a[4], !b[5], !a[6], b[6], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_929(w_eco929, a[4], !b[5], !a[6], b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_930(w_eco930, a[4], !b[5], !a[6], b[6], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_931(w_eco931, a[4], !b[5], !a[6], b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_932(w_eco932, a[4], !b[5], !a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_933(w_eco933, a[4], !b[5], !a[6], b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_934(w_eco934, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_935(w_eco935, a[4], b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_936(w_eco936, a[3], b[4], !a[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_937(w_eco937, !b[3], b[4], !a[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_938(w_eco938, a[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_939(w_eco939, !b[3], a[4], !b[4], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_940(w_eco940, b[3], a[4], !b[5], a[6], !b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_941(w_eco941, b[3], a[4], !b[5], a[6], !b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_942(w_eco942, b[3], a[4], !b[5], a[6], !b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_943(w_eco943, b[3], a[4], !b[5], a[6], !b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_944(w_eco944, a[4], !b[4], !b[5], a[6], !b[6], a[7], !b[7], op[0], !op[1]);
	and _ECO_945(w_eco945, a[4], !b[5], a[6], !b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_946(w_eco946, a[4], !b[5], a[6], !b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_947(w_eco947, a[4], !b[5], a[6], !b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_948(w_eco948, a[3], !a[4], !a[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_949(w_eco949, !b[3], !a[4], !a[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_950(w_eco950, b[3], !b[4], !b[5], !a[6], b[6], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_951(w_eco951, b[3], !b[4], !b[5], !a[6], b[6], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_952(w_eco952, b[3], !b[4], !b[5], !a[6], b[6], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_953(w_eco953, b[3], !b[4], !b[5], !a[6], b[6], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_954(w_eco954, !b[4], !b[5], !a[6], b[6], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_955(w_eco955, !b[4], !b[5], !a[6], b[6], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_956(w_eco956, !b[4], !b[5], !a[6], b[6], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_957(w_eco957, !b[4], !b[5], !a[6], b[6], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_958(w_eco958, !b[4], !b[5], !a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_959(w_eco959, !b[4], !b[5], !a[6], b[6], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_960(w_eco960, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_961(w_eco961, !a[4], !b[4], !a[5], !b[5], a[6], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_962(w_eco962, a[3], !a[4], !a[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_963(w_eco963, !b[3], !a[4], !a[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_964(w_eco964, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_965(w_eco965, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_966(w_eco966, !b[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_967(w_eco967, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_968(w_eco968, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_969(w_eco969, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_970(w_eco970, !a[3], a[4], b[4], a[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_971(w_eco971, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_972(w_eco972, !b[3], a[4], b[4], a[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_973(w_eco973, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_974(w_eco974, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_975(w_eco975, !a[3], a[4], b[4], a[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_976(w_eco976, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_977(w_eco977, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_978(w_eco978, b[3], a[4], a[5], !a[6], b[6], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_979(w_eco979, b[3], a[4], a[5], !a[6], b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_980(w_eco980, b[3], a[4], a[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_981(w_eco981, b[3], a[4], a[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_982(w_eco982, a[4], a[5], !a[6], b[6], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_983(w_eco983, a[4], a[5], !a[6], b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_984(w_eco984, a[4], a[5], !a[6], b[6], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_985(w_eco985, a[4], a[5], !a[6], b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_986(w_eco986, !a[3], a[4], a[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_987(w_eco987, !a[3], a[4], a[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_988(w_eco988, a[4], a[5], !a[6], b[6], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_989(w_eco989, a[4], a[5], !a[6], b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_990(w_eco990, a[4], a[5], !a[6], b[6], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_991(w_eco991, a[4], a[5], !a[6], b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_992(w_eco992, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_993(w_eco993, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_994(w_eco994, !b[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_995(w_eco995, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_996(w_eco996, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_997(w_eco997, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_998(w_eco998, !a[3], a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_999(w_eco999, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1000(w_eco1000, !b[3], a[5], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1001(w_eco1001, !b[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1002(w_eco1002, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1003(w_eco1003, !a[3], a[5], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1004(w_eco1004, !a[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1005(w_eco1005, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1006(w_eco1006, b[3], a[4], a[5], a[6], !b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1007(w_eco1007, b[3], a[4], a[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1008(w_eco1008, a[4], a[5], a[6], !b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1009(w_eco1009, a[4], a[5], a[6], !b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1010(w_eco1010, !a[3], a[4], a[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1011(w_eco1011, a[4], a[5], a[6], !b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1012(w_eco1012, a[4], a[5], a[6], !b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1013(w_eco1013, b[3], !b[4], a[5], !a[6], b[6], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1014(w_eco1014, b[3], !b[4], a[5], !a[6], b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1015(w_eco1015, b[3], !b[4], a[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1016(w_eco1016, b[3], !b[4], a[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1017(w_eco1017, !b[4], a[5], !a[6], b[6], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1018(w_eco1018, !b[4], a[5], !a[6], b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1019(w_eco1019, !b[4], a[5], !a[6], b[6], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1020(w_eco1020, !b[4], a[5], !a[6], b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1021(w_eco1021, !a[3], !b[4], a[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1022(w_eco1022, !a[3], !b[4], a[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1023(w_eco1023, !b[4], a[5], !a[6], b[6], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1024(w_eco1024, !b[4], a[5], !a[6], b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1025(w_eco1025, !b[4], a[5], !a[6], b[6], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1026(w_eco1026, !b[4], a[5], !a[6], b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1027(w_eco1027, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[1]);
	and _ECO_1028(w_eco1028, !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1029(w_eco1029, !b[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1030(w_eco1030, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !b[2], !b[0], !b[7], !op[1]);
	and _ECO_1031(w_eco1031, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1032(w_eco1032, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1033(w_eco1033, !a[3], a[4], b[4], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1034(w_eco1034, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1035(w_eco1035, !b[3], a[4], b[4], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1036(w_eco1036, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[1]);
	and _ECO_1037(w_eco1037, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_1038(w_eco1038, !a[3], a[4], b[4], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1039(w_eco1039, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1040(w_eco1040, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1041(w_eco1041, a[3], !a[5], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1042(w_eco1042, a[3], !a[5], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1043(w_eco1043, a[3], !b[3], !a[5], b[5], a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1044(w_eco1044, !b[3], !a[5], b[5], a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1045(w_eco1045, !b[3], !a[5], b[5], a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1046(w_eco1046, a[3], !a[5], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1047(w_eco1047, a[3], !a[5], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1048(w_eco1048, a[3], !b[3], !a[5], b[5], !a[6], !b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1049(w_eco1049, !b[3], !a[5], b[5], !a[6], !b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1050(w_eco1050, !b[3], !a[5], b[5], !a[6], !b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1051(w_eco1051, a[3], a[5], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1052(w_eco1052, a[3], a[5], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1053(w_eco1053, a[3], !b[3], a[5], !b[5], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1054(w_eco1054, !b[3], a[5], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1055(w_eco1055, !b[3], a[5], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1056(w_eco1056, b[3], a[5], !b[5], a[6], !b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1057(w_eco1057, b[3], a[5], !b[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1058(w_eco1058, a[5], !b[5], a[6], !b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1059(w_eco1059, a[5], !b[5], a[6], !b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1060(w_eco1060, !a[3], a[5], !b[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1061(w_eco1061, a[5], !b[5], a[6], !b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1062(w_eco1062, a[5], !b[5], a[6], !b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1063(w_eco1063, b[3], a[4], !b[5], !a[6], b[6], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1064(w_eco1064, b[3], a[4], !b[5], !a[6], b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1065(w_eco1065, b[3], a[4], !b[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1066(w_eco1066, b[3], a[4], !b[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1067(w_eco1067, a[4], !b[5], !a[6], b[6], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1068(w_eco1068, a[4], !b[5], !a[6], b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1069(w_eco1069, a[4], !b[5], !a[6], b[6], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1070(w_eco1070, a[4], !b[5], !a[6], b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1071(w_eco1071, !a[3], a[4], !b[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1072(w_eco1072, !a[3], a[4], !b[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1073(w_eco1073, a[4], !b[5], !a[6], b[6], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1074(w_eco1074, a[4], !b[5], !a[6], b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1075(w_eco1075, a[4], !b[5], !a[6], b[6], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1076(w_eco1076, a[4], !b[5], !a[6], b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1077(w_eco1077, b[3], a[4], !b[5], a[6], !b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1078(w_eco1078, b[3], a[4], !b[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1079(w_eco1079, a[4], !b[5], a[6], !b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1080(w_eco1080, a[4], !b[5], a[6], !b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1081(w_eco1081, !a[3], a[4], !b[5], a[6], !b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1082(w_eco1082, a[4], !b[5], a[6], !b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1083(w_eco1083, a[4], !b[5], a[6], !b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1084(w_eco1084, b[3], !b[4], !b[5], !a[6], b[6], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1085(w_eco1085, b[3], !b[4], !b[5], !a[6], b[6], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1086(w_eco1086, b[3], !b[4], !b[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1087(w_eco1087, b[3], !b[4], !b[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1088(w_eco1088, !b[4], !b[5], !a[6], b[6], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1089(w_eco1089, !b[4], !b[5], !a[6], b[6], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1090(w_eco1090, !b[4], !b[5], !a[6], b[6], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1091(w_eco1091, !b[4], !b[5], !a[6], b[6], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1092(w_eco1092, !a[3], !b[4], !b[5], !a[6], b[6], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1093(w_eco1093, !a[3], !b[4], !b[5], !a[6], b[6], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1094(w_eco1094, !b[4], !b[5], !a[6], b[6], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1095(w_eco1095, !b[4], !b[5], !a[6], b[6], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1096(w_eco1096, !b[4], !b[5], !a[6], b[6], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1097(w_eco1097, !b[4], !b[5], !a[6], b[6], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1098(w_eco1098, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1099(w_eco1099, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1100(w_eco1100, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1101(w_eco1101, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1102(w_eco1102, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1103(w_eco1103, !b[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1104(w_eco1104, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1105(w_eco1105, !a[3], a[4], b[4], a[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1106(w_eco1106, a[3], a[5], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1107(w_eco1107, !b[3], a[5], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1108(w_eco1108, a[5], !b[5], a[6], !b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1109(w_eco1109, a[5], !b[5], a[6], !b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1110(w_eco1110, a[4], a[5], !a[6], b[6], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1111(w_eco1111, a[4], a[5], !a[6], b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1112(w_eco1112, a[4], a[5], !a[6], b[6], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1113(w_eco1113, a[4], a[5], !a[6], b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1114(w_eco1114, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1115(w_eco1115, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1116(w_eco1116, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1117(w_eco1117, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1118(w_eco1118, !b[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1119(w_eco1119, !b[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1120(w_eco1120, !a[3], a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1121(w_eco1121, !a[3], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1122(w_eco1122, a[4], a[5], a[6], !b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1123(w_eco1123, a[4], a[5], a[6], !b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1124(w_eco1124, !b[4], a[5], !a[6], b[6], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1125(w_eco1125, !b[4], a[5], !a[6], b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1126(w_eco1126, !b[4], a[5], !a[6], b[6], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1127(w_eco1127, !b[4], a[5], !a[6], b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1128(w_eco1128, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[1]);
	and _ECO_1129(w_eco1129, !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1130(w_eco1130, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1131(w_eco1131, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1132(w_eco1132, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[1]);
	and _ECO_1133(w_eco1133, a[3], !b[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_1134(w_eco1134, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1135(w_eco1135, !a[3], a[4], b[4], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1136(w_eco1136, a[3], !a[5], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1137(w_eco1137, !b[3], !a[5], b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1138(w_eco1138, a[3], !a[5], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1139(w_eco1139, !b[3], !a[5], b[5], !a[6], !b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1140(w_eco1140, a[4], !b[5], !a[6], b[6], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1141(w_eco1141, a[4], !b[5], !a[6], b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1142(w_eco1142, a[4], !b[5], !a[6], b[6], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1143(w_eco1143, a[4], !b[5], !a[6], b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1144(w_eco1144, a[4], !b[5], a[6], !b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1145(w_eco1145, a[4], !b[5], a[6], !b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1146(w_eco1146, !b[4], !b[5], !a[6], b[6], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1147(w_eco1147, !b[4], !b[5], !a[6], b[6], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1148(w_eco1148, !b[4], !b[5], !a[6], b[6], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1149(w_eco1149, !b[4], !b[5], !a[6], b[6], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	or _ECO_1150(w_eco1150, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149);
	xor _ECO_out3(y[6], sub_wire3, w_eco1150);
	and _ECO_1151(w_eco1151, !a[4], !b[4], !a[5], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1152(w_eco1152, !a[4], !b[4], a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1153(w_eco1153, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1154(w_eco1154, !a[3], a[4], !a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1155(w_eco1155, !a[3], a[4], !a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1156(w_eco1156, !a[4], !b[4], !a[5], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1157(w_eco1157, !a[3], !b[4], !a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1158(w_eco1158, !a[3], !b[4], !a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1159(w_eco1159, !a[3], a[4], a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1160(w_eco1160, !a[3], a[4], a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1161(w_eco1161, !a[4], !b[4], a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1162(w_eco1162, !a[3], !b[4], a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1163(w_eco1163, !a[3], !b[4], a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1164(w_eco1164, a[4], b[4], !a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1165(w_eco1165, !a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1166(w_eco1166, !a[3], !a[4], b[4], a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1167(w_eco1167, !a[3], !a[4], b[4], a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1168(w_eco1168, !a[3], b[3], a[4], !a[5], b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1169(w_eco1169, !a[3], b[3], a[4], !a[5], b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1170(w_eco1170, b[3], a[4], !a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1171(w_eco1171, b[3], a[4], !a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1172(w_eco1172, !a[3], b[3], !b[4], !a[5], b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1173(w_eco1173, !a[3], b[3], !b[4], !a[5], b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1174(w_eco1174, b[3], !b[4], !a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1175(w_eco1175, b[3], !b[4], !a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1176(w_eco1176, !a[3], b[3], a[4], a[5], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1177(w_eco1177, !a[3], b[3], a[4], a[5], !b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1178(w_eco1178, b[3], a[4], a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1179(w_eco1179, b[3], a[4], a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1180(w_eco1180, !a[3], b[3], !b[4], a[5], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1181(w_eco1181, !a[3], b[3], !b[4], a[5], !b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1182(w_eco1182, b[3], !b[4], a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1183(w_eco1183, b[3], !b[4], a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1184(w_eco1184, !a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1185(w_eco1185, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_1186(w_eco1186, !a[3], b[3], !a[4], b[4], a[5], b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1187(w_eco1187, !a[3], b[3], !a[4], b[4], a[5], b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1188(w_eco1188, b[3], !a[4], b[4], a[5], b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1189(w_eco1189, b[3], !a[4], b[4], a[5], b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1190(w_eco1190, !a[3], !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1191(w_eco1191, !a[3], !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1192(w_eco1192, !a[3], !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1193(w_eco1193, a[4], !b[4], a[5], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1194(w_eco1194, a[4], !b[4], a[5], !b[5], b[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_1195(w_eco1195, !a[3], !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1196(w_eco1196, a[4], !b[4], a[5], !b[5], !a[6], !a[7], b[7], op[0], !op[1]);
	and _ECO_1197(w_eco1197, !a[3], !a[4], b[4], !a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1198(w_eco1198, !a[3], !a[4], b[4], !a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1199(w_eco1199, a[3], b[3], b[4], !a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1200(w_eco1200, a[3], b[3], a[4], !a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1201(w_eco1201, a[3], !b[3], b[4], a[5], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1202(w_eco1202, a[3], !b[3], b[4], a[5], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1203(w_eco1203, a[3], !b[3], b[4], a[5], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1204(w_eco1204, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1205(w_eco1205, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1206(w_eco1206, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_1207(w_eco1207, a[3], !b[3], !a[4], a[5], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1208(w_eco1208, a[3], !b[3], !a[4], a[5], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1209(w_eco1209, a[3], !b[3], !a[4], a[5], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1210(w_eco1210, b[3], a[4], !a[5], b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1211(w_eco1211, b[3], a[4], !a[5], b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1212(w_eco1212, a[4], !a[5], b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1213(w_eco1213, a[4], !a[5], b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1214(w_eco1214, !a[3], !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1215(w_eco1215, !a[3], !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1216(w_eco1216, b[3], !b[4], !a[5], b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1217(w_eco1217, b[3], !b[4], !a[5], b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1218(w_eco1218, !b[4], !a[5], b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1219(w_eco1219, !b[4], !a[5], b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1220(w_eco1220, b[3], a[4], a[5], !b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1221(w_eco1221, b[3], a[4], a[5], !b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1222(w_eco1222, a[4], a[5], !b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1223(w_eco1223, a[4], a[5], !b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1224(w_eco1224, !a[3], !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1225(w_eco1225, !a[3], !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1226(w_eco1226, b[3], !b[4], a[5], !b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1227(w_eco1227, b[3], !b[4], a[5], !b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1228(w_eco1228, !b[4], a[5], !b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1229(w_eco1229, !b[4], a[5], !b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1230(w_eco1230, a[3], !b[3], b[4], !a[5], !b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1231(w_eco1231, a[3], !b[3], b[4], !a[5], !b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1232(w_eco1232, a[3], !b[3], b[4], !a[5], !b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1233(w_eco1233, !a[3], b[3], !a[4], b[4], !a[5], !b[5], a[7], !b[7], op[0], !op[1]);
	and _ECO_1234(w_eco1234, !a[3], b[3], !a[4], b[4], !a[5], !b[5], !a[7], b[7], op[0], !op[1]);
	and _ECO_1235(w_eco1235, b[3], !a[4], b[4], !a[5], !b[5], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1236(w_eco1236, b[3], !a[4], b[4], !a[5], !b[5], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1237(w_eco1237, a[3], b[3], b[4], !a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1238(w_eco1238, a[3], b[3], a[4], !a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1239(w_eco1239, a[3], !b[3], !a[4], !a[5], !b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1240(w_eco1240, a[3], !b[3], !a[4], !a[5], !b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1241(w_eco1241, a[3], !b[3], !a[4], !a[5], !b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1242(w_eco1242, a[3], b[4], a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1243(w_eco1243, a[3], b[4], a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1244(w_eco1244, a[3], !b[3], b[4], a[5], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1245(w_eco1245, !b[3], b[4], a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1246(w_eco1246, !b[3], b[4], a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1247(w_eco1247, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1248(w_eco1248, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1249(w_eco1249, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1250(w_eco1250, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[1]);
	and _ECO_1251(w_eco1251, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1252(w_eco1252, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1253(w_eco1253, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1254(w_eco1254, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1255(w_eco1255, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1256(w_eco1256, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1257(w_eco1257, a[3], !b[3], b[4], a[5], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1258(w_eco1258, a[3], !b[3], b[4], a[5], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1259(w_eco1259, a[3], !b[3], b[4], a[5], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1260(w_eco1260, b[3], !a[4], b[4], a[5], b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1261(w_eco1261, b[3], !a[4], b[4], a[5], b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1262(w_eco1262, !a[4], b[4], a[5], b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1263(w_eco1263, !a[4], b[4], a[5], b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1264(w_eco1264, a[3], !a[4], a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1265(w_eco1265, a[3], !a[4], a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1266(w_eco1266, a[3], !b[3], !a[4], a[5], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1267(w_eco1267, !b[3], !a[4], a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1268(w_eco1268, !b[3], !a[4], a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1269(w_eco1269, a[3], !b[3], !a[4], a[5], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1270(w_eco1270, a[3], !b[3], !a[4], a[5], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1271(w_eco1271, a[3], !b[3], !a[4], a[5], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1272(w_eco1272, b[3], a[4], !a[5], b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1273(w_eco1273, b[3], a[4], !a[5], b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1274(w_eco1274, b[3], a[4], !a[5], b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1275(w_eco1275, b[3], a[4], !a[5], b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1276(w_eco1276, a[4], !a[5], b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1277(w_eco1277, a[4], !a[5], b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1278(w_eco1278, a[4], !a[5], b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1279(w_eco1279, a[4], !a[5], b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1280(w_eco1280, a[4], !a[5], b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1281(w_eco1281, a[4], !a[5], b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1282(w_eco1282, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1283(w_eco1283, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1284(w_eco1284, a[3], !b[3], a[4], !b[4], !a[5], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1285(w_eco1285, a[3], !b[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1286(w_eco1286, a[3], !b[3], a[4], !b[4], !a[5], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1287(w_eco1287, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1288(w_eco1288, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1289(w_eco1289, a[3], !b[3], a[4], !b[4], !a[5], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1290(w_eco1290, a[3], !b[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1291(w_eco1291, a[3], !b[3], a[4], !b[4], !a[5], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1292(w_eco1292, b[3], !b[4], !a[5], b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1293(w_eco1293, b[3], !b[4], !a[5], b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1294(w_eco1294, b[3], !b[4], !a[5], b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1295(w_eco1295, b[3], !b[4], !a[5], b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1296(w_eco1296, !b[4], !a[5], b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1297(w_eco1297, !b[4], !a[5], b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1298(w_eco1298, !b[4], !a[5], b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1299(w_eco1299, !b[4], !a[5], b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1300(w_eco1300, !b[4], !a[5], b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1301(w_eco1301, !b[4], !a[5], b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1302(w_eco1302, b[3], a[4], a[5], !b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1303(w_eco1303, b[3], a[4], a[5], !b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1304(w_eco1304, b[3], a[4], a[5], !b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1305(w_eco1305, b[3], a[4], a[5], !b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1306(w_eco1306, a[4], a[5], !b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1307(w_eco1307, a[4], a[5], !b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1308(w_eco1308, a[4], a[5], !b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1309(w_eco1309, a[4], a[5], !b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1310(w_eco1310, a[4], a[5], !b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1311(w_eco1311, a[4], a[5], !b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1312(w_eco1312, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1313(w_eco1313, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1314(w_eco1314, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1315(w_eco1315, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1316(w_eco1316, b[3], !b[4], a[5], !b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1317(w_eco1317, b[3], !b[4], a[5], !b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1318(w_eco1318, b[3], !b[4], a[5], !b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1319(w_eco1319, b[3], !b[4], a[5], !b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1320(w_eco1320, !b[4], a[5], !b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1321(w_eco1321, !b[4], a[5], !b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1322(w_eco1322, !b[4], a[5], !b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1323(w_eco1323, !b[4], a[5], !b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1324(w_eco1324, !b[4], a[5], !b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1325(w_eco1325, !b[4], a[5], !b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1326(w_eco1326, a[3], b[4], !a[5], !b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1327(w_eco1327, a[3], b[4], !a[5], !b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1328(w_eco1328, a[3], !b[3], b[4], !a[5], !b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1329(w_eco1329, !b[3], b[4], !a[5], !b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1330(w_eco1330, !b[3], b[4], !a[5], !b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1331(w_eco1331, a[3], !b[3], b[4], !a[5], !b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1332(w_eco1332, a[3], !b[3], b[4], !a[5], !b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1333(w_eco1333, a[3], !b[3], b[4], !a[5], !b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1334(w_eco1334, a[3], !a[4], !a[5], !b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1335(w_eco1335, a[3], !a[4], !a[5], !b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1336(w_eco1336, a[3], !b[3], !a[4], !a[5], !b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1337(w_eco1337, !b[3], !a[4], !a[5], !b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1338(w_eco1338, !b[3], !a[4], !a[5], !b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1339(w_eco1339, a[3], !b[3], !a[4], !a[5], !b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1340(w_eco1340, a[3], !b[3], !a[4], !a[5], !b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1341(w_eco1341, a[3], !b[3], !a[4], !a[5], !b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1342(w_eco1342, a[3], b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1343(w_eco1343, !b[3], b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1344(w_eco1344, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1345(w_eco1345, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_1346(w_eco1346, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1347(w_eco1347, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1348(w_eco1348, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1349(w_eco1349, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1350(w_eco1350, !b[3], a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1351(w_eco1351, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1352(w_eco1352, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], !b[7], !op[1]);
	and _ECO_1353(w_eco1353, !a[3], a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1354(w_eco1354, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1355(w_eco1355, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1356(w_eco1356, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1357(w_eco1357, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1358(w_eco1358, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1359(w_eco1359, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1360(w_eco1360, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1361(w_eco1361, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1362(w_eco1362, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1363(w_eco1363, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1364(w_eco1364, a[3], b[4], a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1365(w_eco1365, a[3], b[4], a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1366(w_eco1366, a[3], !b[3], b[4], a[5], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1367(w_eco1367, !b[3], b[4], a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1368(w_eco1368, !b[3], b[4], a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1369(w_eco1369, b[3], !a[4], b[4], a[5], b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1370(w_eco1370, b[3], !a[4], b[4], a[5], b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1371(w_eco1371, b[3], !a[4], b[4], a[5], b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1372(w_eco1372, b[3], !a[4], b[4], a[5], b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1373(w_eco1373, !a[4], b[4], a[5], b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1374(w_eco1374, !a[4], b[4], a[5], b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1375(w_eco1375, !a[4], b[4], a[5], b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1376(w_eco1376, !a[4], b[4], a[5], b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1377(w_eco1377, !a[4], b[4], a[5], b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1378(w_eco1378, !a[4], b[4], a[5], b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1379(w_eco1379, a[3], !a[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1380(w_eco1380, !b[3], !a[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1381(w_eco1381, a[3], !a[4], a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1382(w_eco1382, a[3], !a[4], a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1383(w_eco1383, a[3], !b[3], !a[4], a[5], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1384(w_eco1384, !b[3], !a[4], a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1385(w_eco1385, !b[3], !a[4], a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1386(w_eco1386, b[3], a[4], !a[5], b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1387(w_eco1387, b[3], a[4], !a[5], b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1388(w_eco1388, b[3], a[4], !a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1389(w_eco1389, b[3], a[4], !a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1390(w_eco1390, a[4], !a[5], b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1391(w_eco1391, a[4], !a[5], b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1392(w_eco1392, a[4], !a[5], b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1393(w_eco1393, a[4], !a[5], b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1394(w_eco1394, !a[3], a[4], !a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1395(w_eco1395, !a[3], a[4], !a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1396(w_eco1396, a[4], !a[5], b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1397(w_eco1397, a[4], !a[5], b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1398(w_eco1398, a[4], !a[5], b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1399(w_eco1399, a[4], !a[5], b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1400(w_eco1400, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1401(w_eco1401, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1402(w_eco1402, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1403(w_eco1403, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1404(w_eco1404, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1405(w_eco1405, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1406(w_eco1406, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1407(w_eco1407, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1408(w_eco1408, a[3], a[4], !b[4], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1409(w_eco1409, a[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1410(w_eco1410, a[3], !b[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1411(w_eco1411, !b[3], a[4], !b[4], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1412(w_eco1412, !b[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1413(w_eco1413, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1414(w_eco1414, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1415(w_eco1415, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1416(w_eco1416, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1417(w_eco1417, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1418(w_eco1418, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1419(w_eco1419, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1420(w_eco1420, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1421(w_eco1421, a[3], a[4], !b[4], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1422(w_eco1422, a[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1423(w_eco1423, a[3], !b[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1424(w_eco1424, !b[3], a[4], !b[4], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1425(w_eco1425, !b[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1426(w_eco1426, b[3], !b[4], !a[5], b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1427(w_eco1427, b[3], !b[4], !a[5], b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1428(w_eco1428, b[3], !b[4], !a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1429(w_eco1429, b[3], !b[4], !a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1430(w_eco1430, !b[4], !a[5], b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1431(w_eco1431, !b[4], !a[5], b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1432(w_eco1432, !b[4], !a[5], b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1433(w_eco1433, !b[4], !a[5], b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1434(w_eco1434, !a[3], !b[4], !a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1435(w_eco1435, !a[3], !b[4], !a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1436(w_eco1436, !b[4], !a[5], b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1437(w_eco1437, !b[4], !a[5], b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1438(w_eco1438, !b[4], !a[5], b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1439(w_eco1439, !b[4], !a[5], b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1440(w_eco1440, b[3], a[4], a[5], !b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1441(w_eco1441, b[3], a[4], a[5], !b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1442(w_eco1442, b[3], a[4], a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1443(w_eco1443, b[3], a[4], a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1444(w_eco1444, a[4], a[5], !b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1445(w_eco1445, a[4], a[5], !b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1446(w_eco1446, a[4], a[5], !b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1447(w_eco1447, a[4], a[5], !b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1448(w_eco1448, !a[3], a[4], a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1449(w_eco1449, !a[3], a[4], a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1450(w_eco1450, a[4], a[5], !b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1451(w_eco1451, a[4], a[5], !b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1452(w_eco1452, a[4], a[5], !b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1453(w_eco1453, a[4], a[5], !b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1454(w_eco1454, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1455(w_eco1455, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1456(w_eco1456, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1457(w_eco1457, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1458(w_eco1458, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1459(w_eco1459, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1460(w_eco1460, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1461(w_eco1461, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1462(w_eco1462, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1463(w_eco1463, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1464(w_eco1464, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1465(w_eco1465, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1466(w_eco1466, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1467(w_eco1467, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1468(w_eco1468, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1469(w_eco1469, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1470(w_eco1470, b[3], !b[4], a[5], !b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1471(w_eco1471, b[3], !b[4], a[5], !b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1472(w_eco1472, b[3], !b[4], a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1473(w_eco1473, b[3], !b[4], a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1474(w_eco1474, !b[4], a[5], !b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1475(w_eco1475, !b[4], a[5], !b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1476(w_eco1476, !b[4], a[5], !b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1477(w_eco1477, !b[4], a[5], !b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1478(w_eco1478, !a[3], !b[4], a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1479(w_eco1479, !a[3], !b[4], a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1480(w_eco1480, !b[4], a[5], !b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1481(w_eco1481, !b[4], a[5], !b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1482(w_eco1482, !b[4], a[5], !b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1483(w_eco1483, !b[4], a[5], !b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1484(w_eco1484, a[3], b[4], !a[5], !b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1485(w_eco1485, !b[3], b[4], !a[5], !b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1486(w_eco1486, a[3], b[4], !a[5], !b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1487(w_eco1487, a[3], b[4], !a[5], !b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1488(w_eco1488, a[3], !b[3], b[4], !a[5], !b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1489(w_eco1489, !b[3], b[4], !a[5], !b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1490(w_eco1490, !b[3], b[4], !a[5], !b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1491(w_eco1491, b[3], !a[4], b[4], !a[5], !b[5], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1492(w_eco1492, b[3], !a[4], b[4], !a[5], !b[5], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1493(w_eco1493, !a[4], b[4], !a[5], !b[5], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1494(w_eco1494, !a[4], b[4], !a[5], !b[5], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1495(w_eco1495, a[3], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1496(w_eco1496, a[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1497(w_eco1497, a[3], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1498(w_eco1498, b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1499(w_eco1499, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1500(w_eco1500, b[3], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1501(w_eco1501, a[3], a[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1502(w_eco1502, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1503(w_eco1503, a[3], a[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1504(w_eco1504, b[3], a[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1505(w_eco1505, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1506(w_eco1506, b[3], a[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1507(w_eco1507, a[3], !a[4], !a[5], !b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1508(w_eco1508, !b[3], !a[4], !a[5], !b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1509(w_eco1509, a[3], !a[4], !a[5], !b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1510(w_eco1510, a[3], !a[4], !a[5], !b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1511(w_eco1511, a[3], !b[3], !a[4], !a[5], !b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1512(w_eco1512, !b[3], !a[4], !a[5], !b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1513(w_eco1513, !b[3], !a[4], !a[5], !b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1514(w_eco1514, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[1]);
	and _ECO_1515(w_eco1515, !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1516(w_eco1516, !b[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1517(w_eco1517, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], !b[7], !op[1]);
	and _ECO_1518(w_eco1518, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1519(w_eco1519, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1520(w_eco1520, !a[3], a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1521(w_eco1521, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1522(w_eco1522, !b[3], a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1523(w_eco1523, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[1]);
	and _ECO_1524(w_eco1524, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_1525(w_eco1525, !a[3], a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1526(w_eco1526, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1527(w_eco1527, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1528(w_eco1528, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1529(w_eco1529, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1530(w_eco1530, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1531(w_eco1531, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1532(w_eco1532, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1533(w_eco1533, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1534(w_eco1534, !b[3], a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1535(w_eco1535, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1536(w_eco1536, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1537(w_eco1537, !a[3], a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1538(w_eco1538, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1539(w_eco1539, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1540(w_eco1540, a[3], b[4], a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1541(w_eco1541, !b[3], b[4], a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1542(w_eco1542, b[3], !a[4], b[4], a[5], b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1543(w_eco1543, b[3], !a[4], b[4], a[5], b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1544(w_eco1544, b[3], !a[4], b[4], a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1545(w_eco1545, b[3], !a[4], b[4], a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1546(w_eco1546, !a[4], b[4], a[5], b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1547(w_eco1547, !a[4], b[4], a[5], b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1548(w_eco1548, !a[4], b[4], a[5], b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1549(w_eco1549, !a[4], b[4], a[5], b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1550(w_eco1550, !a[3], !a[4], b[4], a[5], b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1551(w_eco1551, !a[3], !a[4], b[4], a[5], b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1552(w_eco1552, !a[4], b[4], a[5], b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1553(w_eco1553, !a[4], b[4], a[5], b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1554(w_eco1554, !a[4], b[4], a[5], b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1555(w_eco1555, !a[4], b[4], a[5], b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1556(w_eco1556, !a[4], b[4], a[5], b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1557(w_eco1557, !a[4], b[4], a[5], b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1558(w_eco1558, !a[4], b[4], a[5], b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1559(w_eco1559, !a[4], b[4], a[5], b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1560(w_eco1560, a[3], !a[4], a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1561(w_eco1561, !b[3], !a[4], a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1562(w_eco1562, a[4], !a[5], b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1563(w_eco1563, a[4], !a[5], b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1564(w_eco1564, a[4], !a[5], b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1565(w_eco1565, a[4], !a[5], b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1566(w_eco1566, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1567(w_eco1567, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1568(w_eco1568, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1569(w_eco1569, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1570(w_eco1570, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1571(w_eco1571, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1572(w_eco1572, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1573(w_eco1573, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1574(w_eco1574, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1575(w_eco1575, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1576(w_eco1576, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1577(w_eco1577, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1578(w_eco1578, a[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1579(w_eco1579, !b[3], a[4], !b[4], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1580(w_eco1580, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1581(w_eco1581, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1582(w_eco1582, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1583(w_eco1583, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1584(w_eco1584, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1585(w_eco1585, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1586(w_eco1586, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1587(w_eco1587, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1588(w_eco1588, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1589(w_eco1589, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1590(w_eco1590, !a[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1591(w_eco1591, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1592(w_eco1592, a[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1593(w_eco1593, !b[3], a[4], !b[4], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1594(w_eco1594, !b[4], !a[5], b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1595(w_eco1595, !b[4], !a[5], b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1596(w_eco1596, !b[4], !a[5], b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1597(w_eco1597, !b[4], !a[5], b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1598(w_eco1598, a[4], a[5], !b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1599(w_eco1599, a[4], a[5], !b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1600(w_eco1600, a[4], a[5], !b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1601(w_eco1601, a[4], a[5], !b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1602(w_eco1602, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1603(w_eco1603, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1604(w_eco1604, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1605(w_eco1605, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1606(w_eco1606, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1607(w_eco1607, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1608(w_eco1608, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1609(w_eco1609, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1610(w_eco1610, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1611(w_eco1611, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1612(w_eco1612, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1613(w_eco1613, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1614(w_eco1614, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1615(w_eco1615, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1616(w_eco1616, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1617(w_eco1617, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1618(w_eco1618, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1619(w_eco1619, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1620(w_eco1620, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1621(w_eco1621, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1622(w_eco1622, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1623(w_eco1623, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1624(w_eco1624, !a[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1625(w_eco1625, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1626(w_eco1626, a[3], !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1627(w_eco1627, a[3], !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1628(w_eco1628, a[3], !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1629(w_eco1629, !b[4], a[5], !b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1630(w_eco1630, !b[4], a[5], !b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1631(w_eco1631, !b[4], a[5], !b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1632(w_eco1632, !b[4], a[5], !b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1633(w_eco1633, a[3], b[4], !a[5], !b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1634(w_eco1634, !b[3], b[4], !a[5], !b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1635(w_eco1635, b[3], !a[4], b[4], !a[5], !b[5], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1636(w_eco1636, b[3], !a[4], b[4], !a[5], !b[5], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1637(w_eco1637, b[3], !a[4], b[4], !a[5], !b[5], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1638(w_eco1638, b[3], !a[4], b[4], !a[5], !b[5], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1639(w_eco1639, !a[4], b[4], !a[5], !b[5], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1640(w_eco1640, !a[4], b[4], !a[5], !b[5], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1641(w_eco1641, !a[4], b[4], !a[5], !b[5], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1642(w_eco1642, !a[4], b[4], !a[5], !b[5], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1643(w_eco1643, !a[4], b[4], !a[5], !b[5], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1644(w_eco1644, !a[4], b[4], !a[5], !b[5], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1645(w_eco1645, a[3], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1646(w_eco1646, a[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_1647(w_eco1647, a[3], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1648(w_eco1648, b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1649(w_eco1649, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_1650(w_eco1650, b[3], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1651(w_eco1651, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_1652(w_eco1652, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_1653(w_eco1653, b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1654(w_eco1654, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1655(w_eco1655, b[3], !a[4], b[4], !a[5], !b[5], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1656(w_eco1656, b[3], !a[4], b[4], !a[5], !b[5], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1657(w_eco1657, b[3], !a[4], b[4], !a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1658(w_eco1658, b[3], !a[4], b[4], !a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1659(w_eco1659, !a[4], b[4], !a[5], !b[5], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1660(w_eco1660, !a[4], b[4], !a[5], !b[5], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1661(w_eco1661, !a[4], b[4], !a[5], !b[5], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1662(w_eco1662, !a[4], b[4], !a[5], !b[5], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1663(w_eco1663, !a[3], !a[4], b[4], !a[5], !b[5], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1664(w_eco1664, !a[3], !a[4], b[4], !a[5], !b[5], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1665(w_eco1665, !a[4], b[4], !a[5], !b[5], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1666(w_eco1666, !a[4], b[4], !a[5], !b[5], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1667(w_eco1667, !a[4], b[4], !a[5], !b[5], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1668(w_eco1668, !a[4], b[4], !a[5], !b[5], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1669(w_eco1669, a[3], a[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1670(w_eco1670, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_1671(w_eco1671, a[3], a[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1672(w_eco1672, b[3], a[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1673(w_eco1673, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_1674(w_eco1674, b[3], a[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1675(w_eco1675, a[3], a[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1676(w_eco1676, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1677(w_eco1677, b[3], a[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1678(w_eco1678, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1679(w_eco1679, a[3], !a[4], !a[5], !b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1680(w_eco1680, !b[3], !a[4], !a[5], !b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1681(w_eco1681, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[1]);
	and _ECO_1682(w_eco1682, !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1683(w_eco1683, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1684(w_eco1684, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1685(w_eco1685, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[1]);
	and _ECO_1686(w_eco1686, a[3], !b[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_1687(w_eco1687, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1688(w_eco1688, !a[3], a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1689(w_eco1689, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1690(w_eco1690, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1691(w_eco1691, !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1692(w_eco1692, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1693(w_eco1693, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1694(w_eco1694, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1695(w_eco1695, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1696(w_eco1696, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1697(w_eco1697, !b[3], a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1698(w_eco1698, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1699(w_eco1699, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1700(w_eco1700, !a[3], a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1701(w_eco1701, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1702(w_eco1702, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1703(w_eco1703, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1704(w_eco1704, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1705(w_eco1705, !b[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1706(w_eco1706, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1707(w_eco1707, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1708(w_eco1708, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1709(w_eco1709, !a[3], !a[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1710(w_eco1710, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1711(w_eco1711, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1712(w_eco1712, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1713(w_eco1713, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1714(w_eco1714, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1715(w_eco1715, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1716(w_eco1716, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1717(w_eco1717, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1718(w_eco1718, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1719(w_eco1719, !b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1720(w_eco1720, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1721(w_eco1721, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1722(w_eco1722, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1723(w_eco1723, !a[3], b[3], !b[4], !a[5], b[5], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1724(w_eco1724, !a[3], b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1725(w_eco1725, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1726(w_eco1726, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1727(w_eco1727, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1728(w_eco1728, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_1729(w_eco1729, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1730(w_eco1730, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1731(w_eco1731, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1732(w_eco1732, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1733(w_eco1733, !b[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1734(w_eco1734, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1735(w_eco1735, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1736(w_eco1736, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1737(w_eco1737, !a[3], !a[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1738(w_eco1738, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1739(w_eco1739, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1740(w_eco1740, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1741(w_eco1741, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1742(w_eco1742, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1743(w_eco1743, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1744(w_eco1744, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1745(w_eco1745, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1746(w_eco1746, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1747(w_eco1747, !b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1748(w_eco1748, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1749(w_eco1749, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1750(w_eco1750, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1751(w_eco1751, !a[3], b[3], !b[4], a[5], !b[5], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1752(w_eco1752, !a[3], b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1753(w_eco1753, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1754(w_eco1754, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1755(w_eco1755, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1756(w_eco1756, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_1757(w_eco1757, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1758(w_eco1758, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_1759(w_eco1759, a[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1760(w_eco1760, a[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1761(w_eco1761, a[3], !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1762(w_eco1762, !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1763(w_eco1763, !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1764(w_eco1764, a[3], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1765(w_eco1765, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1766(w_eco1766, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_1767(w_eco1767, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_1768(w_eco1768, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_1769(w_eco1769, b[3], b[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1770(w_eco1770, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1771(w_eco1771, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1772(w_eco1772, !a[4], b[4], !a[5], !b[5], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1773(w_eco1773, !a[4], b[4], !a[5], !b[5], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1774(w_eco1774, !a[4], b[4], !a[5], !b[5], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1775(w_eco1775, !a[4], b[4], !a[5], !b[5], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1776(w_eco1776, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1777(w_eco1777, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1778(w_eco1778, a[3], a[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1779(w_eco1779, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1780(w_eco1780, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1781(w_eco1781, b[3], a[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1782(w_eco1782, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1783(w_eco1783, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_1784(w_eco1784, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1785(w_eco1785, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1786(w_eco1786, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1787(w_eco1787, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1788(w_eco1788, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1789(w_eco1789, !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1790(w_eco1790, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1791(w_eco1791, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1792(w_eco1792, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1793(w_eco1793, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1794(w_eco1794, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1795(w_eco1795, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1796(w_eco1796, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1797(w_eco1797, !b[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1798(w_eco1798, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1799(w_eco1799, !a[3], !a[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1800(w_eco1800, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1801(w_eco1801, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_1802(w_eco1802, !a[3], b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1803(w_eco1803, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_1804(w_eco1804, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1805(w_eco1805, !b[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1806(w_eco1806, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1807(w_eco1807, !a[3], !b[4], !a[5], b[5], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_1808(w_eco1808, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1809(w_eco1809, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1810(w_eco1810, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1811(w_eco1811, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_1812(w_eco1812, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1813(w_eco1813, !b[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1814(w_eco1814, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1815(w_eco1815, !a[3], !a[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1816(w_eco1816, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1817(w_eco1817, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_1818(w_eco1818, !a[3], b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1819(w_eco1819, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_1820(w_eco1820, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1821(w_eco1821, !b[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_1822(w_eco1822, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1823(w_eco1823, !a[3], !b[4], a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_1824(w_eco1824, a[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1825(w_eco1825, !b[3], a[4], !b[4], a[5], !b[5], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1826(w_eco1826, a[3], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1827(w_eco1827, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1828(w_eco1828, a[3], !b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_1829(w_eco1829, b[3], b[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1830(w_eco1830, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1831(w_eco1831, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1832(w_eco1832, a[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_1833(w_eco1833, b[3], a[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	or _ECO_1834(w_eco1834, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401, w_eco1402, w_eco1403, w_eco1404, w_eco1405, w_eco1406, w_eco1407, w_eco1408, w_eco1409, w_eco1410, w_eco1411, w_eco1412, w_eco1413, w_eco1414, w_eco1415, w_eco1416, w_eco1417, w_eco1418, w_eco1419, w_eco1420, w_eco1421, w_eco1422, w_eco1423, w_eco1424, w_eco1425, w_eco1426, w_eco1427, w_eco1428, w_eco1429, w_eco1430, w_eco1431, w_eco1432, w_eco1433, w_eco1434, w_eco1435, w_eco1436, w_eco1437, w_eco1438, w_eco1439, w_eco1440, w_eco1441, w_eco1442, w_eco1443, w_eco1444, w_eco1445, w_eco1446, w_eco1447, w_eco1448, w_eco1449, w_eco1450, w_eco1451, w_eco1452, w_eco1453, w_eco1454, w_eco1455, w_eco1456, w_eco1457, w_eco1458, w_eco1459, w_eco1460, w_eco1461, w_eco1462, w_eco1463, w_eco1464, w_eco1465, w_eco1466, w_eco1467, w_eco1468, w_eco1469, w_eco1470, w_eco1471, w_eco1472, w_eco1473, w_eco1474, w_eco1475, w_eco1476, w_eco1477, w_eco1478, w_eco1479, w_eco1480, w_eco1481, w_eco1482, w_eco1483, w_eco1484, w_eco1485, w_eco1486, w_eco1487, w_eco1488, w_eco1489, w_eco1490, w_eco1491, w_eco1492, w_eco1493, w_eco1494, w_eco1495, w_eco1496, w_eco1497, w_eco1498, w_eco1499, w_eco1500, w_eco1501, w_eco1502, w_eco1503, w_eco1504, w_eco1505, w_eco1506, w_eco1507, w_eco1508, w_eco1509, w_eco1510, w_eco1511, w_eco1512, w_eco1513, w_eco1514, w_eco1515, w_eco1516, w_eco1517, w_eco1518, w_eco1519, w_eco1520, w_eco1521, w_eco1522, w_eco1523, w_eco1524, w_eco1525, w_eco1526, w_eco1527, w_eco1528, w_eco1529, w_eco1530, w_eco1531, w_eco1532, w_eco1533, w_eco1534, w_eco1535, w_eco1536, w_eco1537, w_eco1538, w_eco1539, w_eco1540, w_eco1541, w_eco1542, w_eco1543, w_eco1544, w_eco1545, w_eco1546, w_eco1547, w_eco1548, w_eco1549, w_eco1550, w_eco1551, w_eco1552, w_eco1553, w_eco1554, w_eco1555, w_eco1556, w_eco1557, w_eco1558, w_eco1559, w_eco1560, w_eco1561, w_eco1562, w_eco1563, w_eco1564, w_eco1565, w_eco1566, w_eco1567, w_eco1568, w_eco1569, w_eco1570, w_eco1571, w_eco1572, w_eco1573, w_eco1574, w_eco1575, w_eco1576, w_eco1577, w_eco1578, w_eco1579, w_eco1580, w_eco1581, w_eco1582, w_eco1583, w_eco1584, w_eco1585, w_eco1586, w_eco1587, w_eco1588, w_eco1589, w_eco1590, w_eco1591, w_eco1592, w_eco1593, w_eco1594, w_eco1595, w_eco1596, w_eco1597, w_eco1598, w_eco1599, w_eco1600, w_eco1601, w_eco1602, w_eco1603, w_eco1604, w_eco1605, w_eco1606, w_eco1607, w_eco1608, w_eco1609, w_eco1610, w_eco1611, w_eco1612, w_eco1613, w_eco1614, w_eco1615, w_eco1616, w_eco1617, w_eco1618, w_eco1619, w_eco1620, w_eco1621, w_eco1622, w_eco1623, w_eco1624, w_eco1625, w_eco1626, w_eco1627, w_eco1628, w_eco1629, w_eco1630, w_eco1631, w_eco1632, w_eco1633, w_eco1634, w_eco1635, w_eco1636, w_eco1637, w_eco1638, w_eco1639, w_eco1640, w_eco1641, w_eco1642, w_eco1643, w_eco1644, w_eco1645, w_eco1646, w_eco1647, w_eco1648, w_eco1649, w_eco1650, w_eco1651, w_eco1652, w_eco1653, w_eco1654, w_eco1655, w_eco1656, w_eco1657, w_eco1658, w_eco1659, w_eco1660, w_eco1661, w_eco1662, w_eco1663, w_eco1664, w_eco1665, w_eco1666, w_eco1667, w_eco1668, w_eco1669, w_eco1670, w_eco1671, w_eco1672, w_eco1673, w_eco1674, w_eco1675, w_eco1676, w_eco1677, w_eco1678, w_eco1679, w_eco1680, w_eco1681, w_eco1682, w_eco1683, w_eco1684, w_eco1685, w_eco1686, w_eco1687, w_eco1688, w_eco1689, w_eco1690, w_eco1691, w_eco1692, w_eco1693, w_eco1694, w_eco1695, w_eco1696, w_eco1697, w_eco1698, w_eco1699, w_eco1700, w_eco1701, w_eco1702, w_eco1703, w_eco1704, w_eco1705, w_eco1706, w_eco1707, w_eco1708, w_eco1709, w_eco1710, w_eco1711, w_eco1712, w_eco1713, w_eco1714, w_eco1715, w_eco1716, w_eco1717, w_eco1718, w_eco1719, w_eco1720, w_eco1721, w_eco1722, w_eco1723, w_eco1724, w_eco1725, w_eco1726, w_eco1727, w_eco1728, w_eco1729, w_eco1730, w_eco1731, w_eco1732, w_eco1733, w_eco1734, w_eco1735, w_eco1736, w_eco1737, w_eco1738, w_eco1739, w_eco1740, w_eco1741, w_eco1742, w_eco1743, w_eco1744, w_eco1745, w_eco1746, w_eco1747, w_eco1748, w_eco1749, w_eco1750, w_eco1751, w_eco1752, w_eco1753, w_eco1754, w_eco1755, w_eco1756, w_eco1757, w_eco1758, w_eco1759, w_eco1760, w_eco1761, w_eco1762, w_eco1763, w_eco1764, w_eco1765, w_eco1766, w_eco1767, w_eco1768, w_eco1769, w_eco1770, w_eco1771, w_eco1772, w_eco1773, w_eco1774, w_eco1775, w_eco1776, w_eco1777, w_eco1778, w_eco1779, w_eco1780, w_eco1781, w_eco1782, w_eco1783, w_eco1784, w_eco1785, w_eco1786, w_eco1787, w_eco1788, w_eco1789, w_eco1790, w_eco1791, w_eco1792, w_eco1793, w_eco1794, w_eco1795, w_eco1796, w_eco1797, w_eco1798, w_eco1799, w_eco1800, w_eco1801, w_eco1802, w_eco1803, w_eco1804, w_eco1805, w_eco1806, w_eco1807, w_eco1808, w_eco1809, w_eco1810, w_eco1811, w_eco1812, w_eco1813, w_eco1814, w_eco1815, w_eco1816, w_eco1817, w_eco1818, w_eco1819, w_eco1820, w_eco1821, w_eco1822, w_eco1823, w_eco1824, w_eco1825, w_eco1826, w_eco1827, w_eco1828, w_eco1829, w_eco1830, w_eco1831, w_eco1832, w_eco1833);
	xor _ECO_out4(y[5], sub_wire4, w_eco1834);
	and _ECO_1835(w_eco1835, !a[3], !a[4], b[4], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1836(w_eco1836, !a[3], !a[4], b[4], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1837(w_eco1837, !a[3], !b[3], !a[4], b[4], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1838(w_eco1838, !a[3], a[4], !b[4], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1839(w_eco1839, !a[3], a[4], !b[4], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1840(w_eco1840, !a[3], !b[3], a[4], !b[4], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1841(w_eco1841, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1842(w_eco1842, !a[3], b[3], !a[4], b[4], a[7], !b[7], op[0], !op[1]);
	and _ECO_1843(w_eco1843, !a[3], b[3], !a[4], b[4], !a[7], b[7], op[0], !op[1]);
	and _ECO_1844(w_eco1844, b[3], !a[4], b[4], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1845(w_eco1845, b[3], !a[4], b[4], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1846(w_eco1846, !a[3], !b[3], !a[4], b[4], a[5], b[5], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1847(w_eco1847, !a[3], !b[3], !a[4], b[4], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_1848(w_eco1848, !a[3], b[3], a[4], !b[4], a[7], !b[7], op[0], !op[1]);
	and _ECO_1849(w_eco1849, !a[3], b[3], a[4], !b[4], !a[7], b[7], op[0], !op[1]);
	and _ECO_1850(w_eco1850, b[3], a[4], !b[4], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_1851(w_eco1851, b[3], a[4], !b[4], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_1852(w_eco1852, !a[3], !b[3], a[4], !b[4], a[5], b[5], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1853(w_eco1853, !a[3], !b[3], a[4], !b[4], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_1854(w_eco1854, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1855(w_eco1855, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[7], !op[0], !op[1]);
	and _ECO_1856(w_eco1856, !a[3], !b[3], !a[4], b[4], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1857(w_eco1857, !a[3], !b[3], a[4], !b[4], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1858(w_eco1858, a[3], b[3], !a[4], !b[4], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1859(w_eco1859, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], !a[7], !op[0], !op[1]);
	and _ECO_1860(w_eco1860, a[3], !b[3], a[4], b[4], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1861(w_eco1861, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1862(w_eco1862, a[3], !b[3], a[4], b[4], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1863(w_eco1863, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1864(w_eco1864, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1865(w_eco1865, !a[3], !b[3], !a[4], b[4], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_1866(w_eco1866, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1867(w_eco1867, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1868(w_eco1868, !a[3], !b[3], a[4], !b[4], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_1869(w_eco1869, a[3], !b[3], !a[4], !b[4], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1870(w_eco1870, a[3], !b[3], !a[4], !b[4], b[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1871(w_eco1871, a[3], !b[3], !a[4], !b[4], b[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1872(w_eco1872, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[7], !op[0], !op[1]);
	and _ECO_1873(w_eco1873, !a[3], !b[3], !a[4], b[4], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1874(w_eco1874, !a[3], !b[3], a[4], !b[4], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1875(w_eco1875, a[3], b[3], !a[4], !b[4], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1876(w_eco1876, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], !b[7], !op[0], !op[1]);
	and _ECO_1877(w_eco1877, a[3], a[4], b[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1878(w_eco1878, a[3], a[4], b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1879(w_eco1879, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1880(w_eco1880, !b[3], a[4], b[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1881(w_eco1881, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1882(w_eco1882, a[3], !b[3], a[4], b[4], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1883(w_eco1883, a[3], !b[3], a[4], b[4], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1884(w_eco1884, a[3], !b[3], a[4], b[4], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1885(w_eco1885, b[3], !a[4], b[4], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1886(w_eco1886, b[3], !a[4], b[4], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1887(w_eco1887, !a[4], b[4], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1888(w_eco1888, !a[4], b[4], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1889(w_eco1889, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1890(w_eco1890, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1891(w_eco1891, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1892(w_eco1892, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1893(w_eco1893, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1894(w_eco1894, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1895(w_eco1895, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1896(w_eco1896, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1897(w_eco1897, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1898(w_eco1898, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1899(w_eco1899, b[3], a[4], !b[4], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1900(w_eco1900, b[3], a[4], !b[4], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1901(w_eco1901, a[4], !b[4], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1902(w_eco1902, a[4], !b[4], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1903(w_eco1903, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1904(w_eco1904, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1905(w_eco1905, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1906(w_eco1906, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1907(w_eco1907, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1908(w_eco1908, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1909(w_eco1909, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1910(w_eco1910, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1911(w_eco1911, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1912(w_eco1912, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1913(w_eco1913, a[3], !a[4], !b[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1914(w_eco1914, a[3], !a[4], !b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1915(w_eco1915, a[3], !b[3], !a[4], !b[4], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1916(w_eco1916, !b[3], !a[4], !b[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1917(w_eco1917, !b[3], !a[4], !b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1918(w_eco1918, a[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1919(w_eco1919, a[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1920(w_eco1920, a[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1921(w_eco1921, b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_1922(w_eco1922, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_1923(w_eco1923, b[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_1924(w_eco1924, a[3], !b[3], !a[4], !b[4], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1925(w_eco1925, a[3], !b[3], !a[4], !b[4], b[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1926(w_eco1926, a[3], !b[3], !a[4], !b[4], b[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1927(w_eco1927, !b[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1928(w_eco1928, !a[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1929(w_eco1929, !b[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1930(w_eco1930, !a[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1931(w_eco1931, a[3], !b[3], a[4], b[4], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1932(w_eco1932, a[3], !b[3], a[4], b[4], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1933(w_eco1933, a[3], !b[3], a[4], b[4], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1934(w_eco1934, a[3], !b[3], !a[4], !b[4], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1935(w_eco1935, a[3], !b[3], !a[4], !b[4], !a[6], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1936(w_eco1936, a[3], !b[3], !a[4], !b[4], !a[6], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1937(w_eco1937, a[3], !b[3], a[4], b[4], !a[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1938(w_eco1938, a[3], !b[3], a[4], b[4], !a[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1939(w_eco1939, a[3], !b[3], a[4], b[4], !a[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1940(w_eco1940, a[3], !b[3], a[4], b[4], !a[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1941(w_eco1941, a[3], !b[3], a[4], b[4], !a[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1942(w_eco1942, a[3], !b[3], a[4], b[4], !a[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1943(w_eco1943, a[3], !b[3], !a[4], !b[4], !a[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1944(w_eco1944, a[3], !b[3], !a[4], !b[4], !a[5], b[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1945(w_eco1945, a[3], !b[3], !a[4], !b[4], !a[5], b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1946(w_eco1946, a[3], !b[3], !a[4], !b[4], !a[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1947(w_eco1947, a[3], !b[3], !a[4], !b[4], !a[5], !a[6], !a[1], b[1], op[0], !op[1]);
	and _ECO_1948(w_eco1948, a[3], !b[3], !a[4], !b[4], !a[5], !a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_1949(w_eco1949, a[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1950(w_eco1950, !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1951(w_eco1951, a[3], a[4], b[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1952(w_eco1952, a[3], a[4], b[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1953(w_eco1953, a[3], !b[3], a[4], b[4], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_1954(w_eco1954, !b[3], a[4], b[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_1955(w_eco1955, !b[3], a[4], b[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_1956(w_eco1956, b[3], !a[4], b[4], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1957(w_eco1957, b[3], !a[4], b[4], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1958(w_eco1958, b[3], !a[4], b[4], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1959(w_eco1959, b[3], !a[4], b[4], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1960(w_eco1960, !a[4], b[4], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1961(w_eco1961, !a[4], b[4], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1962(w_eco1962, !a[4], b[4], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1963(w_eco1963, !a[4], b[4], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1964(w_eco1964, !a[4], b[4], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1965(w_eco1965, !a[4], b[4], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1966(w_eco1966, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1967(w_eco1967, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1968(w_eco1968, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1969(w_eco1969, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1970(w_eco1970, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1971(w_eco1971, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1972(w_eco1972, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1973(w_eco1973, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_1974(w_eco1974, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1975(w_eco1975, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_1976(w_eco1976, !a[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_1977(w_eco1977, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1978(w_eco1978, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1979(w_eco1979, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1980(w_eco1980, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1981(w_eco1981, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1982(w_eco1982, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_1983(w_eco1983, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1984(w_eco1984, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1985(w_eco1985, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1986(w_eco1986, b[3], a[4], !b[4], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1987(w_eco1987, b[3], a[4], !b[4], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1988(w_eco1988, b[3], a[4], !b[4], a[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1989(w_eco1989, b[3], a[4], !b[4], a[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1990(w_eco1990, a[4], !b[4], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1991(w_eco1991, a[4], !b[4], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1992(w_eco1992, a[4], !b[4], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1993(w_eco1993, a[4], !b[4], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1994(w_eco1994, a[4], !b[4], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_1995(w_eco1995, a[4], !b[4], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_1996(w_eco1996, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_1997(w_eco1997, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_1998(w_eco1998, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_1999(w_eco1999, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2000(w_eco2000, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2001(w_eco2001, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2002(w_eco2002, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2003(w_eco2003, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2004(w_eco2004, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2005(w_eco2005, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2006(w_eco2006, !a[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2007(w_eco2007, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2008(w_eco2008, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2009(w_eco2009, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2010(w_eco2010, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2011(w_eco2011, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2012(w_eco2012, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2013(w_eco2013, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2014(w_eco2014, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2015(w_eco2015, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2016(w_eco2016, a[3], !a[4], !b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2017(w_eco2017, !b[3], !a[4], !b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2018(w_eco2018, a[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2019(w_eco2019, a[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2020(w_eco2020, a[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2021(w_eco2021, b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2022(w_eco2022, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2023(w_eco2023, b[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2024(w_eco2024, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_2025(w_eco2025, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_2026(w_eco2026, b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2027(w_eco2027, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2028(w_eco2028, a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2029(w_eco2029, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2030(w_eco2030, a[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2031(w_eco2031, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2032(w_eco2032, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2033(w_eco2033, b[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2034(w_eco2034, a[3], !a[4], !b[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2035(w_eco2035, a[3], !a[4], !b[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2036(w_eco2036, a[3], !b[3], !a[4], !b[4], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2037(w_eco2037, !b[3], !a[4], !b[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2038(w_eco2038, !b[3], !a[4], !b[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2039(w_eco2039, !b[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2040(w_eco2040, !a[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2041(w_eco2041, !b[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2042(w_eco2042, !b[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2043(w_eco2043, !b[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2044(w_eco2044, !a[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2045(w_eco2045, !a[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2046(w_eco2046, !a[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2047(w_eco2047, !b[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2048(w_eco2048, !a[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2049(w_eco2049, !b[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2050(w_eco2050, !b[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2051(w_eco2051, !b[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2052(w_eco2052, !a[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2053(w_eco2053, !a[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2054(w_eco2054, !a[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2055(w_eco2055, a[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2056(w_eco2056, a[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2057(w_eco2057, a[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2058(w_eco2058, b[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2059(w_eco2059, b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2060(w_eco2060, b[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2061(w_eco2061, a[3], a[4], b[4], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2062(w_eco2062, a[3], a[4], b[4], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2063(w_eco2063, a[3], !b[3], a[4], b[4], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2064(w_eco2064, !b[3], a[4], b[4], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2065(w_eco2065, !b[3], a[4], b[4], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2066(w_eco2066, a[3], !a[4], !b[4], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2067(w_eco2067, a[3], !a[4], !b[4], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2068(w_eco2068, a[3], !b[3], !a[4], !b[4], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2069(w_eco2069, !b[3], !a[4], !b[4], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2070(w_eco2070, !b[3], !a[4], !b[4], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2071(w_eco2071, a[3], a[4], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2072(w_eco2072, a[3], a[4], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2073(w_eco2073, a[3], !b[3], a[4], b[4], !a[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2074(w_eco2074, !b[3], a[4], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2075(w_eco2075, !b[3], a[4], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2076(w_eco2076, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2077(w_eco2077, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2078(w_eco2078, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2079(w_eco2079, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2080(w_eco2080, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2081(w_eco2081, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2082(w_eco2082, a[3], a[4], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2083(w_eco2083, a[3], a[4], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2084(w_eco2084, a[3], !b[3], a[4], b[4], !a[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2085(w_eco2085, !b[3], a[4], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2086(w_eco2086, !b[3], a[4], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2087(w_eco2087, a[3], !a[4], !b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2088(w_eco2088, a[3], !a[4], !b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2089(w_eco2089, a[3], !b[3], !a[4], !b[4], !a[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2090(w_eco2090, !b[3], !a[4], !b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2091(w_eco2091, !b[3], !a[4], !b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2092(w_eco2092, a[3], !a[4], !b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2093(w_eco2093, a[3], !a[4], !b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2094(w_eco2094, a[3], !b[3], !a[4], !b[4], !a[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_2095(w_eco2095, !b[3], !a[4], !b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2096(w_eco2096, !b[3], !a[4], !b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2097(w_eco2097, a[3], a[4], b[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2098(w_eco2098, !b[3], a[4], b[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2099(w_eco2099, b[3], !a[4], b[4], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2100(w_eco2100, b[3], !a[4], b[4], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2101(w_eco2101, b[3], !a[4], b[4], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2102(w_eco2102, b[3], !a[4], b[4], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2103(w_eco2103, !a[4], b[4], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2104(w_eco2104, !a[4], b[4], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2105(w_eco2105, !a[4], b[4], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2106(w_eco2106, !a[4], b[4], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2107(w_eco2107, !a[3], !a[4], b[4], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2108(w_eco2108, !a[3], !a[4], b[4], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2109(w_eco2109, !a[4], b[4], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2110(w_eco2110, !a[4], b[4], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2111(w_eco2111, !a[4], b[4], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2112(w_eco2112, !a[4], b[4], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2113(w_eco2113, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2114(w_eco2114, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2115(w_eco2115, !b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2116(w_eco2116, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2117(w_eco2117, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2118(w_eco2118, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2119(w_eco2119, !a[3], b[3], !a[4], b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2120(w_eco2120, !a[3], b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2121(w_eco2121, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2122(w_eco2122, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2123(w_eco2123, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2124(w_eco2124, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2125(w_eco2125, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2126(w_eco2126, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2127(w_eco2127, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2128(w_eco2128, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2129(w_eco2129, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2130(w_eco2130, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2131(w_eco2131, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2132(w_eco2132, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2133(w_eco2133, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2134(w_eco2134, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2135(w_eco2135, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2136(w_eco2136, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2137(w_eco2137, !a[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2138(w_eco2138, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2139(w_eco2139, b[3], a[4], !b[4], a[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2140(w_eco2140, b[3], a[4], !b[4], a[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2141(w_eco2141, b[3], a[4], !b[4], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2142(w_eco2142, b[3], a[4], !b[4], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2143(w_eco2143, a[4], !b[4], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2144(w_eco2144, a[4], !b[4], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2145(w_eco2145, a[4], !b[4], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2146(w_eco2146, a[4], !b[4], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2147(w_eco2147, !a[3], a[4], !b[4], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2148(w_eco2148, !a[3], a[4], !b[4], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2149(w_eco2149, a[4], !b[4], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2150(w_eco2150, a[4], !b[4], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2151(w_eco2151, a[4], !b[4], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2152(w_eco2152, a[4], !b[4], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2153(w_eco2153, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2154(w_eco2154, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2155(w_eco2155, !b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2156(w_eco2156, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2157(w_eco2157, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2158(w_eco2158, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2159(w_eco2159, !a[3], b[3], a[4], !b[4], a[5], b[5], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2160(w_eco2160, !a[3], b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2161(w_eco2161, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2162(w_eco2162, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2163(w_eco2163, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2164(w_eco2164, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2165(w_eco2165, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2166(w_eco2166, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2167(w_eco2167, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2168(w_eco2168, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2169(w_eco2169, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2170(w_eco2170, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2171(w_eco2171, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2172(w_eco2172, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2173(w_eco2173, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2174(w_eco2174, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2175(w_eco2175, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2176(w_eco2176, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2177(w_eco2177, !a[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2178(w_eco2178, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2179(w_eco2179, a[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2180(w_eco2180, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2181(w_eco2181, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_2182(w_eco2182, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_2183(w_eco2183, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_2184(w_eco2184, b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2185(w_eco2185, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2186(w_eco2186, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2187(w_eco2187, a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2188(w_eco2188, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2189(w_eco2189, a[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2190(w_eco2190, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2191(w_eco2191, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2192(w_eco2192, b[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2193(w_eco2193, a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2194(w_eco2194, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2195(w_eco2195, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2196(w_eco2196, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2197(w_eco2197, a[3], !a[4], !b[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2198(w_eco2198, !b[3], !a[4], !b[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2199(w_eco2199, !b[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2200(w_eco2200, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2201(w_eco2201, !b[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2202(w_eco2202, !a[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2203(w_eco2203, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2204(w_eco2204, !a[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2205(w_eco2205, !b[3], !a[4], b[4], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2206(w_eco2206, !b[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2207(w_eco2207, !b[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2208(w_eco2208, !a[3], !a[4], b[4], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2209(w_eco2209, !a[3], !a[4], b[4], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2210(w_eco2210, !a[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2211(w_eco2211, !b[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2212(w_eco2212, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2213(w_eco2213, !b[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2214(w_eco2214, !a[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2215(w_eco2215, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2216(w_eco2216, !a[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2217(w_eco2217, !b[3], a[4], !b[4], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2218(w_eco2218, !b[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2219(w_eco2219, !b[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2220(w_eco2220, !a[3], a[4], !b[4], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2221(w_eco2221, !a[3], a[4], !b[4], a[6], b[6], !b[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2222(w_eco2222, !a[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2223(w_eco2223, a[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2224(w_eco2224, a[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2225(w_eco2225, a[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2226(w_eco2226, b[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2227(w_eco2227, b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2228(w_eco2228, b[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2229(w_eco2229, a[3], !a[4], !b[4], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2230(w_eco2230, a[3], !a[4], !b[4], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2231(w_eco2231, b[3], !a[4], !b[4], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2232(w_eco2232, b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2233(w_eco2233, a[3], !b[3], a[4], b[4], b[6], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2234(w_eco2234, a[3], !b[3], a[4], b[4], b[6], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2235(w_eco2235, a[3], !b[3], a[4], b[4], b[6], !a[1], b[1], a[7], !b[7], op[0], !op[1]);
	and _ECO_2236(w_eco2236, a[3], !b[3], a[4], b[4], b[6], !a[1], b[1], !a[7], b[7], op[0], !op[1]);
	and _ECO_2237(w_eco2237, a[3], !b[3], a[4], b[4], b[6], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2238(w_eco2238, a[3], !b[3], a[4], b[4], b[6], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2239(w_eco2239, a[3], a[4], b[4], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2240(w_eco2240, !b[3], a[4], b[4], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2241(w_eco2241, a[3], !b[3], a[4], b[4], a[5], !b[5], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2242(w_eco2242, a[3], !b[3], a[4], b[4], a[5], !b[5], !a[1], b[1], a[7], !b[7], op[0], !op[1]);
	and _ECO_2243(w_eco2243, a[3], !b[3], a[4], b[4], a[5], !b[5], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2244(w_eco2244, a[3], !b[3], a[4], b[4], !a[6], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2245(w_eco2245, a[3], !b[3], a[4], b[4], !a[6], !a[1], b[1], !a[7], b[7], op[0], !op[1]);
	and _ECO_2246(w_eco2246, a[3], !b[3], a[4], b[4], !a[6], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2247(w_eco2247, a[3], !b[3], !a[4], !b[4], b[6], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2248(w_eco2248, a[3], !b[3], !a[4], !b[4], b[6], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2249(w_eco2249, a[3], !b[3], !a[4], !b[4], b[6], !a[1], b[1], a[7], !b[7], op[0], !op[1]);
	and _ECO_2250(w_eco2250, a[3], !b[3], !a[4], !b[4], b[6], !a[1], b[1], !a[7], b[7], op[0], !op[1]);
	and _ECO_2251(w_eco2251, a[3], !b[3], !a[4], !b[4], b[6], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2252(w_eco2252, a[3], !b[3], !a[4], !b[4], b[6], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2253(w_eco2253, a[3], !a[4], !b[4], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2254(w_eco2254, !b[3], !a[4], !b[4], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2255(w_eco2255, a[3], !b[3], !a[4], !b[4], a[5], !b[5], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2256(w_eco2256, a[3], !b[3], !a[4], !b[4], a[5], !b[5], !a[1], b[1], a[7], !b[7], op[0], !op[1]);
	and _ECO_2257(w_eco2257, a[3], !b[3], !a[4], !b[4], a[5], !b[5], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2258(w_eco2258, a[3], !b[3], !a[4], !b[4], !a[6], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2259(w_eco2259, a[3], !b[3], !a[4], !b[4], !a[6], !a[1], b[1], !a[7], b[7], op[0], !op[1]);
	and _ECO_2260(w_eco2260, a[3], !b[3], !a[4], !b[4], !a[6], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2261(w_eco2261, a[3], a[4], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2262(w_eco2262, !b[3], a[4], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2263(w_eco2263, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2264(w_eco2264, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2265(w_eco2265, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2266(w_eco2266, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2267(w_eco2267, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2268(w_eco2268, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2269(w_eco2269, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_2270(w_eco2270, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_2271(w_eco2271, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2272(w_eco2272, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2273(w_eco2273, a[3], a[4], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2274(w_eco2274, !b[3], a[4], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2275(w_eco2275, a[3], !a[4], !b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2276(w_eco2276, !b[3], !a[4], !b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2277(w_eco2277, a[3], !a[4], !b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2278(w_eco2278, !b[3], !a[4], !b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2279(w_eco2279, !a[4], b[4], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2280(w_eco2280, !a[4], b[4], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2281(w_eco2281, !a[4], b[4], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2282(w_eco2282, !a[4], b[4], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2283(w_eco2283, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2284(w_eco2284, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2285(w_eco2285, !a[3], b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2286(w_eco2286, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2287(w_eco2287, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2288(w_eco2288, !b[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2289(w_eco2289, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2290(w_eco2290, !a[3], !a[4], b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2291(w_eco2291, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2292(w_eco2292, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2293(w_eco2293, !b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2294(w_eco2294, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2295(w_eco2295, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2296(w_eco2296, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2297(w_eco2297, !a[3], b[3], !a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2298(w_eco2298, !a[3], b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2299(w_eco2299, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2300(w_eco2300, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2301(w_eco2301, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2302(w_eco2302, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2303(w_eco2303, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2304(w_eco2304, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2305(w_eco2305, a[4], !b[4], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2306(w_eco2306, a[4], !b[4], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2307(w_eco2307, a[4], !b[4], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2308(w_eco2308, a[4], !b[4], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2309(w_eco2309, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2310(w_eco2310, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2311(w_eco2311, !a[3], b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2312(w_eco2312, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2313(w_eco2313, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2314(w_eco2314, !b[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2315(w_eco2315, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2316(w_eco2316, !a[3], a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2317(w_eco2317, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2318(w_eco2318, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2319(w_eco2319, !b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2320(w_eco2320, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2321(w_eco2321, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2322(w_eco2322, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2323(w_eco2323, !a[3], b[3], a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2324(w_eco2324, !a[3], b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2325(w_eco2325, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2326(w_eco2326, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2327(w_eco2327, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2328(w_eco2328, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2329(w_eco2329, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2330(w_eco2330, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2331(w_eco2331, a[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2332(w_eco2332, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2333(w_eco2333, a[3], !b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_2334(w_eco2334, b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2335(w_eco2335, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2336(w_eco2336, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2337(w_eco2337, a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2338(w_eco2338, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2339(w_eco2339, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2340(w_eco2340, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2341(w_eco2341, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2342(w_eco2342, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2343(w_eco2343, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2344(w_eco2344, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2345(w_eco2345, !b[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2346(w_eco2346, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2347(w_eco2347, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2348(w_eco2348, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2349(w_eco2349, !a[3], b[3], !a[4], b[4], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2350(w_eco2350, !a[3], b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2351(w_eco2351, !b[3], !a[4], b[4], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2352(w_eco2352, !b[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2353(w_eco2353, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2354(w_eco2354, !a[3], !a[4], b[4], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2355(w_eco2355, !a[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2356(w_eco2356, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2357(w_eco2357, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2358(w_eco2358, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2359(w_eco2359, !b[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2360(w_eco2360, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2361(w_eco2361, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2362(w_eco2362, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2363(w_eco2363, !a[3], b[3], a[4], !b[4], a[6], b[6], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2364(w_eco2364, !a[3], b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2365(w_eco2365, !b[3], a[4], !b[4], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2366(w_eco2366, !b[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2367(w_eco2367, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2368(w_eco2368, !a[3], a[4], !b[4], a[6], b[6], !a[2], !b[2], a[7], !b[7], !op[1]);
	and _ECO_2369(w_eco2369, !a[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2370(w_eco2370, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2371(w_eco2371, a[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2372(w_eco2372, b[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2373(w_eco2373, a[3], !b[3], !a[4], !b[4], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_2374(w_eco2374, a[3], !a[4], !b[4], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2375(w_eco2375, a[3], !b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_2376(w_eco2376, b[3], !a[4], !b[4], a[6], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2377(w_eco2377, b[3], !a[4], !b[4], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2378(w_eco2378, b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2379(w_eco2379, a[3], a[4], b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2380(w_eco2380, a[3], a[4], b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2381(w_eco2381, a[3], a[4], b[4], b[6], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2382(w_eco2382, a[3], a[4], b[4], b[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2383(w_eco2383, a[3], !b[3], a[4], b[4], b[6], !a[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2384(w_eco2384, a[3], !b[3], a[4], b[4], b[6], !a[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2385(w_eco2385, !b[3], a[4], b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2386(w_eco2386, !b[3], a[4], b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2387(w_eco2387, !b[3], a[4], b[4], b[6], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2388(w_eco2388, !b[3], a[4], b[4], b[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2389(w_eco2389, a[3], a[4], b[4], a[5], !b[5], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2390(w_eco2390, a[3], a[4], b[4], a[5], !b[5], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2391(w_eco2391, a[3], !b[3], a[4], b[4], a[5], !b[5], !a[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2392(w_eco2392, !b[3], a[4], b[4], a[5], !b[5], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2393(w_eco2393, !b[3], a[4], b[4], a[5], !b[5], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2394(w_eco2394, a[3], a[4], b[4], !a[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2395(w_eco2395, a[3], a[4], b[4], !a[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2396(w_eco2396, a[3], !b[3], a[4], b[4], !a[6], !a[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2397(w_eco2397, !b[3], a[4], b[4], !a[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2398(w_eco2398, !b[3], a[4], b[4], !a[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2399(w_eco2399, a[3], !a[4], !b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2400(w_eco2400, a[3], !a[4], !b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2401(w_eco2401, a[3], !a[4], !b[4], b[6], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2402(w_eco2402, a[3], !a[4], !b[4], b[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2403(w_eco2403, a[3], !b[3], !a[4], !b[4], b[6], !a[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2404(w_eco2404, a[3], !b[3], !a[4], !b[4], b[6], !a[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2405(w_eco2405, !b[3], !a[4], !b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2406(w_eco2406, !b[3], !a[4], !b[4], b[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2407(w_eco2407, !b[3], !a[4], !b[4], b[6], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2408(w_eco2408, !b[3], !a[4], !b[4], b[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2409(w_eco2409, a[3], !a[4], !b[4], a[5], !b[5], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2410(w_eco2410, a[3], !a[4], !b[4], a[5], !b[5], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2411(w_eco2411, a[3], !b[3], !a[4], !b[4], a[5], !b[5], !a[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2412(w_eco2412, !b[3], !a[4], !b[4], a[5], !b[5], b[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2413(w_eco2413, !b[3], !a[4], !b[4], a[5], !b[5], !a[1], b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2414(w_eco2414, a[3], !a[4], !b[4], !a[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2415(w_eco2415, a[3], !a[4], !b[4], !a[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2416(w_eco2416, a[3], !b[3], !a[4], !b[4], !a[6], !a[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2417(w_eco2417, !b[3], !a[4], !b[4], !a[6], b[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2418(w_eco2418, !b[3], !a[4], !b[4], !a[6], !a[1], b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2419(w_eco2419, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2420(w_eco2420, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2421(w_eco2421, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_2422(w_eco2422, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_2423(w_eco2423, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_2424(w_eco2424, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2425(w_eco2425, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2426(w_eco2426, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2427(w_eco2427, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2428(w_eco2428, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2429(w_eco2429, !a[3], b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2430(w_eco2430, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2431(w_eco2431, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2432(w_eco2432, !b[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2433(w_eco2433, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2434(w_eco2434, !a[3], !a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2435(w_eco2435, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2436(w_eco2436, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2437(w_eco2437, !a[3], b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2438(w_eco2438, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2439(w_eco2439, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2440(w_eco2440, !b[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2441(w_eco2441, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2442(w_eco2442, !a[3], a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2443(w_eco2443, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2444(w_eco2444, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2445(w_eco2445, a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2446(w_eco2446, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2447(w_eco2447, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2448(w_eco2448, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2449(w_eco2449, !a[3], b[3], !a[4], b[4], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2450(w_eco2450, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2451(w_eco2451, !b[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2452(w_eco2452, !b[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2453(w_eco2453, !a[3], !a[4], b[4], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2454(w_eco2454, !a[3], !a[4], b[4], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2455(w_eco2455, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2456(w_eco2456, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2457(w_eco2457, !a[3], b[3], a[4], !b[4], a[6], b[6], !a[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2458(w_eco2458, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_2459(w_eco2459, !b[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2460(w_eco2460, !b[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_2461(w_eco2461, !a[3], a[4], !b[4], a[6], b[6], !a[1], !a[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2462(w_eco2462, !a[3], a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], a[7], !b[7], !op[1]);
	and _ECO_2463(w_eco2463, a[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2464(w_eco2464, b[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2465(w_eco2465, a[3], !b[3], !a[4], !b[4], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_2466(w_eco2466, b[3], !a[4], !b[4], a[6], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2467(w_eco2467, a[3], a[4], b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2468(w_eco2468, a[3], a[4], b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2469(w_eco2469, !b[3], a[4], b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2470(w_eco2470, !b[3], a[4], b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2471(w_eco2471, a[3], a[4], b[4], a[5], !b[5], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2472(w_eco2472, !b[3], a[4], b[4], a[5], !b[5], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2473(w_eco2473, a[3], a[4], b[4], !a[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2474(w_eco2474, !b[3], a[4], b[4], !a[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2475(w_eco2475, a[3], !a[4], !b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2476(w_eco2476, a[3], !a[4], !b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2477(w_eco2477, !b[3], !a[4], !b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2478(w_eco2478, !b[3], !a[4], !b[4], b[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2479(w_eco2479, a[3], !a[4], !b[4], a[5], !b[5], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2480(w_eco2480, !b[3], !a[4], !b[4], a[5], !b[5], !a[1], a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2481(w_eco2481, a[3], !a[4], !b[4], !a[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2482(w_eco2482, !b[3], !a[4], !b[4], !a[6], !a[1], a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2483(w_eco2483, a[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2484(w_eco2484, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2485(w_eco2485, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_2486(w_eco2486, b[3], a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	or _ECO_2487(w_eco2487, w_eco1835, w_eco1836, w_eco1837, w_eco1838, w_eco1839, w_eco1840, w_eco1841, w_eco1842, w_eco1843, w_eco1844, w_eco1845, w_eco1846, w_eco1847, w_eco1848, w_eco1849, w_eco1850, w_eco1851, w_eco1852, w_eco1853, w_eco1854, w_eco1855, w_eco1856, w_eco1857, w_eco1858, w_eco1859, w_eco1860, w_eco1861, w_eco1862, w_eco1863, w_eco1864, w_eco1865, w_eco1866, w_eco1867, w_eco1868, w_eco1869, w_eco1870, w_eco1871, w_eco1872, w_eco1873, w_eco1874, w_eco1875, w_eco1876, w_eco1877, w_eco1878, w_eco1879, w_eco1880, w_eco1881, w_eco1882, w_eco1883, w_eco1884, w_eco1885, w_eco1886, w_eco1887, w_eco1888, w_eco1889, w_eco1890, w_eco1891, w_eco1892, w_eco1893, w_eco1894, w_eco1895, w_eco1896, w_eco1897, w_eco1898, w_eco1899, w_eco1900, w_eco1901, w_eco1902, w_eco1903, w_eco1904, w_eco1905, w_eco1906, w_eco1907, w_eco1908, w_eco1909, w_eco1910, w_eco1911, w_eco1912, w_eco1913, w_eco1914, w_eco1915, w_eco1916, w_eco1917, w_eco1918, w_eco1919, w_eco1920, w_eco1921, w_eco1922, w_eco1923, w_eco1924, w_eco1925, w_eco1926, w_eco1927, w_eco1928, w_eco1929, w_eco1930, w_eco1931, w_eco1932, w_eco1933, w_eco1934, w_eco1935, w_eco1936, w_eco1937, w_eco1938, w_eco1939, w_eco1940, w_eco1941, w_eco1942, w_eco1943, w_eco1944, w_eco1945, w_eco1946, w_eco1947, w_eco1948, w_eco1949, w_eco1950, w_eco1951, w_eco1952, w_eco1953, w_eco1954, w_eco1955, w_eco1956, w_eco1957, w_eco1958, w_eco1959, w_eco1960, w_eco1961, w_eco1962, w_eco1963, w_eco1964, w_eco1965, w_eco1966, w_eco1967, w_eco1968, w_eco1969, w_eco1970, w_eco1971, w_eco1972, w_eco1973, w_eco1974, w_eco1975, w_eco1976, w_eco1977, w_eco1978, w_eco1979, w_eco1980, w_eco1981, w_eco1982, w_eco1983, w_eco1984, w_eco1985, w_eco1986, w_eco1987, w_eco1988, w_eco1989, w_eco1990, w_eco1991, w_eco1992, w_eco1993, w_eco1994, w_eco1995, w_eco1996, w_eco1997, w_eco1998, w_eco1999, w_eco2000, w_eco2001, w_eco2002, w_eco2003, w_eco2004, w_eco2005, w_eco2006, w_eco2007, w_eco2008, w_eco2009, w_eco2010, w_eco2011, w_eco2012, w_eco2013, w_eco2014, w_eco2015, w_eco2016, w_eco2017, w_eco2018, w_eco2019, w_eco2020, w_eco2021, w_eco2022, w_eco2023, w_eco2024, w_eco2025, w_eco2026, w_eco2027, w_eco2028, w_eco2029, w_eco2030, w_eco2031, w_eco2032, w_eco2033, w_eco2034, w_eco2035, w_eco2036, w_eco2037, w_eco2038, w_eco2039, w_eco2040, w_eco2041, w_eco2042, w_eco2043, w_eco2044, w_eco2045, w_eco2046, w_eco2047, w_eco2048, w_eco2049, w_eco2050, w_eco2051, w_eco2052, w_eco2053, w_eco2054, w_eco2055, w_eco2056, w_eco2057, w_eco2058, w_eco2059, w_eco2060, w_eco2061, w_eco2062, w_eco2063, w_eco2064, w_eco2065, w_eco2066, w_eco2067, w_eco2068, w_eco2069, w_eco2070, w_eco2071, w_eco2072, w_eco2073, w_eco2074, w_eco2075, w_eco2076, w_eco2077, w_eco2078, w_eco2079, w_eco2080, w_eco2081, w_eco2082, w_eco2083, w_eco2084, w_eco2085, w_eco2086, w_eco2087, w_eco2088, w_eco2089, w_eco2090, w_eco2091, w_eco2092, w_eco2093, w_eco2094, w_eco2095, w_eco2096, w_eco2097, w_eco2098, w_eco2099, w_eco2100, w_eco2101, w_eco2102, w_eco2103, w_eco2104, w_eco2105, w_eco2106, w_eco2107, w_eco2108, w_eco2109, w_eco2110, w_eco2111, w_eco2112, w_eco2113, w_eco2114, w_eco2115, w_eco2116, w_eco2117, w_eco2118, w_eco2119, w_eco2120, w_eco2121, w_eco2122, w_eco2123, w_eco2124, w_eco2125, w_eco2126, w_eco2127, w_eco2128, w_eco2129, w_eco2130, w_eco2131, w_eco2132, w_eco2133, w_eco2134, w_eco2135, w_eco2136, w_eco2137, w_eco2138, w_eco2139, w_eco2140, w_eco2141, w_eco2142, w_eco2143, w_eco2144, w_eco2145, w_eco2146, w_eco2147, w_eco2148, w_eco2149, w_eco2150, w_eco2151, w_eco2152, w_eco2153, w_eco2154, w_eco2155, w_eco2156, w_eco2157, w_eco2158, w_eco2159, w_eco2160, w_eco2161, w_eco2162, w_eco2163, w_eco2164, w_eco2165, w_eco2166, w_eco2167, w_eco2168, w_eco2169, w_eco2170, w_eco2171, w_eco2172, w_eco2173, w_eco2174, w_eco2175, w_eco2176, w_eco2177, w_eco2178, w_eco2179, w_eco2180, w_eco2181, w_eco2182, w_eco2183, w_eco2184, w_eco2185, w_eco2186, w_eco2187, w_eco2188, w_eco2189, w_eco2190, w_eco2191, w_eco2192, w_eco2193, w_eco2194, w_eco2195, w_eco2196, w_eco2197, w_eco2198, w_eco2199, w_eco2200, w_eco2201, w_eco2202, w_eco2203, w_eco2204, w_eco2205, w_eco2206, w_eco2207, w_eco2208, w_eco2209, w_eco2210, w_eco2211, w_eco2212, w_eco2213, w_eco2214, w_eco2215, w_eco2216, w_eco2217, w_eco2218, w_eco2219, w_eco2220, w_eco2221, w_eco2222, w_eco2223, w_eco2224, w_eco2225, w_eco2226, w_eco2227, w_eco2228, w_eco2229, w_eco2230, w_eco2231, w_eco2232, w_eco2233, w_eco2234, w_eco2235, w_eco2236, w_eco2237, w_eco2238, w_eco2239, w_eco2240, w_eco2241, w_eco2242, w_eco2243, w_eco2244, w_eco2245, w_eco2246, w_eco2247, w_eco2248, w_eco2249, w_eco2250, w_eco2251, w_eco2252, w_eco2253, w_eco2254, w_eco2255, w_eco2256, w_eco2257, w_eco2258, w_eco2259, w_eco2260, w_eco2261, w_eco2262, w_eco2263, w_eco2264, w_eco2265, w_eco2266, w_eco2267, w_eco2268, w_eco2269, w_eco2270, w_eco2271, w_eco2272, w_eco2273, w_eco2274, w_eco2275, w_eco2276, w_eco2277, w_eco2278, w_eco2279, w_eco2280, w_eco2281, w_eco2282, w_eco2283, w_eco2284, w_eco2285, w_eco2286, w_eco2287, w_eco2288, w_eco2289, w_eco2290, w_eco2291, w_eco2292, w_eco2293, w_eco2294, w_eco2295, w_eco2296, w_eco2297, w_eco2298, w_eco2299, w_eco2300, w_eco2301, w_eco2302, w_eco2303, w_eco2304, w_eco2305, w_eco2306, w_eco2307, w_eco2308, w_eco2309, w_eco2310, w_eco2311, w_eco2312, w_eco2313, w_eco2314, w_eco2315, w_eco2316, w_eco2317, w_eco2318, w_eco2319, w_eco2320, w_eco2321, w_eco2322, w_eco2323, w_eco2324, w_eco2325, w_eco2326, w_eco2327, w_eco2328, w_eco2329, w_eco2330, w_eco2331, w_eco2332, w_eco2333, w_eco2334, w_eco2335, w_eco2336, w_eco2337, w_eco2338, w_eco2339, w_eco2340, w_eco2341, w_eco2342, w_eco2343, w_eco2344, w_eco2345, w_eco2346, w_eco2347, w_eco2348, w_eco2349, w_eco2350, w_eco2351, w_eco2352, w_eco2353, w_eco2354, w_eco2355, w_eco2356, w_eco2357, w_eco2358, w_eco2359, w_eco2360, w_eco2361, w_eco2362, w_eco2363, w_eco2364, w_eco2365, w_eco2366, w_eco2367, w_eco2368, w_eco2369, w_eco2370, w_eco2371, w_eco2372, w_eco2373, w_eco2374, w_eco2375, w_eco2376, w_eco2377, w_eco2378, w_eco2379, w_eco2380, w_eco2381, w_eco2382, w_eco2383, w_eco2384, w_eco2385, w_eco2386, w_eco2387, w_eco2388, w_eco2389, w_eco2390, w_eco2391, w_eco2392, w_eco2393, w_eco2394, w_eco2395, w_eco2396, w_eco2397, w_eco2398, w_eco2399, w_eco2400, w_eco2401, w_eco2402, w_eco2403, w_eco2404, w_eco2405, w_eco2406, w_eco2407, w_eco2408, w_eco2409, w_eco2410, w_eco2411, w_eco2412, w_eco2413, w_eco2414, w_eco2415, w_eco2416, w_eco2417, w_eco2418, w_eco2419, w_eco2420, w_eco2421, w_eco2422, w_eco2423, w_eco2424, w_eco2425, w_eco2426, w_eco2427, w_eco2428, w_eco2429, w_eco2430, w_eco2431, w_eco2432, w_eco2433, w_eco2434, w_eco2435, w_eco2436, w_eco2437, w_eco2438, w_eco2439, w_eco2440, w_eco2441, w_eco2442, w_eco2443, w_eco2444, w_eco2445, w_eco2446, w_eco2447, w_eco2448, w_eco2449, w_eco2450, w_eco2451, w_eco2452, w_eco2453, w_eco2454, w_eco2455, w_eco2456, w_eco2457, w_eco2458, w_eco2459, w_eco2460, w_eco2461, w_eco2462, w_eco2463, w_eco2464, w_eco2465, w_eco2466, w_eco2467, w_eco2468, w_eco2469, w_eco2470, w_eco2471, w_eco2472, w_eco2473, w_eco2474, w_eco2475, w_eco2476, w_eco2477, w_eco2478, w_eco2479, w_eco2480, w_eco2481, w_eco2482, w_eco2483, w_eco2484, w_eco2485, w_eco2486);
	xor _ECO_out5(y[4], sub_wire5, w_eco2487);
	and _ECO_2488(w_eco2488, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2489(w_eco2489, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2490(w_eco2490, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2491(w_eco2491, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2492(w_eco2492, a[3], !b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2493(w_eco2493, !a[3], b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2494(w_eco2494, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2495(w_eco2495, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2496(w_eco2496, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2497(w_eco2497, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2498(w_eco2498, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2499(w_eco2499, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2500(w_eco2500, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2501(w_eco2501, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2502(w_eco2502, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2503(w_eco2503, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2504(w_eco2504, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2505(w_eco2505, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2506(w_eco2506, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2507(w_eco2507, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2508(w_eco2508, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2509(w_eco2509, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2510(w_eco2510, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2511(w_eco2511, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2512(w_eco2512, a[3], b[3], a[4], b[4], a[5], b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2513(w_eco2513, a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2514(w_eco2514, a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2515(w_eco2515, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2516(w_eco2516, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2517(w_eco2517, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2518(w_eco2518, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2519(w_eco2519, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2520(w_eco2520, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2521(w_eco2521, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2522(w_eco2522, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2523(w_eco2523, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2524(w_eco2524, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2525(w_eco2525, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2526(w_eco2526, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2527(w_eco2527, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2528(w_eco2528, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2529(w_eco2529, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2530(w_eco2530, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2531(w_eco2531, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2532(w_eco2532, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2533(w_eco2533, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2534(w_eco2534, a[3], !b[3], !a[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2535(w_eco2535, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2536(w_eco2536, a[3], !b[3], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2537(w_eco2537, a[3], !b[3], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2538(w_eco2538, !a[3], b[3], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2539(w_eco2539, !a[3], b[3], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2540(w_eco2540, a[3], !b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2541(w_eco2541, !a[3], b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2542(w_eco2542, !a[3], !b[3], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2543(w_eco2543, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2544(w_eco2544, !a[3], !b[3], a[5], b[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2545(w_eco2545, a[3], !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2546(w_eco2546, a[3], !b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2547(w_eco2547, a[3], !b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2548(w_eco2548, !a[3], b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2549(w_eco2549, !a[3], b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2550(w_eco2550, !a[3], b[3], a[5], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2551(w_eco2551, a[3], !b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2552(w_eco2552, !a[3], b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2553(w_eco2553, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2554(w_eco2554, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2555(w_eco2555, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2556(w_eco2556, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2557(w_eco2557, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2558(w_eco2558, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2559(w_eco2559, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2560(w_eco2560, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2561(w_eco2561, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2562(w_eco2562, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2563(w_eco2563, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2564(w_eco2564, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2565(w_eco2565, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2566(w_eco2566, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2567(w_eco2567, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2568(w_eco2568, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2569(w_eco2569, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2570(w_eco2570, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2571(w_eco2571, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2572(w_eco2572, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2573(w_eco2573, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2574(w_eco2574, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2575(w_eco2575, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2576(w_eco2576, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2577(w_eco2577, a[3], !b[3], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2578(w_eco2578, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2579(w_eco2579, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2580(w_eco2580, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2581(w_eco2581, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2582(w_eco2582, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2583(w_eco2583, !a[3], !b[3], a[4], b[4], b[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2584(w_eco2584, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2585(w_eco2585, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2586(w_eco2586, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2587(w_eco2587, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2588(w_eco2588, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2589(w_eco2589, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2590(w_eco2590, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2591(w_eco2591, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2592(w_eco2592, a[3], !b[3], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2593(w_eco2593, !a[3], b[3], a[6], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2594(w_eco2594, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2595(w_eco2595, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2596(w_eco2596, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2597(w_eco2597, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2598(w_eco2598, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2599(w_eco2599, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2600(w_eco2600, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2601(w_eco2601, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2602(w_eco2602, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2603(w_eco2603, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2604(w_eco2604, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2605(w_eco2605, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2606(w_eco2606, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2607(w_eco2607, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2608(w_eco2608, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2609(w_eco2609, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2610(w_eco2610, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2611(w_eco2611, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2612(w_eco2612, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2613(w_eco2613, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2614(w_eco2614, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2615(w_eco2615, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2616(w_eco2616, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2617(w_eco2617, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2618(w_eco2618, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2619(w_eco2619, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2620(w_eco2620, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2621(w_eco2621, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2622(w_eco2622, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2623(w_eco2623, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2624(w_eco2624, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2625(w_eco2625, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2626(w_eco2626, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2627(w_eco2627, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2628(w_eco2628, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2629(w_eco2629, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2630(w_eco2630, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2631(w_eco2631, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2632(w_eco2632, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2633(w_eco2633, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2634(w_eco2634, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2635(w_eco2635, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_2636(w_eco2636, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2637(w_eco2637, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2638(w_eco2638, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2639(w_eco2639, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2640(w_eco2640, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2641(w_eco2641, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2642(w_eco2642, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[1], !a[2], op[0], !op[1]);
	and _ECO_2643(w_eco2643, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[2], b[2], op[0], !op[1]);
	and _ECO_2644(w_eco2644, a[3], b[3], a[4], b[4], a[5], b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2645(w_eco2645, a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2646(w_eco2646, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2647(w_eco2647, a[3], !b[3], b[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2648(w_eco2648, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2649(w_eco2649, a[3], !b[3], b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2650(w_eco2650, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2651(w_eco2651, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2652(w_eco2652, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2653(w_eco2653, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2654(w_eco2654, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2655(w_eco2655, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2656(w_eco2656, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2657(w_eco2657, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2658(w_eco2658, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2659(w_eco2659, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2660(w_eco2660, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2661(w_eco2661, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2662(w_eco2662, !a[3], !b[3], a[4], b[4], a[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2663(w_eco2663, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2664(w_eco2664, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2665(w_eco2665, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2666(w_eco2666, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2667(w_eco2667, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2668(w_eco2668, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2669(w_eco2669, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2670(w_eco2670, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2671(w_eco2671, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2672(w_eco2672, a[3], !b[3], b[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2673(w_eco2673, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2674(w_eco2674, a[3], !b[3], b[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2675(w_eco2675, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2676(w_eco2676, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2677(w_eco2677, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2678(w_eco2678, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2679(w_eco2679, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2680(w_eco2680, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2681(w_eco2681, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2682(w_eco2682, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2683(w_eco2683, a[3], !b[3], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2684(w_eco2684, a[3], !b[3], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2685(w_eco2685, a[3], !b[3], !a[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2686(w_eco2686, a[3], !b[3], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2687(w_eco2687, a[3], !b[3], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2688(w_eco2688, !a[3], b[3], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2689(w_eco2689, !a[3], b[3], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2690(w_eco2690, !a[3], b[3], a[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2691(w_eco2691, !a[3], b[3], a[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2692(w_eco2692, a[3], b[3], b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2693(w_eco2693, a[3], b[3], b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2694(w_eco2694, a[3], b[3], !a[1], b[1], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2695(w_eco2695, a[3], b[3], !a[1], b[1], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2696(w_eco2696, a[3], b[3], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2697(w_eco2697, a[3], b[3], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2698(w_eco2698, a[3], !b[3], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2699(w_eco2699, a[3], !b[3], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2700(w_eco2700, !a[3], b[3], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2701(w_eco2701, !a[3], b[3], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2702(w_eco2702, !a[3], !b[3], b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2703(w_eco2703, !a[3], !b[3], b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2704(w_eco2704, !a[3], !b[3], !a[1], b[1], !a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2705(w_eco2705, !a[3], !b[3], !a[1], b[1], !a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2706(w_eco2706, !a[3], !b[3], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2707(w_eco2707, !a[3], !b[3], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2708(w_eco2708, a[3], !b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2709(w_eco2709, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2710(w_eco2710, a[3], !b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2711(w_eco2711, !a[3], b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2712(w_eco2712, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2713(w_eco2713, !a[3], b[3], a[5], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2714(w_eco2714, !a[3], !b[3], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2715(w_eco2715, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2716(w_eco2716, !a[3], !b[3], a[5], b[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2717(w_eco2717, a[3], !b[3], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2718(w_eco2718, a[3], !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2719(w_eco2719, a[3], !b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2720(w_eco2720, !a[3], b[3], a[5], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2721(w_eco2721, !a[3], b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2722(w_eco2722, !a[3], b[3], a[5], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2723(w_eco2723, !a[3], !b[3], a[5], b[5], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2724(w_eco2724, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2725(w_eco2725, a[3], !b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2726(w_eco2726, !a[3], b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2727(w_eco2727, !a[3], !b[3], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2728(w_eco2728, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2729(w_eco2729, !a[3], !b[3], a[5], b[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2730(w_eco2730, a[3], !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2731(w_eco2731, a[3], !b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2732(w_eco2732, a[3], !b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2733(w_eco2733, !a[3], b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2734(w_eco2734, !a[3], b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2735(w_eco2735, !a[3], b[3], a[5], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2736(w_eco2736, a[3], !b[3], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2737(w_eco2737, a[3], !b[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2738(w_eco2738, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2739(w_eco2739, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2740(w_eco2740, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2741(w_eco2741, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2742(w_eco2742, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2743(w_eco2743, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2744(w_eco2744, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2745(w_eco2745, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2746(w_eco2746, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2747(w_eco2747, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2748(w_eco2748, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2749(w_eco2749, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2750(w_eco2750, a[3], b[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2751(w_eco2751, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2752(w_eco2752, a[3], b[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2753(w_eco2753, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2754(w_eco2754, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2755(w_eco2755, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2756(w_eco2756, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2757(w_eco2757, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2758(w_eco2758, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2759(w_eco2759, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2760(w_eco2760, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2761(w_eco2761, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2762(w_eco2762, a[3], !b[3], !a[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2763(w_eco2763, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2764(w_eco2764, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2765(w_eco2765, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2766(w_eco2766, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2767(w_eco2767, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2768(w_eco2768, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2769(w_eco2769, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2770(w_eco2770, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2771(w_eco2771, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2772(w_eco2772, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2773(w_eco2773, a[3], !b[3], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2774(w_eco2774, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2775(w_eco2775, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_2776(w_eco2776, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2777(w_eco2777, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2778(w_eco2778, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2779(w_eco2779, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2780(w_eco2780, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2781(w_eco2781, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2782(w_eco2782, !a[3], !b[3], a[4], b[4], b[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2783(w_eco2783, a[3], !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2784(w_eco2784, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2785(w_eco2785, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2786(w_eco2786, !a[3], b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2787(w_eco2787, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2788(w_eco2788, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2789(w_eco2789, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2790(w_eco2790, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2791(w_eco2791, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2792(w_eco2792, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2793(w_eco2793, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2794(w_eco2794, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2795(w_eco2795, !a[3], !b[3], a[4], b[4], b[5], a[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2796(w_eco2796, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2797(w_eco2797, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2798(w_eco2798, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2799(w_eco2799, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2800(w_eco2800, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2801(w_eco2801, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2802(w_eco2802, a[3], !b[3], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2803(w_eco2803, !a[3], b[3], a[6], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2804(w_eco2804, !a[3], !b[3], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2805(w_eco2805, !a[3], !b[3], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2806(w_eco2806, !a[3], !b[3], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2807(w_eco2807, a[3], !b[3], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2808(w_eco2808, a[3], !b[3], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2809(w_eco2809, a[3], !b[3], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2810(w_eco2810, !a[3], b[3], a[6], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2811(w_eco2811, !a[3], b[3], a[6], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2812(w_eco2812, !a[3], b[3], a[6], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2813(w_eco2813, a[3], !b[3], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2814(w_eco2814, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2815(w_eco2815, a[3], !b[3], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2816(w_eco2816, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2817(w_eco2817, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2818(w_eco2818, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2819(w_eco2819, !a[3], !b[3], a[4], b[4], a[5], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2820(w_eco2820, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2821(w_eco2821, !a[3], !b[3], a[4], b[4], a[5], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2822(w_eco2822, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2823(w_eco2823, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2824(w_eco2824, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2825(w_eco2825, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2826(w_eco2826, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2827(w_eco2827, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2828(w_eco2828, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2829(w_eco2829, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2830(w_eco2830, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2831(w_eco2831, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2832(w_eco2832, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2833(w_eco2833, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2834(w_eco2834, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2835(w_eco2835, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2836(w_eco2836, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2837(w_eco2837, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2838(w_eco2838, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2839(w_eco2839, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2840(w_eco2840, a[3], b[3], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2841(w_eco2841, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !a[7], !op[0], !op[1]);
	and _ECO_2842(w_eco2842, a[3], b[3], !a[5], !b[5], a[6], b[6], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2843(w_eco2843, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2844(w_eco2844, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2845(w_eco2845, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2846(w_eco2846, a[3], !b[3], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2847(w_eco2847, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2848(w_eco2848, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2849(w_eco2849, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2850(w_eco2850, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2851(w_eco2851, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2852(w_eco2852, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2853(w_eco2853, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2854(w_eco2854, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2855(w_eco2855, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2856(w_eco2856, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2857(w_eco2857, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2858(w_eco2858, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2859(w_eco2859, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2860(w_eco2860, a[3], !b[3], !a[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2861(w_eco2861, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2862(w_eco2862, a[3], !b[3], !a[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2863(w_eco2863, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2864(w_eco2864, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2865(w_eco2865, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2866(w_eco2866, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2867(w_eco2867, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2868(w_eco2868, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2869(w_eco2869, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2870(w_eco2870, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2871(w_eco2871, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2872(w_eco2872, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2873(w_eco2873, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2874(w_eco2874, a[3], !b[3], !a[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2875(w_eco2875, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2876(w_eco2876, a[3], !b[3], !a[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_2877(w_eco2877, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], a[0], op[0], !op[1]);
	and _ECO_2878(w_eco2878, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[2], !b[2], op[0], !op[1]);
	and _ECO_2879(w_eco2879, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2880(w_eco2880, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[1], b[2], op[0], !op[1]);
	and _ECO_2881(w_eco2881, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2882(w_eco2882, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2883(w_eco2883, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2884(w_eco2884, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_2885(w_eco2885, a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2886(w_eco2886, a[3], !b[3], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2887(w_eco2887, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2888(w_eco2888, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2889(w_eco2889, a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2890(w_eco2890, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2891(w_eco2891, a[3], !b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2892(w_eco2892, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2893(w_eco2893, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2894(w_eco2894, !a[3], !b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2895(w_eco2895, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2896(w_eco2896, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2897(w_eco2897, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2898(w_eco2898, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2899(w_eco2899, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2900(w_eco2900, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2901(w_eco2901, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2902(w_eco2902, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2903(w_eco2903, !a[3], !b[3], a[4], b[4], a[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2904(w_eco2904, a[3], !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2905(w_eco2905, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2906(w_eco2906, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2907(w_eco2907, !a[3], b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2908(w_eco2908, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2909(w_eco2909, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2910(w_eco2910, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2911(w_eco2911, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2912(w_eco2912, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2913(w_eco2913, a[3], !b[3], b[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2914(w_eco2914, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2915(w_eco2915, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2916(w_eco2916, a[3], b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2917(w_eco2917, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2918(w_eco2918, a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2919(w_eco2919, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2920(w_eco2920, !a[3], b[3], a[4], b[4], a[5], b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2921(w_eco2921, !a[3], !b[3], a[4], b[4], a[5], b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2922(w_eco2922, a[3], b[3], b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2923(w_eco2923, a[3], b[3], b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2924(w_eco2924, a[3], b[3], !a[1], b[1], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2925(w_eco2925, a[3], b[3], !a[1], b[1], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2926(w_eco2926, a[3], !b[3], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2927(w_eco2927, a[3], !b[3], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2928(w_eco2928, a[3], !b[3], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2929(w_eco2929, a[3], !b[3], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2930(w_eco2930, !a[3], b[3], a[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2931(w_eco2931, !a[3], b[3], a[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2932(w_eco2932, !a[3], b[3], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2933(w_eco2933, !a[3], b[3], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2934(w_eco2934, !a[3], !b[3], b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2935(w_eco2935, !a[3], !b[3], b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2936(w_eco2936, !a[3], !b[3], !a[1], b[1], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_2937(w_eco2937, !a[3], !b[3], !a[1], b[1], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_2938(w_eco2938, a[3], !b[3], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2939(w_eco2939, a[3], !b[3], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2940(w_eco2940, a[3], !b[3], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2941(w_eco2941, a[3], !b[3], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2942(w_eco2942, !a[3], b[3], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2943(w_eco2943, !a[3], b[3], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2944(w_eco2944, !a[3], b[3], a[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_2945(w_eco2945, !a[3], b[3], a[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_2946(w_eco2946, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2947(w_eco2947, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2948(w_eco2948, a[3], !b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2949(w_eco2949, a[3], !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2950(w_eco2950, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2951(w_eco2951, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2952(w_eco2952, !a[3], b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_2953(w_eco2953, !a[3], b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2954(w_eco2954, !a[3], !b[3], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2955(w_eco2955, a[3], !b[3], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2956(w_eco2956, a[3], !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2957(w_eco2957, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2958(w_eco2958, !a[3], b[3], a[5], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_2959(w_eco2959, !a[3], b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2960(w_eco2960, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_2961(w_eco2961, !a[3], !b[3], a[5], b[5], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_2962(w_eco2962, !a[3], !b[3], a[5], b[5], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2963(w_eco2963, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_2964(w_eco2964, a[3], !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2965(w_eco2965, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2966(w_eco2966, a[3], !b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2967(w_eco2967, !a[3], b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_2968(w_eco2968, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_2969(w_eco2969, !a[3], b[3], a[5], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_2970(w_eco2970, !a[3], !b[3], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2971(w_eco2971, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2972(w_eco2972, !a[3], !b[3], a[5], b[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2973(w_eco2973, a[3], !b[3], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2974(w_eco2974, a[3], !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2975(w_eco2975, a[3], !b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2976(w_eco2976, !a[3], b[3], a[5], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_2977(w_eco2977, !a[3], b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_2978(w_eco2978, !a[3], b[3], a[5], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_2979(w_eco2979, !a[3], !b[3], a[5], b[5], a[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2980(w_eco2980, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2981(w_eco2981, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2982(w_eco2982, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_2983(w_eco2983, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2984(w_eco2984, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2985(w_eco2985, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2986(w_eco2986, a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2987(w_eco2987, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_2988(w_eco2988, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_2989(w_eco2989, !a[3], !b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_2990(w_eco2990, a[3], b[3], !a[4], !b[4], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2991(w_eco2991, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2992(w_eco2992, a[3], b[3], !a[4], !b[4], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2993(w_eco2993, a[3], b[3], !a[4], !b[4], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2994(w_eco2994, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_2995(w_eco2995, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_2996(w_eco2996, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_2997(w_eco2997, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_2998(w_eco2998, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_2999(w_eco2999, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3000(w_eco3000, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3001(w_eco3001, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_3002(w_eco3002, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3003(w_eco3003, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_3004(w_eco3004, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], b[2], !a[7], !op[1]);
	and _ECO_3005(w_eco3005, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3006(w_eco3006, a[3], !b[3], !a[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3007(w_eco3007, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_3008(w_eco3008, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3009(w_eco3009, a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3010(w_eco3010, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3011(w_eco3011, a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3012(w_eco3012, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3013(w_eco3013, !a[3], b[3], !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3014(w_eco3014, !a[3], !b[3], !a[4], !b[4], a[5], b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3015(w_eco3015, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], a[2], !b[2], !a[0], !a[7], !op[1]);
	and _ECO_3016(w_eco3016, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3017(w_eco3017, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3018(w_eco3018, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3019(w_eco3019, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3020(w_eco3020, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3021(w_eco3021, !a[3], b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3022(w_eco3022, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3023(w_eco3023, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3024(w_eco3024, a[3], !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3025(w_eco3025, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3026(w_eco3026, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3027(w_eco3027, !a[3], b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3028(w_eco3028, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3029(w_eco3029, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3030(w_eco3030, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3031(w_eco3031, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3032(w_eco3032, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3033(w_eco3033, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3034(w_eco3034, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3035(w_eco3035, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3036(w_eco3036, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3037(w_eco3037, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3038(w_eco3038, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3039(w_eco3039, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3040(w_eco3040, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_3041(w_eco3041, !a[3], !b[3], a[4], b[4], b[5], a[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3042(w_eco3042, a[3], !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3043(w_eco3043, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3044(w_eco3044, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3045(w_eco3045, !a[3], b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3046(w_eco3046, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3047(w_eco3047, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3048(w_eco3048, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3049(w_eco3049, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3050(w_eco3050, a[3], !b[3], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3051(w_eco3051, a[3], !b[3], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3052(w_eco3052, a[3], !b[3], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3053(w_eco3053, !a[3], b[3], a[6], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3054(w_eco3054, !a[3], b[3], a[6], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3055(w_eco3055, !a[3], b[3], a[6], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3056(w_eco3056, !a[3], !b[3], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3057(w_eco3057, !a[3], !b[3], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_3058(w_eco3058, !a[3], !b[3], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3059(w_eco3059, a[3], !b[3], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3060(w_eco3060, a[3], !b[3], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3061(w_eco3061, a[3], !b[3], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3062(w_eco3062, !a[3], b[3], a[6], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3063(w_eco3063, !a[3], b[3], a[6], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3064(w_eco3064, !a[3], b[3], a[6], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3065(w_eco3065, !a[3], !b[3], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3066(w_eco3066, !a[3], !b[3], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3067(w_eco3067, a[3], !b[3], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3068(w_eco3068, a[3], !b[3], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3069(w_eco3069, a[3], !b[3], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3070(w_eco3070, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3071(w_eco3071, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3072(w_eco3072, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3073(w_eco3073, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3074(w_eco3074, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3075(w_eco3075, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3076(w_eco3076, !a[3], !b[3], a[4], b[4], a[5], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3077(w_eco3077, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_3078(w_eco3078, !a[3], !b[3], a[4], b[4], a[5], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3079(w_eco3079, a[3], !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3080(w_eco3080, a[3], !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3081(w_eco3081, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3082(w_eco3082, !a[3], b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3083(w_eco3083, !a[3], b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3084(w_eco3084, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3085(w_eco3085, !a[3], !b[3], a[4], b[4], a[5], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3086(w_eco3086, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3087(w_eco3087, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3088(w_eco3088, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_3089(w_eco3089, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3090(w_eco3090, a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3091(w_eco3091, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3092(w_eco3092, a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3093(w_eco3093, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3094(w_eco3094, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3095(w_eco3095, !a[3], !b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3096(w_eco3096, a[3], b[3], !a[5], !b[5], a[6], b[6], b[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3097(w_eco3097, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], !b[7], !op[0], !op[1]);
	and _ECO_3098(w_eco3098, a[3], b[3], !a[5], !b[5], a[6], b[6], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3099(w_eco3099, a[3], b[3], !a[5], !b[5], a[6], b[6], b[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3100(w_eco3100, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], b[1], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3101(w_eco3101, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3102(w_eco3102, a[3], !b[3], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3103(w_eco3103, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_3104(w_eco3104, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3105(w_eco3105, a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3106(w_eco3106, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3107(w_eco3107, a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3108(w_eco3108, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3109(w_eco3109, !a[3], b[3], a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3110(w_eco3110, !a[3], !b[3], a[4], b[4], !a[5], !b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3111(w_eco3111, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3112(w_eco3112, a[3], !b[3], !a[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3113(w_eco3113, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_3114(w_eco3114, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3115(w_eco3115, a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3116(w_eco3116, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3117(w_eco3117, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3118(w_eco3118, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3119(w_eco3119, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3120(w_eco3120, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3121(w_eco3121, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3122(w_eco3122, a[3], !b[3], !a[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3123(w_eco3123, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], op[0], !op[1]);
	and _ECO_3124(w_eco3124, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3125(w_eco3125, a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3126(w_eco3126, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3127(w_eco3127, a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3128(w_eco3128, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_3129(w_eco3129, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[1], !b[2], op[0], !op[1]);
	and _ECO_3130(w_eco3130, !a[3], !b[3], !a[4], !b[4], !a[5], !b[5], !b[6], !a[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3131(w_eco3131, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3132(w_eco3132, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3133(w_eco3133, a[3], !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3134(w_eco3134, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3135(w_eco3135, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3136(w_eco3136, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3137(w_eco3137, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3138(w_eco3138, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3139(w_eco3139, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3140(w_eco3140, a[3], !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3141(w_eco3141, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3142(w_eco3142, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3143(w_eco3143, !a[3], b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3144(w_eco3144, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3145(w_eco3145, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3146(w_eco3146, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3147(w_eco3147, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3148(w_eco3148, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3149(w_eco3149, a[3], b[3], !a[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3150(w_eco3150, a[3], b[3], !a[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3151(w_eco3151, !a[3], b[3], a[1], !b[1], a[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3152(w_eco3152, !a[3], b[3], a[1], !b[1], a[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3153(w_eco3153, !a[3], !b[3], !a[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3154(w_eco3154, !a[3], !b[3], !a[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3155(w_eco3155, a[3], b[3], !a[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3156(w_eco3156, a[3], b[3], !a[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3157(w_eco3157, a[3], !b[3], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3158(w_eco3158, a[3], !b[3], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3159(w_eco3159, a[3], !b[3], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3160(w_eco3160, a[3], !b[3], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3161(w_eco3161, !a[3], b[3], a[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3162(w_eco3162, !a[3], b[3], a[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3163(w_eco3163, !a[3], b[3], a[1], !b[1], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3164(w_eco3164, !a[3], b[3], a[1], !b[1], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3165(w_eco3165, !a[3], !b[3], !a[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3166(w_eco3166, !a[3], !b[3], !a[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3167(w_eco3167, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3168(w_eco3168, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3169(w_eco3169, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3170(w_eco3170, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3171(w_eco3171, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3172(w_eco3172, a[3], !b[3], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3173(w_eco3173, a[3], !b[3], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3174(w_eco3174, a[3], !b[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3175(w_eco3175, a[3], !b[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3176(w_eco3176, !a[3], b[3], a[6], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3177(w_eco3177, !a[3], b[3], a[6], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3178(w_eco3178, !a[3], b[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3179(w_eco3179, !a[3], b[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3180(w_eco3180, !a[3], !b[3], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3181(w_eco3181, a[3], b[3], !a[5], !b[5], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3182(w_eco3182, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3183(w_eco3183, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3184(w_eco3184, a[3], !b[3], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3185(w_eco3185, a[3], !b[3], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3186(w_eco3186, a[3], !b[3], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3187(w_eco3187, !a[3], b[3], a[6], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3188(w_eco3188, !a[3], b[3], a[6], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3189(w_eco3189, !a[3], b[3], a[6], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3190(w_eco3190, !a[3], !b[3], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3191(w_eco3191, !a[3], !b[3], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3192(w_eco3192, !a[3], !b[3], a[6], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3193(w_eco3193, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3194(w_eco3194, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3195(w_eco3195, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3196(w_eco3196, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3197(w_eco3197, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3198(w_eco3198, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3199(w_eco3199, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3200(w_eco3200, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3201(w_eco3201, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3202(w_eco3202, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3203(w_eco3203, a[3], !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3204(w_eco3204, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3205(w_eco3205, !a[3], b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3206(w_eco3206, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3207(w_eco3207, !a[3], !b[3], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3208(w_eco3208, a[3], !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3209(w_eco3209, a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3210(w_eco3210, !a[3], b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3211(w_eco3211, !a[3], b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3212(w_eco3212, !a[3], !b[3], a[5], b[5], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3213(w_eco3213, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3214(w_eco3214, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3215(w_eco3215, a[3], !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3216(w_eco3216, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3217(w_eco3217, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3218(w_eco3218, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3219(w_eco3219, !a[3], b[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3220(w_eco3220, !a[3], b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3221(w_eco3221, !a[3], !b[3], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3222(w_eco3222, a[3], !b[3], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3223(w_eco3223, a[3], !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3224(w_eco3224, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3225(w_eco3225, !a[3], b[3], a[5], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3226(w_eco3226, !a[3], b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3227(w_eco3227, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3228(w_eco3228, !a[3], !b[3], a[5], b[5], a[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3229(w_eco3229, !a[3], !b[3], a[5], b[5], a[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3230(w_eco3230, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3231(w_eco3231, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3232(w_eco3232, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3233(w_eco3233, !a[3], b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3234(w_eco3234, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3235(w_eco3235, !a[3], !b[3], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3236(w_eco3236, a[3], !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3237(w_eco3237, a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3238(w_eco3238, !a[3], b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3239(w_eco3239, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3240(w_eco3240, !a[3], !b[3], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3241(w_eco3241, a[3], !b[3], b[6], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3242(w_eco3242, a[3], !b[3], a[4], !b[4], a[5], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3243(w_eco3243, a[3], !b[3], !a[6], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3244(w_eco3244, a[3], !b[3], a[5], !b[5], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3245(w_eco3245, a[3], !b[3], a[4], !b[4], !b[5], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3246(w_eco3246, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3247(w_eco3247, a[3], !b[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3248(w_eco3248, a[3], !b[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3249(w_eco3249, !a[3], b[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3250(w_eco3250, !a[3], b[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3251(w_eco3251, !a[3], !b[3], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3252(w_eco3252, a[3], b[3], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3253(w_eco3253, a[3], !b[3], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3254(w_eco3254, a[3], !b[3], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3255(w_eco3255, !a[3], b[3], a[6], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3256(w_eco3256, !a[3], b[3], a[6], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3257(w_eco3257, !a[3], !b[3], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3258(w_eco3258, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3259(w_eco3259, a[3], b[3], !a[4], !b[4], a[5], b[5], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3260(w_eco3260, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3261(w_eco3261, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_3262(w_eco3262, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], b[0], !a[7], !op[1]);
	and _ECO_3263(w_eco3263, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], b[2], !b[7], !op[1]);
	and _ECO_3264(w_eco3264, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3265(w_eco3265, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3266(w_eco3266, a[3], !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3267(w_eco3267, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3268(w_eco3268, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3269(w_eco3269, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3270(w_eco3270, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3271(w_eco3271, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3272(w_eco3272, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3273(w_eco3273, a[3], !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3274(w_eco3274, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3275(w_eco3275, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3276(w_eco3276, !a[3], b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3277(w_eco3277, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3278(w_eco3278, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3279(w_eco3279, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3280(w_eco3280, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3281(w_eco3281, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3282(w_eco3282, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3283(w_eco3283, a[3], b[3], !a[4], !b[4], a[6], b[6], b[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3284(w_eco3284, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3285(w_eco3285, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3286(w_eco3286, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3287(w_eco3287, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3288(w_eco3288, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3289(w_eco3289, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3290(w_eco3290, a[3], !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3291(w_eco3291, !a[3], b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3292(w_eco3292, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3293(w_eco3293, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], b[2], a[7], !b[7], !op[1]);
	and _ECO_3294(w_eco3294, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3295(w_eco3295, a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], b[0], !b[7], !op[1]);
	and _ECO_3296(w_eco3296, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3297(w_eco3297, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3298(w_eco3298, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3299(w_eco3299, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3300(w_eco3300, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3301(w_eco3301, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3302(w_eco3302, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3303(w_eco3303, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3304(w_eco3304, !a[3], b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3305(w_eco3305, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3306(w_eco3306, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3307(w_eco3307, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3308(w_eco3308, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3309(w_eco3309, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3310(w_eco3310, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3311(w_eco3311, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3312(w_eco3312, a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3313(w_eco3313, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3314(w_eco3314, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3315(w_eco3315, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3316(w_eco3316, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3317(w_eco3317, a[3], b[3], !a[4], !b[4], a[6], b[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3318(w_eco3318, a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3319(w_eco3319, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3320(w_eco3320, !a[3], b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3321(w_eco3321, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3322(w_eco3322, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3323(w_eco3323, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3324(w_eco3324, a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3325(w_eco3325, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3326(w_eco3326, !a[3], b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], !a[7], !op[0], !op[1]);
	and _ECO_3327(w_eco3327, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_3328(w_eco3328, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3329(w_eco3329, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3330(w_eco3330, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !a[0], a[7], !b[7], !op[1]);
	and _ECO_3331(w_eco3331, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3332(w_eco3332, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3333(w_eco3333, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3334(w_eco3334, a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3335(w_eco3335, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3336(w_eco3336, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], !b[7], !op[0], !op[1]);
	and _ECO_3337(w_eco3337, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], b[2], a[0], b[0], a[7], !b[7], !op[1]);
	or _ECO_3338(w_eco3338, w_eco2488, w_eco2489, w_eco2490, w_eco2491, w_eco2492, w_eco2493, w_eco2494, w_eco2495, w_eco2496, w_eco2497, w_eco2498, w_eco2499, w_eco2500, w_eco2501, w_eco2502, w_eco2503, w_eco2504, w_eco2505, w_eco2506, w_eco2507, w_eco2508, w_eco2509, w_eco2510, w_eco2511, w_eco2512, w_eco2513, w_eco2514, w_eco2515, w_eco2516, w_eco2517, w_eco2518, w_eco2519, w_eco2520, w_eco2521, w_eco2522, w_eco2523, w_eco2524, w_eco2525, w_eco2526, w_eco2527, w_eco2528, w_eco2529, w_eco2530, w_eco2531, w_eco2532, w_eco2533, w_eco2534, w_eco2535, w_eco2536, w_eco2537, w_eco2538, w_eco2539, w_eco2540, w_eco2541, w_eco2542, w_eco2543, w_eco2544, w_eco2545, w_eco2546, w_eco2547, w_eco2548, w_eco2549, w_eco2550, w_eco2551, w_eco2552, w_eco2553, w_eco2554, w_eco2555, w_eco2556, w_eco2557, w_eco2558, w_eco2559, w_eco2560, w_eco2561, w_eco2562, w_eco2563, w_eco2564, w_eco2565, w_eco2566, w_eco2567, w_eco2568, w_eco2569, w_eco2570, w_eco2571, w_eco2572, w_eco2573, w_eco2574, w_eco2575, w_eco2576, w_eco2577, w_eco2578, w_eco2579, w_eco2580, w_eco2581, w_eco2582, w_eco2583, w_eco2584, w_eco2585, w_eco2586, w_eco2587, w_eco2588, w_eco2589, w_eco2590, w_eco2591, w_eco2592, w_eco2593, w_eco2594, w_eco2595, w_eco2596, w_eco2597, w_eco2598, w_eco2599, w_eco2600, w_eco2601, w_eco2602, w_eco2603, w_eco2604, w_eco2605, w_eco2606, w_eco2607, w_eco2608, w_eco2609, w_eco2610, w_eco2611, w_eco2612, w_eco2613, w_eco2614, w_eco2615, w_eco2616, w_eco2617, w_eco2618, w_eco2619, w_eco2620, w_eco2621, w_eco2622, w_eco2623, w_eco2624, w_eco2625, w_eco2626, w_eco2627, w_eco2628, w_eco2629, w_eco2630, w_eco2631, w_eco2632, w_eco2633, w_eco2634, w_eco2635, w_eco2636, w_eco2637, w_eco2638, w_eco2639, w_eco2640, w_eco2641, w_eco2642, w_eco2643, w_eco2644, w_eco2645, w_eco2646, w_eco2647, w_eco2648, w_eco2649, w_eco2650, w_eco2651, w_eco2652, w_eco2653, w_eco2654, w_eco2655, w_eco2656, w_eco2657, w_eco2658, w_eco2659, w_eco2660, w_eco2661, w_eco2662, w_eco2663, w_eco2664, w_eco2665, w_eco2666, w_eco2667, w_eco2668, w_eco2669, w_eco2670, w_eco2671, w_eco2672, w_eco2673, w_eco2674, w_eco2675, w_eco2676, w_eco2677, w_eco2678, w_eco2679, w_eco2680, w_eco2681, w_eco2682, w_eco2683, w_eco2684, w_eco2685, w_eco2686, w_eco2687, w_eco2688, w_eco2689, w_eco2690, w_eco2691, w_eco2692, w_eco2693, w_eco2694, w_eco2695, w_eco2696, w_eco2697, w_eco2698, w_eco2699, w_eco2700, w_eco2701, w_eco2702, w_eco2703, w_eco2704, w_eco2705, w_eco2706, w_eco2707, w_eco2708, w_eco2709, w_eco2710, w_eco2711, w_eco2712, w_eco2713, w_eco2714, w_eco2715, w_eco2716, w_eco2717, w_eco2718, w_eco2719, w_eco2720, w_eco2721, w_eco2722, w_eco2723, w_eco2724, w_eco2725, w_eco2726, w_eco2727, w_eco2728, w_eco2729, w_eco2730, w_eco2731, w_eco2732, w_eco2733, w_eco2734, w_eco2735, w_eco2736, w_eco2737, w_eco2738, w_eco2739, w_eco2740, w_eco2741, w_eco2742, w_eco2743, w_eco2744, w_eco2745, w_eco2746, w_eco2747, w_eco2748, w_eco2749, w_eco2750, w_eco2751, w_eco2752, w_eco2753, w_eco2754, w_eco2755, w_eco2756, w_eco2757, w_eco2758, w_eco2759, w_eco2760, w_eco2761, w_eco2762, w_eco2763, w_eco2764, w_eco2765, w_eco2766, w_eco2767, w_eco2768, w_eco2769, w_eco2770, w_eco2771, w_eco2772, w_eco2773, w_eco2774, w_eco2775, w_eco2776, w_eco2777, w_eco2778, w_eco2779, w_eco2780, w_eco2781, w_eco2782, w_eco2783, w_eco2784, w_eco2785, w_eco2786, w_eco2787, w_eco2788, w_eco2789, w_eco2790, w_eco2791, w_eco2792, w_eco2793, w_eco2794, w_eco2795, w_eco2796, w_eco2797, w_eco2798, w_eco2799, w_eco2800, w_eco2801, w_eco2802, w_eco2803, w_eco2804, w_eco2805, w_eco2806, w_eco2807, w_eco2808, w_eco2809, w_eco2810, w_eco2811, w_eco2812, w_eco2813, w_eco2814, w_eco2815, w_eco2816, w_eco2817, w_eco2818, w_eco2819, w_eco2820, w_eco2821, w_eco2822, w_eco2823, w_eco2824, w_eco2825, w_eco2826, w_eco2827, w_eco2828, w_eco2829, w_eco2830, w_eco2831, w_eco2832, w_eco2833, w_eco2834, w_eco2835, w_eco2836, w_eco2837, w_eco2838, w_eco2839, w_eco2840, w_eco2841, w_eco2842, w_eco2843, w_eco2844, w_eco2845, w_eco2846, w_eco2847, w_eco2848, w_eco2849, w_eco2850, w_eco2851, w_eco2852, w_eco2853, w_eco2854, w_eco2855, w_eco2856, w_eco2857, w_eco2858, w_eco2859, w_eco2860, w_eco2861, w_eco2862, w_eco2863, w_eco2864, w_eco2865, w_eco2866, w_eco2867, w_eco2868, w_eco2869, w_eco2870, w_eco2871, w_eco2872, w_eco2873, w_eco2874, w_eco2875, w_eco2876, w_eco2877, w_eco2878, w_eco2879, w_eco2880, w_eco2881, w_eco2882, w_eco2883, w_eco2884, w_eco2885, w_eco2886, w_eco2887, w_eco2888, w_eco2889, w_eco2890, w_eco2891, w_eco2892, w_eco2893, w_eco2894, w_eco2895, w_eco2896, w_eco2897, w_eco2898, w_eco2899, w_eco2900, w_eco2901, w_eco2902, w_eco2903, w_eco2904, w_eco2905, w_eco2906, w_eco2907, w_eco2908, w_eco2909, w_eco2910, w_eco2911, w_eco2912, w_eco2913, w_eco2914, w_eco2915, w_eco2916, w_eco2917, w_eco2918, w_eco2919, w_eco2920, w_eco2921, w_eco2922, w_eco2923, w_eco2924, w_eco2925, w_eco2926, w_eco2927, w_eco2928, w_eco2929, w_eco2930, w_eco2931, w_eco2932, w_eco2933, w_eco2934, w_eco2935, w_eco2936, w_eco2937, w_eco2938, w_eco2939, w_eco2940, w_eco2941, w_eco2942, w_eco2943, w_eco2944, w_eco2945, w_eco2946, w_eco2947, w_eco2948, w_eco2949, w_eco2950, w_eco2951, w_eco2952, w_eco2953, w_eco2954, w_eco2955, w_eco2956, w_eco2957, w_eco2958, w_eco2959, w_eco2960, w_eco2961, w_eco2962, w_eco2963, w_eco2964, w_eco2965, w_eco2966, w_eco2967, w_eco2968, w_eco2969, w_eco2970, w_eco2971, w_eco2972, w_eco2973, w_eco2974, w_eco2975, w_eco2976, w_eco2977, w_eco2978, w_eco2979, w_eco2980, w_eco2981, w_eco2982, w_eco2983, w_eco2984, w_eco2985, w_eco2986, w_eco2987, w_eco2988, w_eco2989, w_eco2990, w_eco2991, w_eco2992, w_eco2993, w_eco2994, w_eco2995, w_eco2996, w_eco2997, w_eco2998, w_eco2999, w_eco3000, w_eco3001, w_eco3002, w_eco3003, w_eco3004, w_eco3005, w_eco3006, w_eco3007, w_eco3008, w_eco3009, w_eco3010, w_eco3011, w_eco3012, w_eco3013, w_eco3014, w_eco3015, w_eco3016, w_eco3017, w_eco3018, w_eco3019, w_eco3020, w_eco3021, w_eco3022, w_eco3023, w_eco3024, w_eco3025, w_eco3026, w_eco3027, w_eco3028, w_eco3029, w_eco3030, w_eco3031, w_eco3032, w_eco3033, w_eco3034, w_eco3035, w_eco3036, w_eco3037, w_eco3038, w_eco3039, w_eco3040, w_eco3041, w_eco3042, w_eco3043, w_eco3044, w_eco3045, w_eco3046, w_eco3047, w_eco3048, w_eco3049, w_eco3050, w_eco3051, w_eco3052, w_eco3053, w_eco3054, w_eco3055, w_eco3056, w_eco3057, w_eco3058, w_eco3059, w_eco3060, w_eco3061, w_eco3062, w_eco3063, w_eco3064, w_eco3065, w_eco3066, w_eco3067, w_eco3068, w_eco3069, w_eco3070, w_eco3071, w_eco3072, w_eco3073, w_eco3074, w_eco3075, w_eco3076, w_eco3077, w_eco3078, w_eco3079, w_eco3080, w_eco3081, w_eco3082, w_eco3083, w_eco3084, w_eco3085, w_eco3086, w_eco3087, w_eco3088, w_eco3089, w_eco3090, w_eco3091, w_eco3092, w_eco3093, w_eco3094, w_eco3095, w_eco3096, w_eco3097, w_eco3098, w_eco3099, w_eco3100, w_eco3101, w_eco3102, w_eco3103, w_eco3104, w_eco3105, w_eco3106, w_eco3107, w_eco3108, w_eco3109, w_eco3110, w_eco3111, w_eco3112, w_eco3113, w_eco3114, w_eco3115, w_eco3116, w_eco3117, w_eco3118, w_eco3119, w_eco3120, w_eco3121, w_eco3122, w_eco3123, w_eco3124, w_eco3125, w_eco3126, w_eco3127, w_eco3128, w_eco3129, w_eco3130, w_eco3131, w_eco3132, w_eco3133, w_eco3134, w_eco3135, w_eco3136, w_eco3137, w_eco3138, w_eco3139, w_eco3140, w_eco3141, w_eco3142, w_eco3143, w_eco3144, w_eco3145, w_eco3146, w_eco3147, w_eco3148, w_eco3149, w_eco3150, w_eco3151, w_eco3152, w_eco3153, w_eco3154, w_eco3155, w_eco3156, w_eco3157, w_eco3158, w_eco3159, w_eco3160, w_eco3161, w_eco3162, w_eco3163, w_eco3164, w_eco3165, w_eco3166, w_eco3167, w_eco3168, w_eco3169, w_eco3170, w_eco3171, w_eco3172, w_eco3173, w_eco3174, w_eco3175, w_eco3176, w_eco3177, w_eco3178, w_eco3179, w_eco3180, w_eco3181, w_eco3182, w_eco3183, w_eco3184, w_eco3185, w_eco3186, w_eco3187, w_eco3188, w_eco3189, w_eco3190, w_eco3191, w_eco3192, w_eco3193, w_eco3194, w_eco3195, w_eco3196, w_eco3197, w_eco3198, w_eco3199, w_eco3200, w_eco3201, w_eco3202, w_eco3203, w_eco3204, w_eco3205, w_eco3206, w_eco3207, w_eco3208, w_eco3209, w_eco3210, w_eco3211, w_eco3212, w_eco3213, w_eco3214, w_eco3215, w_eco3216, w_eco3217, w_eco3218, w_eco3219, w_eco3220, w_eco3221, w_eco3222, w_eco3223, w_eco3224, w_eco3225, w_eco3226, w_eco3227, w_eco3228, w_eco3229, w_eco3230, w_eco3231, w_eco3232, w_eco3233, w_eco3234, w_eco3235, w_eco3236, w_eco3237, w_eco3238, w_eco3239, w_eco3240, w_eco3241, w_eco3242, w_eco3243, w_eco3244, w_eco3245, w_eco3246, w_eco3247, w_eco3248, w_eco3249, w_eco3250, w_eco3251, w_eco3252, w_eco3253, w_eco3254, w_eco3255, w_eco3256, w_eco3257, w_eco3258, w_eco3259, w_eco3260, w_eco3261, w_eco3262, w_eco3263, w_eco3264, w_eco3265, w_eco3266, w_eco3267, w_eco3268, w_eco3269, w_eco3270, w_eco3271, w_eco3272, w_eco3273, w_eco3274, w_eco3275, w_eco3276, w_eco3277, w_eco3278, w_eco3279, w_eco3280, w_eco3281, w_eco3282, w_eco3283, w_eco3284, w_eco3285, w_eco3286, w_eco3287, w_eco3288, w_eco3289, w_eco3290, w_eco3291, w_eco3292, w_eco3293, w_eco3294, w_eco3295, w_eco3296, w_eco3297, w_eco3298, w_eco3299, w_eco3300, w_eco3301, w_eco3302, w_eco3303, w_eco3304, w_eco3305, w_eco3306, w_eco3307, w_eco3308, w_eco3309, w_eco3310, w_eco3311, w_eco3312, w_eco3313, w_eco3314, w_eco3315, w_eco3316, w_eco3317, w_eco3318, w_eco3319, w_eco3320, w_eco3321, w_eco3322, w_eco3323, w_eco3324, w_eco3325, w_eco3326, w_eco3327, w_eco3328, w_eco3329, w_eco3330, w_eco3331, w_eco3332, w_eco3333, w_eco3334, w_eco3335, w_eco3336, w_eco3337);
	xor _ECO_out6(y[3], sub_wire6, w_eco3338);
	and _ECO_3339(w_eco3339, a[4], b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3340(w_eco3340, a[4], b[4], a[5], b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3341(w_eco3341, a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3342(w_eco3342, a[4], b[4], a[5], b[5], !a[6], !b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3343(w_eco3343, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3344(w_eco3344, !a[4], !b[4], a[5], b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3345(w_eco3345, !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3346(w_eco3346, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3347(w_eco3347, a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3348(w_eco3348, a[4], b[4], !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3349(w_eco3349, a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3350(w_eco3350, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3351(w_eco3351, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3352(w_eco3352, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3353(w_eco3353, !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3354(w_eco3354, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3355(w_eco3355, a[4], b[4], a[5], b[5], a[6], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3356(w_eco3356, a[4], b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3357(w_eco3357, a[4], b[4], a[5], b[5], a[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3358(w_eco3358, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3359(w_eco3359, a[4], b[4], a[5], b[5], a[6], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3360(w_eco3360, a[4], b[4], a[5], b[5], a[6], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3361(w_eco3361, a[4], b[4], a[5], b[5], a[6], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3362(w_eco3362, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3363(w_eco3363, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3364(w_eco3364, a[4], b[4], a[5], b[5], !a[6], !b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3365(w_eco3365, a[4], b[4], a[5], b[5], !b[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3366(w_eco3366, a[4], b[4], a[5], b[5], !b[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3367(w_eco3367, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3368(w_eco3368, a[4], b[4], a[5], b[5], !a[6], !b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3369(w_eco3369, a[4], b[4], a[5], b[5], !a[6], !b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3370(w_eco3370, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3371(w_eco3371, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3372(w_eco3372, a[3], !b[3], !a[4], b[5], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3373(w_eco3373, !a[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3374(w_eco3374, !a[4], !b[4], a[5], b[5], a[6], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3375(w_eco3375, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3376(w_eco3376, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3377(w_eco3377, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3378(w_eco3378, !a[4], !b[4], a[5], b[5], a[6], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3379(w_eco3379, !a[4], !b[4], a[5], b[5], a[6], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3380(w_eco3380, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3381(w_eco3381, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3382(w_eco3382, !a[4], !b[4], a[6], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3383(w_eco3383, !a[4], !b[4], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3384(w_eco3384, !a[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3385(w_eco3385, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_3386(w_eco3386, !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3387(w_eco3387, !a[4], !b[4], a[5], b[5], !a[6], !b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3388(w_eco3388, !a[4], !b[4], a[5], b[5], !b[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3389(w_eco3389, !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3390(w_eco3390, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3391(w_eco3391, !a[4], !b[4], a[5], b[5], !a[6], !b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3392(w_eco3392, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3393(w_eco3393, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3394(w_eco3394, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3395(w_eco3395, a[3], !b[3], b[4], !a[5], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3396(w_eco3396, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3397(w_eco3397, !a[4], !b[4], a[6], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3398(w_eco3398, a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3399(w_eco3399, a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3400(w_eco3400, a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3401(w_eco3401, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3402(w_eco3402, a[4], b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3403(w_eco3403, a[4], b[4], !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3404(w_eco3404, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3405(w_eco3405, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3406(w_eco3406, !a[5], !b[5], a[6], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3407(w_eco3407, !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3408(w_eco3408, !a[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3409(w_eco3409, a[4], b[4], !a[5], !b[5], !a[6], !b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3410(w_eco3410, a[4], b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3411(w_eco3411, a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3412(w_eco3412, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3413(w_eco3413, a[4], b[4], !a[5], !b[5], !a[6], !b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3414(w_eco3414, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3415(w_eco3415, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3416(w_eco3416, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3417(w_eco3417, !a[4], !b[4], !a[5], !b[5], a[6], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3418(w_eco3418, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3419(w_eco3419, !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3420(w_eco3420, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3421(w_eco3421, !a[4], !b[4], !a[5], !b[5], a[6], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3422(w_eco3422, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3423(w_eco3423, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3424(w_eco3424, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3425(w_eco3425, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3426(w_eco3426, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3427(w_eco3427, !a[4], !b[4], !a[5], !b[5], !b[6], !b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3428(w_eco3428, !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_3429(w_eco3429, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3430(w_eco3430, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3431(w_eco3431, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3432(w_eco3432, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3433(w_eco3433, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3434(w_eco3434, a[4], b[4], a[5], b[5], a[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3435(w_eco3435, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3436(w_eco3436, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3437(w_eco3437, a[4], b[4], a[5], b[5], a[6], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3438(w_eco3438, a[4], b[4], a[5], b[5], a[6], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3439(w_eco3439, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3440(w_eco3440, a[3], !b[3], !a[6], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3441(w_eco3441, !a[3], a[4], b[4], a[5], b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3442(w_eco3442, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3443(w_eco3443, b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3444(w_eco3444, !a[3], a[4], b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3445(w_eco3445, !a[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3446(w_eco3446, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3447(w_eco3447, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3448(w_eco3448, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3449(w_eco3449, a[4], b[4], a[5], b[5], !b[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3450(w_eco3450, a[4], b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3451(w_eco3451, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3452(w_eco3452, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3453(w_eco3453, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3454(w_eco3454, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3455(w_eco3455, a[3], !b[3], !a[4], b[5], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3456(w_eco3456, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3457(w_eco3457, !b[1], a[2], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3458(w_eco3458, !b[1], a[2], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3459(w_eco3459, a[3], !b[3], !a[4], b[5], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3460(w_eco3460, a[3], !b[3], !a[4], b[5], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3461(w_eco3461, a[3], !b[3], !a[4], b[5], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3462(w_eco3462, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3463(w_eco3463, !a[3], !b[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3464(w_eco3464, !a[3], !b[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3465(w_eco3465, !b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3466(w_eco3466, !a[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3467(w_eco3467, !b[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3468(w_eco3468, !a[3], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3469(w_eco3469, !a[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3470(w_eco3470, !a[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3471(w_eco3471, !a[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3472(w_eco3472, !a[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3473(w_eco3473, !a[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3474(w_eco3474, a[3], !b[3], !a[4], b[5], !a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3475(w_eco3475, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3476(w_eco3476, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3477(w_eco3477, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3478(w_eco3478, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3479(w_eco3479, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3480(w_eco3480, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3481(w_eco3481, !a[4], !b[4], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3482(w_eco3482, !a[4], !b[4], a[6], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3483(w_eco3483, !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3484(w_eco3484, !a[4], !b[4], a[6], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3485(w_eco3485, !a[4], !b[4], a[6], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3486(w_eco3486, !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3487(w_eco3487, !a[4], !b[4], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3488(w_eco3488, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3489(w_eco3489, !a[4], !b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3490(w_eco3490, !a[4], !b[4], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3491(w_eco3491, !a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3492(w_eco3492, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3493(w_eco3493, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3494(w_eco3494, !a[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3495(w_eco3495, !a[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3496(w_eco3496, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3497(w_eco3497, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3498(w_eco3498, !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3499(w_eco3499, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3500(w_eco3500, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3501(w_eco3501, !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3502(w_eco3502, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], !b[7], !op[1]);
	and _ECO_3503(w_eco3503, !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3504(w_eco3504, !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3505(w_eco3505, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3506(w_eco3506, !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3507(w_eco3507, !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3508(w_eco3508, !a[4], !b[4], a[5], b[5], !b[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3509(w_eco3509, !a[4], !b[4], a[5], b[5], !b[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3510(w_eco3510, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3511(w_eco3511, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3512(w_eco3512, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3513(w_eco3513, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3514(w_eco3514, a[3], !b[3], b[4], !a[5], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3515(w_eco3515, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3516(w_eco3516, a[3], !b[3], b[4], !a[5], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3517(w_eco3517, a[3], !b[3], b[4], !a[5], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3518(w_eco3518, a[3], !b[3], b[4], !a[5], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3519(w_eco3519, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3520(w_eco3520, !b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3521(w_eco3521, !a[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3522(w_eco3522, a[3], !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[1]);
	and _ECO_3523(w_eco3523, !a[3], a[4], b[4], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3524(w_eco3524, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3525(w_eco3525, !a[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3526(w_eco3526, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3527(w_eco3527, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3528(w_eco3528, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3529(w_eco3529, a[3], !b[3], b[4], !a[5], !a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3530(w_eco3530, !a[3], a[6], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3531(w_eco3531, a[3], !b[3], !a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3532(w_eco3532, a[3], !b[3], !a[5], b[5], !a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3533(w_eco3533, !a[4], !b[4], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3534(w_eco3534, !a[4], !b[4], a[6], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3535(w_eco3535, !a[4], !b[4], a[6], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3536(w_eco3536, !a[4], !b[4], a[6], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3537(w_eco3537, !a[4], !b[4], a[6], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3538(w_eco3538, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3539(w_eco3539, a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3540(w_eco3540, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3541(w_eco3541, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3542(w_eco3542, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3543(w_eco3543, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3544(w_eco3544, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3545(w_eco3545, !a[5], !b[5], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3546(w_eco3546, !a[5], !b[5], a[6], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3547(w_eco3547, !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3548(w_eco3548, !a[5], !b[5], a[6], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3549(w_eco3549, !a[5], !b[5], a[6], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3550(w_eco3550, !a[5], !b[5], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3551(w_eco3551, !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3552(w_eco3552, !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3553(w_eco3553, !a[5], !b[5], a[6], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3554(w_eco3554, !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3555(w_eco3555, !a[3], a[4], b[4], !a[5], !b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3556(w_eco3556, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3557(w_eco3557, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3558(w_eco3558, !a[3], a[4], b[4], !a[5], !b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3559(w_eco3559, !a[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3560(w_eco3560, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3561(w_eco3561, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3562(w_eco3562, a[4], b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3563(w_eco3563, a[4], b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3564(w_eco3564, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3565(w_eco3565, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3566(w_eco3566, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3567(w_eco3567, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3568(w_eco3568, !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3569(w_eco3569, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3570(w_eco3570, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3571(w_eco3571, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3572(w_eco3572, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3573(w_eco3573, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3574(w_eco3574, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3575(w_eco3575, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3576(w_eco3576, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3577(w_eco3577, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3578(w_eco3578, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3579(w_eco3579, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3580(w_eco3580, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3581(w_eco3581, !a[4], !b[4], !a[5], !b[5], !b[6], a[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_3582(w_eco3582, !a[4], !b[4], !a[5], !b[5], !b[6], a[1], !b[1], a[2], !b[2], op[0], !op[1]);
	and _ECO_3583(w_eco3583, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3584(w_eco3584, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3585(w_eco3585, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3586(w_eco3586, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3587(w_eco3587, a[3], !b[3], !a[6], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3588(w_eco3588, a[3], !b[3], !a[6], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3589(w_eco3589, a[3], !b[3], !a[6], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3590(w_eco3590, a[3], !b[3], !a[6], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3591(w_eco3591, a[3], !b[3], !a[6], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3592(w_eco3592, a[3], !b[3], !a[6], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3593(w_eco3593, b[3], a[4], b[4], a[5], b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3594(w_eco3594, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3595(w_eco3595, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3596(w_eco3596, b[3], a[4], b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3597(w_eco3597, b[3], a[4], b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3598(w_eco3598, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3599(w_eco3599, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3600(w_eco3600, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3601(w_eco3601, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3602(w_eco3602, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3603(w_eco3603, !b[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3604(w_eco3604, !a[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3605(w_eco3605, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3606(w_eco3606, !a[3], a[4], b[4], a[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3607(w_eco3607, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3608(w_eco3608, !a[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3609(w_eco3609, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3610(w_eco3610, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3611(w_eco3611, a[3], !b[3], !a[4], b[5], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3612(w_eco3612, !a[3], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3613(w_eco3613, !a[3], b[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3614(w_eco3614, !b[1], a[2], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3615(w_eco3615, !b[1], a[2], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3616(w_eco3616, a[1], a[2], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3617(w_eco3617, a[1], a[2], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3618(w_eco3618, !a[3], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3619(w_eco3619, !a[3], !a[1], b[1], a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3620(w_eco3620, b[3], !b[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3621(w_eco3621, b[3], !b[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3622(w_eco3622, a[3], !b[3], !a[4], b[5], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3623(w_eco3623, a[3], !b[3], !a[4], b[5], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3624(w_eco3624, a[3], !b[3], !a[4], b[5], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3625(w_eco3625, !a[3], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3626(w_eco3626, !a[3], b[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3627(w_eco3627, !a[3], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3628(w_eco3628, !a[3], !b[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3629(w_eco3629, !a[3], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3630(w_eco3630, !a[3], a[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3631(w_eco3631, !a[3], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3632(w_eco3632, !a[3], !a[1], b[1], !a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3633(w_eco3633, !b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3634(w_eco3634, !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3635(w_eco3635, !b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3636(w_eco3636, !a[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3637(w_eco3637, !a[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3638(w_eco3638, !a[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3639(w_eco3639, !a[3], !b[3], a[5], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3640(w_eco3640, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3641(w_eco3641, !b[3], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3642(w_eco3642, !b[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3643(w_eco3643, !b[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3644(w_eco3644, !b[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3645(w_eco3645, !b[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3646(w_eco3646, !a[3], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3647(w_eco3647, !a[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3648(w_eco3648, !a[3], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3649(w_eco3649, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3650(w_eco3650, !a[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3651(w_eco3651, !a[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3652(w_eco3652, !a[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3653(w_eco3653, !b[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3654(w_eco3654, !a[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3655(w_eco3655, !b[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3656(w_eco3656, !a[3], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3657(w_eco3657, !a[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3658(w_eco3658, !a[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3659(w_eco3659, !a[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3660(w_eco3660, !a[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3661(w_eco3661, a[3], !b[3], !a[4], b[5], !a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3662(w_eco3662, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3663(w_eco3663, a[3], !b[3], !a[4], b[5], !a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3664(w_eco3664, a[3], !b[3], !a[4], b[5], !a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3665(w_eco3665, a[3], !b[3], !a[4], b[5], !a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3666(w_eco3666, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3667(w_eco3667, !a[4], !b[4], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3668(w_eco3668, !a[4], !b[4], a[6], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3669(w_eco3669, !a[4], !b[4], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3670(w_eco3670, !a[4], !b[4], a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3671(w_eco3671, !a[4], !b[4], a[6], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3672(w_eco3672, !a[4], !b[4], a[6], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3673(w_eco3673, !a[4], !b[4], a[6], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3674(w_eco3674, !a[4], !b[4], a[5], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3675(w_eco3675, !a[4], !b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3676(w_eco3676, !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3677(w_eco3677, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3678(w_eco3678, !a[4], !b[4], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3679(w_eco3679, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3680(w_eco3680, !a[4], !b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3681(w_eco3681, !a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3682(w_eco3682, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3683(w_eco3683, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3684(w_eco3684, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3685(w_eco3685, b[3], !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3686(w_eco3686, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3687(w_eco3687, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3688(w_eco3688, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3689(w_eco3689, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3690(w_eco3690, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3691(w_eco3691, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3692(w_eco3692, !a[4], !b[4], a[5], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3693(w_eco3693, !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3694(w_eco3694, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3695(w_eco3695, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], !a[7], !op[1]);
	and _ECO_3696(w_eco3696, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3697(w_eco3697, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3698(w_eco3698, !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3699(w_eco3699, !a[4], !b[4], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3700(w_eco3700, !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3701(w_eco3701, !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3702(w_eco3702, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3703(w_eco3703, !a[4], !b[4], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3704(w_eco3704, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3705(w_eco3705, !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3706(w_eco3706, a[3], !b[3], b[4], !a[5], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3707(w_eco3707, a[3], !b[3], b[4], !a[5], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3708(w_eco3708, a[3], !b[3], b[4], !a[5], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3709(w_eco3709, a[3], !b[3], b[4], !a[5], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3710(w_eco3710, !b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3711(w_eco3711, !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3712(w_eco3712, !b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3713(w_eco3713, !a[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3714(w_eco3714, !a[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3715(w_eco3715, !a[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3716(w_eco3716, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3717(w_eco3717, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3718(w_eco3718, !b[3], a[4], b[4], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3719(w_eco3719, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3720(w_eco3720, !b[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3721(w_eco3721, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3722(w_eco3722, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3723(w_eco3723, !a[3], a[4], b[4], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3724(w_eco3724, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3725(w_eco3725, !a[3], a[4], b[4], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3726(w_eco3726, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3727(w_eco3727, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3728(w_eco3728, !a[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3729(w_eco3729, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3730(w_eco3730, !b[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3731(w_eco3731, !a[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3732(w_eco3732, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3733(w_eco3733, !a[3], a[4], b[4], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3734(w_eco3734, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3735(w_eco3735, !a[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3736(w_eco3736, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3737(w_eco3737, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3738(w_eco3738, a[3], !b[3], b[4], !a[5], !a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3739(w_eco3739, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3740(w_eco3740, a[3], !b[3], b[4], !a[5], !a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3741(w_eco3741, a[3], !b[3], b[4], !a[5], !a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3742(w_eco3742, a[3], !b[3], b[4], !a[5], !a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3743(w_eco3743, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3744(w_eco3744, !b[3], a[6], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3745(w_eco3745, !a[3], a[6], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3746(w_eco3746, !b[3], a[6], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3747(w_eco3747, !a[3], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3748(w_eco3748, !a[3], a[6], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3749(w_eco3749, !a[3], a[6], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3750(w_eco3750, !a[3], a[6], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3751(w_eco3751, !a[3], a[6], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3752(w_eco3752, a[3], !b[3], !a[5], b[5], b[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3753(w_eco3753, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3754(w_eco3754, a[3], !b[3], !a[5], b[5], b[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3755(w_eco3755, a[3], !b[3], !a[5], b[5], b[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3756(w_eco3756, a[3], !b[3], !a[5], b[5], b[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3757(w_eco3757, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3758(w_eco3758, a[3], !b[3], !a[5], b[5], !a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3759(w_eco3759, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3760(w_eco3760, a[3], !b[3], !a[5], b[5], !a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3761(w_eco3761, a[3], !b[3], !a[5], b[5], !a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3762(w_eco3762, a[3], !b[3], !a[5], b[5], !a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3763(w_eco3763, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3764(w_eco3764, !a[4], !b[4], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3765(w_eco3765, !a[4], !b[4], a[6], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3766(w_eco3766, !a[4], !b[4], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3767(w_eco3767, !a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3768(w_eco3768, !a[4], !b[4], a[6], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3769(w_eco3769, !a[4], !b[4], a[6], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3770(w_eco3770, !a[4], !b[4], a[6], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3771(w_eco3771, !b[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3772(w_eco3772, !a[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3773(w_eco3773, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3774(w_eco3774, !a[3], a[4], b[4], a[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3775(w_eco3775, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3776(w_eco3776, !a[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3777(w_eco3777, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3778(w_eco3778, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3779(w_eco3779, !a[5], !b[5], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3780(w_eco3780, !a[5], !b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3781(w_eco3781, !a[5], !b[5], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3782(w_eco3782, !a[5], !b[5], a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3783(w_eco3783, !a[5], !b[5], a[6], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3784(w_eco3784, !a[5], !b[5], a[6], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3785(w_eco3785, !a[5], !b[5], a[6], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3786(w_eco3786, !a[5], !b[5], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3787(w_eco3787, !a[5], !b[5], a[6], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3788(w_eco3788, !a[5], !b[5], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3789(w_eco3789, !a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3790(w_eco3790, !a[5], !b[5], a[6], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3791(w_eco3791, !a[5], !b[5], a[6], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3792(w_eco3792, !a[5], !b[5], a[6], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3793(w_eco3793, b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3794(w_eco3794, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3795(w_eco3795, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3796(w_eco3796, b[3], a[4], b[4], !a[5], !b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3797(w_eco3797, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3798(w_eco3798, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3799(w_eco3799, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3800(w_eco3800, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3801(w_eco3801, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3802(w_eco3802, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3803(w_eco3803, b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3804(w_eco3804, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], a[2], b[2], op[0], !op[1]);
	and _ECO_3805(w_eco3805, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3806(w_eco3806, b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3807(w_eco3807, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3808(w_eco3808, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_3809(w_eco3809, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[2], op[0], !op[1]);
	and _ECO_3810(w_eco3810, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3811(w_eco3811, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3812(w_eco3812, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3813(w_eco3813, a[3], !b[3], !a[6], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3814(w_eco3814, a[3], !b[3], !a[6], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3815(w_eco3815, a[3], !b[3], !a[6], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3816(w_eco3816, a[3], !b[3], !a[6], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3817(w_eco3817, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3818(w_eco3818, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3819(w_eco3819, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3820(w_eco3820, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3821(w_eco3821, !b[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3822(w_eco3822, !b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3823(w_eco3823, !b[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3824(w_eco3824, !a[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3825(w_eco3825, !a[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3826(w_eco3826, !a[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3827(w_eco3827, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3828(w_eco3828, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3829(w_eco3829, !b[3], a[4], b[4], a[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3830(w_eco3830, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3831(w_eco3831, !b[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3832(w_eco3832, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3833(w_eco3833, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3834(w_eco3834, !a[3], a[4], b[4], a[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3835(w_eco3835, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3836(w_eco3836, !a[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3837(w_eco3837, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3838(w_eco3838, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3839(w_eco3839, !a[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3840(w_eco3840, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3841(w_eco3841, b[3], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3842(w_eco3842, b[3], b[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3843(w_eco3843, b[3], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3844(w_eco3844, b[3], !a[1], b[1], a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3845(w_eco3845, a[1], a[2], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3846(w_eco3846, a[1], a[2], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3847(w_eco3847, a[1], !b[1], a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3848(w_eco3848, a[1], !b[1], a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3849(w_eco3849, !a[3], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3850(w_eco3850, !a[3], !a[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3851(w_eco3851, b[3], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3852(w_eco3852, b[3], b[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3853(w_eco3853, b[3], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3854(w_eco3854, b[3], !b[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3855(w_eco3855, b[3], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3856(w_eco3856, b[3], a[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3857(w_eco3857, b[3], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3858(w_eco3858, b[3], !a[1], b[1], !a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3859(w_eco3859, !a[3], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3860(w_eco3860, !a[3], a[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3861(w_eco3861, !a[3], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_3862(w_eco3862, !a[3], a[1], !b[1], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_3863(w_eco3863, !a[3], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3864(w_eco3864, !a[3], !a[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3865(w_eco3865, !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3866(w_eco3866, !b[3], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3867(w_eco3867, !b[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3868(w_eco3868, !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3869(w_eco3869, !a[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3870(w_eco3870, !a[3], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3871(w_eco3871, !a[3], a[5], b[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3872(w_eco3872, !a[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3873(w_eco3873, !a[3], !b[3], a[5], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3874(w_eco3874, !a[3], !b[3], a[5], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3875(w_eco3875, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3876(w_eco3876, !b[3], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3877(w_eco3877, !b[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3878(w_eco3878, !b[3], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3879(w_eco3879, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3880(w_eco3880, !b[3], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3881(w_eco3881, !b[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3882(w_eco3882, !b[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3883(w_eco3883, !a[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3884(w_eco3884, !a[3], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3885(w_eco3885, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3886(w_eco3886, !b[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3887(w_eco3887, !b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3888(w_eco3888, !b[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3889(w_eco3889, !a[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3890(w_eco3890, !a[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3891(w_eco3891, !a[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3892(w_eco3892, !a[3], !b[3], a[5], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3893(w_eco3893, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3894(w_eco3894, !b[3], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3895(w_eco3895, !b[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3896(w_eco3896, !b[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3897(w_eco3897, !b[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3898(w_eco3898, !b[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3899(w_eco3899, !a[3], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3900(w_eco3900, !a[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3901(w_eco3901, !a[3], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3902(w_eco3902, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3903(w_eco3903, !a[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3904(w_eco3904, !a[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3905(w_eco3905, !a[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3906(w_eco3906, a[3], !b[3], !a[4], b[5], !a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3907(w_eco3907, a[3], !b[3], !a[4], b[5], !a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3908(w_eco3908, a[3], !b[3], !a[4], b[5], !a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3909(w_eco3909, a[3], !b[3], !a[4], b[5], !a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3910(w_eco3910, b[6], !b[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3911(w_eco3911, a[4], !b[4], a[5], !b[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_3912(w_eco3912, !a[6], !b[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_3913(w_eco3913, !a[4], !b[4], a[6], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3914(w_eco3914, !a[4], !b[4], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3915(w_eco3915, !a[4], !b[4], a[6], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3916(w_eco3916, !a[4], !b[4], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3917(w_eco3917, !a[4], !b[4], a[5], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3918(w_eco3918, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3919(w_eco3919, !a[4], !b[4], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3920(w_eco3920, !a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3921(w_eco3921, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3922(w_eco3922, !a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3923(w_eco3923, !a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3924(w_eco3924, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3925(w_eco3925, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3926(w_eco3926, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3927(w_eco3927, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3928(w_eco3928, !a[4], !b[4], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3929(w_eco3929, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3930(w_eco3930, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], !b[7], !op[1]);
	and _ECO_3931(w_eco3931, !a[4], !b[4], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3932(w_eco3932, !a[4], !b[4], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3933(w_eco3933, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3934(w_eco3934, !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3935(w_eco3935, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3936(w_eco3936, !b[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3937(w_eco3937, !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3938(w_eco3938, !a[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3939(w_eco3939, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3940(w_eco3940, !a[3], a[4], b[4], b[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3941(w_eco3941, !a[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3942(w_eco3942, !a[3], !b[3], a[4], b[4], b[5], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3943(w_eco3943, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3944(w_eco3944, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_3945(w_eco3945, !b[3], a[4], b[4], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3946(w_eco3946, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3947(w_eco3947, !b[3], a[4], b[4], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3948(w_eco3948, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], !a[7], !op[1]);
	and _ECO_3949(w_eco3949, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3950(w_eco3950, !b[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3951(w_eco3951, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3952(w_eco3952, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3953(w_eco3953, !a[3], a[4], b[4], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3954(w_eco3954, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_3955(w_eco3955, !b[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3956(w_eco3956, !b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3957(w_eco3957, !b[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3958(w_eco3958, !a[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3959(w_eco3959, !a[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3960(w_eco3960, !a[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3961(w_eco3961, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3962(w_eco3962, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3963(w_eco3963, !b[3], a[4], b[4], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3964(w_eco3964, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3965(w_eco3965, !b[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3966(w_eco3966, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3967(w_eco3967, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3968(w_eco3968, !a[3], a[4], b[4], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3969(w_eco3969, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3970(w_eco3970, !a[3], a[4], b[4], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3971(w_eco3971, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3972(w_eco3972, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3973(w_eco3973, !a[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3974(w_eco3974, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3975(w_eco3975, a[3], !b[3], b[4], !a[5], !a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3976(w_eco3976, a[3], !b[3], b[4], !a[5], !a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_3977(w_eco3977, a[3], !b[3], b[4], !a[5], !a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_3978(w_eco3978, a[3], !b[3], b[4], !a[5], !a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_3979(w_eco3979, !b[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3980(w_eco3980, !b[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3981(w_eco3981, !b[3], a[6], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3982(w_eco3982, !a[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3983(w_eco3983, !a[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3984(w_eco3984, !a[3], a[6], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3985(w_eco3985, !a[3], !b[3], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3986(w_eco3986, !a[3], !b[3], a[6], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3987(w_eco3987, !b[3], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3988(w_eco3988, !b[3], a[6], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3989(w_eco3989, !b[3], a[6], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_3990(w_eco3990, !b[3], a[6], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_3991(w_eco3991, !b[3], a[6], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_3992(w_eco3992, !a[3], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_3993(w_eco3993, !a[3], a[6], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_3994(w_eco3994, !a[3], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_3995(w_eco3995, !a[3], a[6], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_3996(w_eco3996, !a[3], a[6], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_3997(w_eco3997, !a[3], a[6], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_3998(w_eco3998, !a[3], a[6], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_3999(w_eco3999, a[3], !b[3], !a[5], b[5], b[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4000(w_eco4000, a[3], !b[3], !a[5], b[5], b[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4001(w_eco4001, a[3], !b[3], !a[5], b[5], b[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_4002(w_eco4002, a[3], !b[3], !a[5], b[5], b[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4003(w_eco4003, a[3], !b[3], !a[5], b[5], !a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4004(w_eco4004, a[3], !b[3], !a[5], b[5], !a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4005(w_eco4005, a[3], !b[3], !a[5], b[5], !a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_4006(w_eco4006, a[3], !b[3], !a[5], b[5], !a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4007(w_eco4007, !a[4], !b[4], a[6], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4008(w_eco4008, !a[4], !b[4], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4009(w_eco4009, !a[4], !b[4], a[6], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4010(w_eco4010, b[3], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4011(w_eco4011, b[3], !a[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4012(w_eco4012, b[3], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4013(w_eco4013, b[3], a[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4014(w_eco4014, b[3], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4015(w_eco4015, b[3], a[1], !b[1], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4016(w_eco4016, b[3], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4017(w_eco4017, b[3], !a[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4018(w_eco4018, !b[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4019(w_eco4019, !b[3], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4020(w_eco4020, !a[3], a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4021(w_eco4021, !a[3], a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4022(w_eco4022, !a[3], !b[3], a[5], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4023(w_eco4023, !b[3], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4024(w_eco4024, !b[3], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4025(w_eco4025, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4026(w_eco4026, !b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4027(w_eco4027, !b[3], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4028(w_eco4028, !b[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4029(w_eco4029, !b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4030(w_eco4030, !a[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4031(w_eco4031, !a[3], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4032(w_eco4032, !a[3], a[5], b[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4033(w_eco4033, !a[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4034(w_eco4034, !a[3], !b[3], a[5], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4035(w_eco4035, !a[3], !b[3], a[5], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4036(w_eco4036, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4037(w_eco4037, !b[3], a[5], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4038(w_eco4038, !b[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4039(w_eco4039, !b[3], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4040(w_eco4040, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4041(w_eco4041, !b[3], a[5], b[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4042(w_eco4042, !b[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4043(w_eco4043, !b[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4044(w_eco4044, !a[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4045(w_eco4045, !a[3], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4046(w_eco4046, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4047(w_eco4047, !b[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4048(w_eco4048, !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4049(w_eco4049, !b[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4050(w_eco4050, !a[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4051(w_eco4051, !a[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4052(w_eco4052, !a[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4053(w_eco4053, !a[3], !b[3], a[4], b[4], a[5], b[6], b[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4054(w_eco4054, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4055(w_eco4055, !b[3], a[4], b[4], a[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4056(w_eco4056, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4057(w_eco4057, !b[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4058(w_eco4058, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4059(w_eco4059, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4060(w_eco4060, !a[3], a[4], b[4], a[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4061(w_eco4061, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4062(w_eco4062, !a[3], a[4], b[4], a[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4063(w_eco4063, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4064(w_eco4064, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4065(w_eco4065, !a[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4066(w_eco4066, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4067(w_eco4067, a[5], !b[5], !b[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4068(w_eco4068, !a[5], !b[5], a[6], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4069(w_eco4069, !a[5], !b[5], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4070(w_eco4070, !a[5], !b[5], a[6], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4071(w_eco4071, !a[5], !b[5], a[6], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4072(w_eco4072, !a[5], !b[5], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4073(w_eco4073, !a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4074(w_eco4074, a[4], !b[4], !b[5], !b[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4075(w_eco4075, !b[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4076(w_eco4076, !b[3], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4077(w_eco4077, !a[3], a[5], b[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4078(w_eco4078, !a[3], a[5], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4079(w_eco4079, !a[3], !b[3], a[5], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4080(w_eco4080, !b[3], a[5], b[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4081(w_eco4081, !b[3], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4082(w_eco4082, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4083(w_eco4083, b[6], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4084(w_eco4084, b[6], b[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4085(w_eco4085, b[6], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4086(w_eco4086, b[6], !a[1], b[1], a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4087(w_eco4087, b[6], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4088(w_eco4088, b[6], b[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4089(w_eco4089, b[6], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4090(w_eco4090, b[6], a[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4091(w_eco4091, b[6], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4092(w_eco4092, b[6], !a[1], b[1], !a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4093(w_eco4093, a[4], !b[4], a[5], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4094(w_eco4094, a[4], !b[4], a[5], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4095(w_eco4095, a[4], !b[4], a[5], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4096(w_eco4096, a[4], !b[4], a[5], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4097(w_eco4097, b[6], !b[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4098(w_eco4098, a[4], !b[4], a[5], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4099(w_eco4099, a[4], !b[4], a[5], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4100(w_eco4100, !a[6], b[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4101(w_eco4101, !a[6], !a[1], b[1], a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4102(w_eco4102, !a[6], b[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4103(w_eco4103, !a[6], !b[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4104(w_eco4104, !a[6], a[1], !a[2], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4105(w_eco4105, !a[6], !a[1], b[1], !a[2], !b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4106(w_eco4106, !a[4], !b[4], a[5], b[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4107(w_eco4107, !a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4108(w_eco4108, !a[4], !b[4], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4109(w_eco4109, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4110(w_eco4110, !a[4], !b[4], a[5], b[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4111(w_eco4111, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4112(w_eco4112, !a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4113(w_eco4113, !b[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4114(w_eco4114, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4115(w_eco4115, !a[3], a[4], b[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4116(w_eco4116, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4117(w_eco4117, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4118(w_eco4118, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4119(w_eco4119, !b[3], a[4], b[4], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4120(w_eco4120, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4121(w_eco4121, !b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4122(w_eco4122, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4123(w_eco4123, !b[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4124(w_eco4124, !b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4125(w_eco4125, !a[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4126(w_eco4126, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4127(w_eco4127, !a[3], a[4], b[4], b[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4128(w_eco4128, !a[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4129(w_eco4129, !a[3], !b[3], a[4], b[4], b[5], a[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4130(w_eco4130, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4131(w_eco4131, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4132(w_eco4132, !b[3], a[4], b[4], b[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4133(w_eco4133, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4134(w_eco4134, !b[3], a[4], b[4], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4135(w_eco4135, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4136(w_eco4136, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4137(w_eco4137, !b[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4138(w_eco4138, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4139(w_eco4139, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4140(w_eco4140, !a[3], a[4], b[4], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4141(w_eco4141, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4142(w_eco4142, !b[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4143(w_eco4143, !b[3], a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4144(w_eco4144, !b[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4145(w_eco4145, !b[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4146(w_eco4146, !a[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4147(w_eco4147, !a[3], a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4148(w_eco4148, !a[3], a[6], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4149(w_eco4149, !a[3], a[6], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4150(w_eco4150, !a[3], !b[3], a[6], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4151(w_eco4151, !a[3], !b[3], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4152(w_eco4152, !a[3], !b[3], a[6], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4153(w_eco4153, !b[3], a[6], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4154(w_eco4154, !b[3], a[6], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4155(w_eco4155, !b[3], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4156(w_eco4156, !b[3], a[6], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4157(w_eco4157, !b[3], a[6], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4158(w_eco4158, !b[3], a[6], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4159(w_eco4159, !b[3], a[6], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4160(w_eco4160, !a[3], a[6], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4161(w_eco4161, !a[3], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4162(w_eco4162, !a[3], a[6], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4163(w_eco4163, b[6], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4164(w_eco4164, !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4165(w_eco4165, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4166(w_eco4166, !b[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4167(w_eco4167, !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4168(w_eco4168, !a[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4169(w_eco4169, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4170(w_eco4170, !a[3], a[4], b[4], a[5], b[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4171(w_eco4171, !a[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4172(w_eco4172, !a[3], !b[3], a[4], b[4], a[5], b[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4173(w_eco4173, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4174(w_eco4174, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4175(w_eco4175, !b[3], a[4], b[4], a[5], b[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4176(w_eco4176, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4177(w_eco4177, !b[3], a[4], b[4], a[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4178(w_eco4178, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4179(w_eco4179, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4180(w_eco4180, !b[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4181(w_eco4181, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4182(w_eco4182, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4183(w_eco4183, !a[3], a[4], b[4], a[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4184(w_eco4184, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4185(w_eco4185, a[5], !b[5], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4186(w_eco4186, a[5], !b[5], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4187(w_eco4187, a[5], !b[5], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4188(w_eco4188, a[5], !b[5], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4189(w_eco4189, a[5], !b[5], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4190(w_eco4190, a[5], !b[5], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4191(w_eco4191, !b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4192(w_eco4192, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4193(w_eco4193, !b[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4194(w_eco4194, !b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4195(w_eco4195, !a[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4196(w_eco4196, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[2], !b[2], !a[7], !op[0], !op[1]);
	and _ECO_4197(w_eco4197, !a[3], a[4], b[4], a[5], a[6], !b[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4198(w_eco4198, !a[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4199(w_eco4199, !a[3], !b[3], a[4], b[4], a[5], a[6], b[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4200(w_eco4200, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], a[2], b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4201(w_eco4201, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4202(w_eco4202, !b[3], a[4], b[4], a[5], a[6], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4203(w_eco4203, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4204(w_eco4204, !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4205(w_eco4205, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], b[2], !a[7], !op[0], !op[1]);
	and _ECO_4206(w_eco4206, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4207(w_eco4207, !b[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], !b[7], !op[0], !op[1]);
	and _ECO_4208(w_eco4208, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4209(w_eco4209, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4210(w_eco4210, !a[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4211(w_eco4211, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4212(w_eco4212, a[4], !b[4], !b[5], b[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4213(w_eco4213, a[4], !b[4], !b[5], !a[1], b[1], a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4214(w_eco4214, a[4], !b[4], !b[5], b[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4215(w_eco4215, a[4], !b[4], !b[5], !b[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4216(w_eco4216, a[4], !b[4], !b[5], a[1], !a[2], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4217(w_eco4217, a[4], !b[4], !b[5], !a[1], b[1], !a[2], !b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4218(w_eco4218, b[6], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4219(w_eco4219, b[6], !a[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4220(w_eco4220, b[6], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4221(w_eco4221, b[6], a[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4222(w_eco4222, b[6], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4223(w_eco4223, b[6], a[1], !b[1], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4224(w_eco4224, b[6], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4225(w_eco4225, b[6], !a[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4226(w_eco4226, !b[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4227(w_eco4227, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4228(w_eco4228, !a[3], a[4], b[4], a[5], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4229(w_eco4229, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4230(w_eco4230, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4231(w_eco4231, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4232(w_eco4232, !b[3], a[4], b[4], a[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4233(w_eco4233, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4234(w_eco4234, a[4], !b[4], a[5], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4235(w_eco4235, a[4], !b[4], a[5], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4236(w_eco4236, a[4], !b[4], a[5], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4237(w_eco4237, a[4], !b[4], a[5], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4238(w_eco4238, !a[6], !a[1], a[2], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4239(w_eco4239, !a[6], a[1], !a[2], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4240(w_eco4240, !a[6], a[1], !b[1], !a[2], b[2], !a[7], b[7], op[0], !op[1]);
	and _ECO_4241(w_eco4241, !a[6], !a[1], !a[2], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4242(w_eco4242, a[5], !b[5], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4243(w_eco4243, a[5], !b[5], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4244(w_eco4244, a[5], !b[5], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4245(w_eco4245, a[5], !b[5], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4246(w_eco4246, a[4], !b[4], !b[5], !a[1], a[2], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4247(w_eco4247, a[4], !b[4], !b[5], a[1], !a[2], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4248(w_eco4248, a[4], !b[4], !b[5], a[1], !b[1], !a[2], b[2], a[7], !b[7], op[0], !op[1]);
	and _ECO_4249(w_eco4249, a[4], !b[4], !b[5], !a[1], !a[2], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4250(w_eco4250, !a[4], !b[4], a[5], b[5], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4251(w_eco4251, !a[4], !b[4], a[5], b[5], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4252(w_eco4252, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4253(w_eco4253, !b[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4254(w_eco4254, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4255(w_eco4255, !a[3], a[4], b[4], b[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4256(w_eco4256, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4257(w_eco4257, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4258(w_eco4258, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4259(w_eco4259, !b[3], a[4], b[4], b[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4260(w_eco4260, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4261(w_eco4261, !b[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4262(w_eco4262, !b[3], a[6], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4263(w_eco4263, !a[3], a[6], b[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4264(w_eco4264, !a[3], a[6], b[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4265(w_eco4265, !a[3], !b[3], a[6], b[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4266(w_eco4266, !b[3], a[6], b[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4267(w_eco4267, !b[3], a[6], b[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4268(w_eco4268, !b[3], a[6], b[6], !a[1], !b[1], !a[2], b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4269(w_eco4269, !b[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4270(w_eco4270, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4271(w_eco4271, !a[3], a[4], b[4], a[5], a[6], !a[1], a[2], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4272(w_eco4272, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[2], !b[2], a[0], a[7], !b[7], !op[1]);
	and _ECO_4273(w_eco4273, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], a[2], b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4274(w_eco4274, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4275(w_eco4275, !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4276(w_eco4276, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], b[2], !b[7], !op[0], !op[1]);
	and _ECO_4277(w_eco4277, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4278(w_eco4278, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4279(w_eco4279, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_4280(w_eco4280, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4281(w_eco4281, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4282(w_eco4282, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4283(w_eco4283, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !a[2], b[2], op[0], !op[1]);
	and _ECO_4284(w_eco4284, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	or _ECO_4285(w_eco4285, w_eco3339, w_eco3340, w_eco3341, w_eco3342, w_eco3343, w_eco3344, w_eco3345, w_eco3346, w_eco3347, w_eco3348, w_eco3349, w_eco3350, w_eco3351, w_eco3352, w_eco3353, w_eco3354, w_eco3355, w_eco3356, w_eco3357, w_eco3358, w_eco3359, w_eco3360, w_eco3361, w_eco3362, w_eco3363, w_eco3364, w_eco3365, w_eco3366, w_eco3367, w_eco3368, w_eco3369, w_eco3370, w_eco3371, w_eco3372, w_eco3373, w_eco3374, w_eco3375, w_eco3376, w_eco3377, w_eco3378, w_eco3379, w_eco3380, w_eco3381, w_eco3382, w_eco3383, w_eco3384, w_eco3385, w_eco3386, w_eco3387, w_eco3388, w_eco3389, w_eco3390, w_eco3391, w_eco3392, w_eco3393, w_eco3394, w_eco3395, w_eco3396, w_eco3397, w_eco3398, w_eco3399, w_eco3400, w_eco3401, w_eco3402, w_eco3403, w_eco3404, w_eco3405, w_eco3406, w_eco3407, w_eco3408, w_eco3409, w_eco3410, w_eco3411, w_eco3412, w_eco3413, w_eco3414, w_eco3415, w_eco3416, w_eco3417, w_eco3418, w_eco3419, w_eco3420, w_eco3421, w_eco3422, w_eco3423, w_eco3424, w_eco3425, w_eco3426, w_eco3427, w_eco3428, w_eco3429, w_eco3430, w_eco3431, w_eco3432, w_eco3433, w_eco3434, w_eco3435, w_eco3436, w_eco3437, w_eco3438, w_eco3439, w_eco3440, w_eco3441, w_eco3442, w_eco3443, w_eco3444, w_eco3445, w_eco3446, w_eco3447, w_eco3448, w_eco3449, w_eco3450, w_eco3451, w_eco3452, w_eco3453, w_eco3454, w_eco3455, w_eco3456, w_eco3457, w_eco3458, w_eco3459, w_eco3460, w_eco3461, w_eco3462, w_eco3463, w_eco3464, w_eco3465, w_eco3466, w_eco3467, w_eco3468, w_eco3469, w_eco3470, w_eco3471, w_eco3472, w_eco3473, w_eco3474, w_eco3475, w_eco3476, w_eco3477, w_eco3478, w_eco3479, w_eco3480, w_eco3481, w_eco3482, w_eco3483, w_eco3484, w_eco3485, w_eco3486, w_eco3487, w_eco3488, w_eco3489, w_eco3490, w_eco3491, w_eco3492, w_eco3493, w_eco3494, w_eco3495, w_eco3496, w_eco3497, w_eco3498, w_eco3499, w_eco3500, w_eco3501, w_eco3502, w_eco3503, w_eco3504, w_eco3505, w_eco3506, w_eco3507, w_eco3508, w_eco3509, w_eco3510, w_eco3511, w_eco3512, w_eco3513, w_eco3514, w_eco3515, w_eco3516, w_eco3517, w_eco3518, w_eco3519, w_eco3520, w_eco3521, w_eco3522, w_eco3523, w_eco3524, w_eco3525, w_eco3526, w_eco3527, w_eco3528, w_eco3529, w_eco3530, w_eco3531, w_eco3532, w_eco3533, w_eco3534, w_eco3535, w_eco3536, w_eco3537, w_eco3538, w_eco3539, w_eco3540, w_eco3541, w_eco3542, w_eco3543, w_eco3544, w_eco3545, w_eco3546, w_eco3547, w_eco3548, w_eco3549, w_eco3550, w_eco3551, w_eco3552, w_eco3553, w_eco3554, w_eco3555, w_eco3556, w_eco3557, w_eco3558, w_eco3559, w_eco3560, w_eco3561, w_eco3562, w_eco3563, w_eco3564, w_eco3565, w_eco3566, w_eco3567, w_eco3568, w_eco3569, w_eco3570, w_eco3571, w_eco3572, w_eco3573, w_eco3574, w_eco3575, w_eco3576, w_eco3577, w_eco3578, w_eco3579, w_eco3580, w_eco3581, w_eco3582, w_eco3583, w_eco3584, w_eco3585, w_eco3586, w_eco3587, w_eco3588, w_eco3589, w_eco3590, w_eco3591, w_eco3592, w_eco3593, w_eco3594, w_eco3595, w_eco3596, w_eco3597, w_eco3598, w_eco3599, w_eco3600, w_eco3601, w_eco3602, w_eco3603, w_eco3604, w_eco3605, w_eco3606, w_eco3607, w_eco3608, w_eco3609, w_eco3610, w_eco3611, w_eco3612, w_eco3613, w_eco3614, w_eco3615, w_eco3616, w_eco3617, w_eco3618, w_eco3619, w_eco3620, w_eco3621, w_eco3622, w_eco3623, w_eco3624, w_eco3625, w_eco3626, w_eco3627, w_eco3628, w_eco3629, w_eco3630, w_eco3631, w_eco3632, w_eco3633, w_eco3634, w_eco3635, w_eco3636, w_eco3637, w_eco3638, w_eco3639, w_eco3640, w_eco3641, w_eco3642, w_eco3643, w_eco3644, w_eco3645, w_eco3646, w_eco3647, w_eco3648, w_eco3649, w_eco3650, w_eco3651, w_eco3652, w_eco3653, w_eco3654, w_eco3655, w_eco3656, w_eco3657, w_eco3658, w_eco3659, w_eco3660, w_eco3661, w_eco3662, w_eco3663, w_eco3664, w_eco3665, w_eco3666, w_eco3667, w_eco3668, w_eco3669, w_eco3670, w_eco3671, w_eco3672, w_eco3673, w_eco3674, w_eco3675, w_eco3676, w_eco3677, w_eco3678, w_eco3679, w_eco3680, w_eco3681, w_eco3682, w_eco3683, w_eco3684, w_eco3685, w_eco3686, w_eco3687, w_eco3688, w_eco3689, w_eco3690, w_eco3691, w_eco3692, w_eco3693, w_eco3694, w_eco3695, w_eco3696, w_eco3697, w_eco3698, w_eco3699, w_eco3700, w_eco3701, w_eco3702, w_eco3703, w_eco3704, w_eco3705, w_eco3706, w_eco3707, w_eco3708, w_eco3709, w_eco3710, w_eco3711, w_eco3712, w_eco3713, w_eco3714, w_eco3715, w_eco3716, w_eco3717, w_eco3718, w_eco3719, w_eco3720, w_eco3721, w_eco3722, w_eco3723, w_eco3724, w_eco3725, w_eco3726, w_eco3727, w_eco3728, w_eco3729, w_eco3730, w_eco3731, w_eco3732, w_eco3733, w_eco3734, w_eco3735, w_eco3736, w_eco3737, w_eco3738, w_eco3739, w_eco3740, w_eco3741, w_eco3742, w_eco3743, w_eco3744, w_eco3745, w_eco3746, w_eco3747, w_eco3748, w_eco3749, w_eco3750, w_eco3751, w_eco3752, w_eco3753, w_eco3754, w_eco3755, w_eco3756, w_eco3757, w_eco3758, w_eco3759, w_eco3760, w_eco3761, w_eco3762, w_eco3763, w_eco3764, w_eco3765, w_eco3766, w_eco3767, w_eco3768, w_eco3769, w_eco3770, w_eco3771, w_eco3772, w_eco3773, w_eco3774, w_eco3775, w_eco3776, w_eco3777, w_eco3778, w_eco3779, w_eco3780, w_eco3781, w_eco3782, w_eco3783, w_eco3784, w_eco3785, w_eco3786, w_eco3787, w_eco3788, w_eco3789, w_eco3790, w_eco3791, w_eco3792, w_eco3793, w_eco3794, w_eco3795, w_eco3796, w_eco3797, w_eco3798, w_eco3799, w_eco3800, w_eco3801, w_eco3802, w_eco3803, w_eco3804, w_eco3805, w_eco3806, w_eco3807, w_eco3808, w_eco3809, w_eco3810, w_eco3811, w_eco3812, w_eco3813, w_eco3814, w_eco3815, w_eco3816, w_eco3817, w_eco3818, w_eco3819, w_eco3820, w_eco3821, w_eco3822, w_eco3823, w_eco3824, w_eco3825, w_eco3826, w_eco3827, w_eco3828, w_eco3829, w_eco3830, w_eco3831, w_eco3832, w_eco3833, w_eco3834, w_eco3835, w_eco3836, w_eco3837, w_eco3838, w_eco3839, w_eco3840, w_eco3841, w_eco3842, w_eco3843, w_eco3844, w_eco3845, w_eco3846, w_eco3847, w_eco3848, w_eco3849, w_eco3850, w_eco3851, w_eco3852, w_eco3853, w_eco3854, w_eco3855, w_eco3856, w_eco3857, w_eco3858, w_eco3859, w_eco3860, w_eco3861, w_eco3862, w_eco3863, w_eco3864, w_eco3865, w_eco3866, w_eco3867, w_eco3868, w_eco3869, w_eco3870, w_eco3871, w_eco3872, w_eco3873, w_eco3874, w_eco3875, w_eco3876, w_eco3877, w_eco3878, w_eco3879, w_eco3880, w_eco3881, w_eco3882, w_eco3883, w_eco3884, w_eco3885, w_eco3886, w_eco3887, w_eco3888, w_eco3889, w_eco3890, w_eco3891, w_eco3892, w_eco3893, w_eco3894, w_eco3895, w_eco3896, w_eco3897, w_eco3898, w_eco3899, w_eco3900, w_eco3901, w_eco3902, w_eco3903, w_eco3904, w_eco3905, w_eco3906, w_eco3907, w_eco3908, w_eco3909, w_eco3910, w_eco3911, w_eco3912, w_eco3913, w_eco3914, w_eco3915, w_eco3916, w_eco3917, w_eco3918, w_eco3919, w_eco3920, w_eco3921, w_eco3922, w_eco3923, w_eco3924, w_eco3925, w_eco3926, w_eco3927, w_eco3928, w_eco3929, w_eco3930, w_eco3931, w_eco3932, w_eco3933, w_eco3934, w_eco3935, w_eco3936, w_eco3937, w_eco3938, w_eco3939, w_eco3940, w_eco3941, w_eco3942, w_eco3943, w_eco3944, w_eco3945, w_eco3946, w_eco3947, w_eco3948, w_eco3949, w_eco3950, w_eco3951, w_eco3952, w_eco3953, w_eco3954, w_eco3955, w_eco3956, w_eco3957, w_eco3958, w_eco3959, w_eco3960, w_eco3961, w_eco3962, w_eco3963, w_eco3964, w_eco3965, w_eco3966, w_eco3967, w_eco3968, w_eco3969, w_eco3970, w_eco3971, w_eco3972, w_eco3973, w_eco3974, w_eco3975, w_eco3976, w_eco3977, w_eco3978, w_eco3979, w_eco3980, w_eco3981, w_eco3982, w_eco3983, w_eco3984, w_eco3985, w_eco3986, w_eco3987, w_eco3988, w_eco3989, w_eco3990, w_eco3991, w_eco3992, w_eco3993, w_eco3994, w_eco3995, w_eco3996, w_eco3997, w_eco3998, w_eco3999, w_eco4000, w_eco4001, w_eco4002, w_eco4003, w_eco4004, w_eco4005, w_eco4006, w_eco4007, w_eco4008, w_eco4009, w_eco4010, w_eco4011, w_eco4012, w_eco4013, w_eco4014, w_eco4015, w_eco4016, w_eco4017, w_eco4018, w_eco4019, w_eco4020, w_eco4021, w_eco4022, w_eco4023, w_eco4024, w_eco4025, w_eco4026, w_eco4027, w_eco4028, w_eco4029, w_eco4030, w_eco4031, w_eco4032, w_eco4033, w_eco4034, w_eco4035, w_eco4036, w_eco4037, w_eco4038, w_eco4039, w_eco4040, w_eco4041, w_eco4042, w_eco4043, w_eco4044, w_eco4045, w_eco4046, w_eco4047, w_eco4048, w_eco4049, w_eco4050, w_eco4051, w_eco4052, w_eco4053, w_eco4054, w_eco4055, w_eco4056, w_eco4057, w_eco4058, w_eco4059, w_eco4060, w_eco4061, w_eco4062, w_eco4063, w_eco4064, w_eco4065, w_eco4066, w_eco4067, w_eco4068, w_eco4069, w_eco4070, w_eco4071, w_eco4072, w_eco4073, w_eco4074, w_eco4075, w_eco4076, w_eco4077, w_eco4078, w_eco4079, w_eco4080, w_eco4081, w_eco4082, w_eco4083, w_eco4084, w_eco4085, w_eco4086, w_eco4087, w_eco4088, w_eco4089, w_eco4090, w_eco4091, w_eco4092, w_eco4093, w_eco4094, w_eco4095, w_eco4096, w_eco4097, w_eco4098, w_eco4099, w_eco4100, w_eco4101, w_eco4102, w_eco4103, w_eco4104, w_eco4105, w_eco4106, w_eco4107, w_eco4108, w_eco4109, w_eco4110, w_eco4111, w_eco4112, w_eco4113, w_eco4114, w_eco4115, w_eco4116, w_eco4117, w_eco4118, w_eco4119, w_eco4120, w_eco4121, w_eco4122, w_eco4123, w_eco4124, w_eco4125, w_eco4126, w_eco4127, w_eco4128, w_eco4129, w_eco4130, w_eco4131, w_eco4132, w_eco4133, w_eco4134, w_eco4135, w_eco4136, w_eco4137, w_eco4138, w_eco4139, w_eco4140, w_eco4141, w_eco4142, w_eco4143, w_eco4144, w_eco4145, w_eco4146, w_eco4147, w_eco4148, w_eco4149, w_eco4150, w_eco4151, w_eco4152, w_eco4153, w_eco4154, w_eco4155, w_eco4156, w_eco4157, w_eco4158, w_eco4159, w_eco4160, w_eco4161, w_eco4162, w_eco4163, w_eco4164, w_eco4165, w_eco4166, w_eco4167, w_eco4168, w_eco4169, w_eco4170, w_eco4171, w_eco4172, w_eco4173, w_eco4174, w_eco4175, w_eco4176, w_eco4177, w_eco4178, w_eco4179, w_eco4180, w_eco4181, w_eco4182, w_eco4183, w_eco4184, w_eco4185, w_eco4186, w_eco4187, w_eco4188, w_eco4189, w_eco4190, w_eco4191, w_eco4192, w_eco4193, w_eco4194, w_eco4195, w_eco4196, w_eco4197, w_eco4198, w_eco4199, w_eco4200, w_eco4201, w_eco4202, w_eco4203, w_eco4204, w_eco4205, w_eco4206, w_eco4207, w_eco4208, w_eco4209, w_eco4210, w_eco4211, w_eco4212, w_eco4213, w_eco4214, w_eco4215, w_eco4216, w_eco4217, w_eco4218, w_eco4219, w_eco4220, w_eco4221, w_eco4222, w_eco4223, w_eco4224, w_eco4225, w_eco4226, w_eco4227, w_eco4228, w_eco4229, w_eco4230, w_eco4231, w_eco4232, w_eco4233, w_eco4234, w_eco4235, w_eco4236, w_eco4237, w_eco4238, w_eco4239, w_eco4240, w_eco4241, w_eco4242, w_eco4243, w_eco4244, w_eco4245, w_eco4246, w_eco4247, w_eco4248, w_eco4249, w_eco4250, w_eco4251, w_eco4252, w_eco4253, w_eco4254, w_eco4255, w_eco4256, w_eco4257, w_eco4258, w_eco4259, w_eco4260, w_eco4261, w_eco4262, w_eco4263, w_eco4264, w_eco4265, w_eco4266, w_eco4267, w_eco4268, w_eco4269, w_eco4270, w_eco4271, w_eco4272, w_eco4273, w_eco4274, w_eco4275, w_eco4276, w_eco4277, w_eco4278, w_eco4279, w_eco4280, w_eco4281, w_eco4282, w_eco4283, w_eco4284);
	xor _ECO_out7(y[2], sub_wire7, w_eco4285);
	and _ECO_4286(w_eco4286, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4287(w_eco4287, a[4], b[4], a[5], b[5], a[6], b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4288(w_eco4288, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4289(w_eco4289, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4290(w_eco4290, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4291(w_eco4291, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4292(w_eco4292, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4293(w_eco4293, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4294(w_eco4294, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4295(w_eco4295, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4296(w_eco4296, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4297(w_eco4297, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4298(w_eco4298, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4299(w_eco4299, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4300(w_eco4300, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4301(w_eco4301, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4302(w_eco4302, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4303(w_eco4303, a[4], b[4], a[5], b[5], a[6], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4304(w_eco4304, a[4], b[4], a[5], b[5], a[6], b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4305(w_eco4305, a[4], b[4], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4306(w_eco4306, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4307(w_eco4307, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4308(w_eco4308, a[4], b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4309(w_eco4309, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4310(w_eco4310, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4311(w_eco4311, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4312(w_eco4312, !a[4], !b[4], a[5], b[5], a[6], b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4313(w_eco4313, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4314(w_eco4314, !a[4], !b[4], a[6], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4315(w_eco4315, !a[4], !b[4], a[6], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4316(w_eco4316, !a[4], !b[4], a[5], b[5], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4317(w_eco4317, !a[4], !b[4], a[5], b[5], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4318(w_eco4318, !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4319(w_eco4319, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4320(w_eco4320, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4321(w_eco4321, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4322(w_eco4322, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4323(w_eco4323, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4324(w_eco4324, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4325(w_eco4325, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4326(w_eco4326, a[4], b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4327(w_eco4327, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4328(w_eco4328, !a[5], !b[5], a[6], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4329(w_eco4329, !a[5], !b[5], a[6], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4330(w_eco4330, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4331(w_eco4331, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4332(w_eco4332, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4333(w_eco4333, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4334(w_eco4334, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4335(w_eco4335, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4336(w_eco4336, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4337(w_eco4337, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4338(w_eco4338, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4339(w_eco4339, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4340(w_eco4340, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4341(w_eco4341, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4342(w_eco4342, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4343(w_eco4343, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4344(w_eco4344, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4345(w_eco4345, b[6], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4346(w_eco4346, b[6], !a[1], b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4347(w_eco4347, b[6], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4348(w_eco4348, b[6], a[1], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4349(w_eco4349, !a[6], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4350(w_eco4350, !a[6], !a[1], b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4351(w_eco4351, !a[6], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4352(w_eco4352, !a[6], a[1], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4353(w_eco4353, !a[4], !b[4], a[6], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4354(w_eco4354, !a[4], !b[4], a[6], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4355(w_eco4355, !a[4], !b[4], a[6], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4356(w_eco4356, !a[4], !b[4], a[6], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4357(w_eco4357, !a[4], !b[4], a[6], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4358(w_eco4358, !a[4], !b[4], a[6], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4359(w_eco4359, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4360(w_eco4360, !a[4], !b[4], a[5], b[5], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4361(w_eco4361, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4362(w_eco4362, !a[4], !b[4], a[5], b[5], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4363(w_eco4363, !a[4], !b[4], a[5], b[5], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4364(w_eco4364, !a[4], !b[4], a[5], b[5], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4365(w_eco4365, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4366(w_eco4366, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4367(w_eco4367, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4368(w_eco4368, !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4369(w_eco4369, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4370(w_eco4370, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4371(w_eco4371, !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4372(w_eco4372, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4373(w_eco4373, !a[5], !b[5], a[6], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4374(w_eco4374, !a[5], !b[5], a[6], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4375(w_eco4375, !a[5], !b[5], a[6], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4376(w_eco4376, !a[5], !b[5], a[6], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4377(w_eco4377, !a[5], !b[5], a[6], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4378(w_eco4378, !a[5], !b[5], a[6], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4379(w_eco4379, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4380(w_eco4380, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4381(w_eco4381, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4382(w_eco4382, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4383(w_eco4383, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4384(w_eco4384, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_4385(w_eco4385, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4386(w_eco4386, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4387(w_eco4387, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4388(w_eco4388, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4389(w_eco4389, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4390(w_eco4390, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4391(w_eco4391, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4392(w_eco4392, a[3], !b[3], !a[4], b[5], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4393(w_eco4393, a[3], !b[3], !a[4], b[5], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4394(w_eco4394, !a[3], !b[3], a[5], b[5], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4395(w_eco4395, !a[3], !b[3], a[5], b[5], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4396(w_eco4396, !b[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4397(w_eco4397, !b[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4398(w_eco4398, !a[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4399(w_eco4399, !a[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4400(w_eco4400, b[6], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4401(w_eco4401, b[6], !a[1], b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4402(w_eco4402, b[6], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4403(w_eco4403, b[6], a[1], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4404(w_eco4404, b[6], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4405(w_eco4405, b[6], a[1], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4406(w_eco4406, b[6], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4407(w_eco4407, b[6], !a[1], !b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4408(w_eco4408, !a[6], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4409(w_eco4409, !a[6], !a[1], b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4410(w_eco4410, !a[6], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4411(w_eco4411, !a[6], a[1], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4412(w_eco4412, !a[6], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4413(w_eco4413, !a[6], a[1], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4414(w_eco4414, !a[6], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4415(w_eco4415, !a[6], !a[1], !b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4416(w_eco4416, !a[4], !b[4], a[6], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4417(w_eco4417, !a[4], !b[4], a[6], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4418(w_eco4418, !a[4], !b[4], a[6], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4419(w_eco4419, !a[4], !b[4], a[6], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4420(w_eco4420, !a[4], !b[4], a[5], b[5], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4421(w_eco4421, !a[4], !b[4], a[5], b[5], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4422(w_eco4422, !a[4], !b[4], a[5], b[5], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4423(w_eco4423, !a[4], !b[4], a[5], b[5], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4424(w_eco4424, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4425(w_eco4425, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_4426(w_eco4426, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4427(w_eco4427, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4428(w_eco4428, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4429(w_eco4429, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4430(w_eco4430, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4431(w_eco4431, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4432(w_eco4432, !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4433(w_eco4433, !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4434(w_eco4434, !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4435(w_eco4435, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4436(w_eco4436, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4437(w_eco4437, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4438(w_eco4438, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[1]);
	and _ECO_4439(w_eco4439, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4440(w_eco4440, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4441(w_eco4441, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4442(w_eco4442, !a[5], !b[5], a[6], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4443(w_eco4443, !a[5], !b[5], a[6], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4444(w_eco4444, !a[5], !b[5], a[6], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4445(w_eco4445, !a[5], !b[5], a[6], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4446(w_eco4446, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4447(w_eco4447, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_4448(w_eco4448, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4449(w_eco4449, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4450(w_eco4450, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4451(w_eco4451, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4452(w_eco4452, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4453(w_eco4453, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4454(w_eco4454, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[0], op[0], !op[1]);
	and _ECO_4455(w_eco4455, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !b[0], op[0], !op[1]);
	and _ECO_4456(w_eco4456, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4457(w_eco4457, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], !b[0], op[0], !op[1]);
	and _ECO_4458(w_eco4458, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4459(w_eco4459, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4460(w_eco4460, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4461(w_eco4461, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4462(w_eco4462, b[3], a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4463(w_eco4463, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4464(w_eco4464, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_4465(w_eco4465, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4466(w_eco4466, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4467(w_eco4467, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4468(w_eco4468, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4469(w_eco4469, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4470(w_eco4470, b[3], a[4], b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4471(w_eco4471, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4472(w_eco4472, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4473(w_eco4473, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4474(w_eco4474, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4475(w_eco4475, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4476(w_eco4476, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4477(w_eco4477, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4478(w_eco4478, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4479(w_eco4479, !b[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4480(w_eco4480, !b[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4481(w_eco4481, !a[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4482(w_eco4482, !a[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4483(w_eco4483, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4484(w_eco4484, !a[3], !b[3], a[5], b[5], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4485(w_eco4485, !a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4486(w_eco4486, !a[3], !b[3], a[5], b[5], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4487(w_eco4487, !a[3], !b[3], a[5], b[5], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4488(w_eco4488, !a[3], !b[3], a[5], b[5], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4489(w_eco4489, !b[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4490(w_eco4490, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4491(w_eco4491, !b[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4492(w_eco4492, !b[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4493(w_eco4493, !b[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4494(w_eco4494, !a[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4495(w_eco4495, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4496(w_eco4496, !a[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4497(w_eco4497, !a[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4498(w_eco4498, !a[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4499(w_eco4499, !a[3], !a[1], b[1], !a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4500(w_eco4500, !a[3], !a[1], b[1], !a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4501(w_eco4501, !a[3], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4502(w_eco4502, !a[3], a[1], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4503(w_eco4503, !a[3], !b[3], a[5], b[5], a[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4504(w_eco4504, !a[3], !b[3], a[5], b[5], a[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4505(w_eco4505, !b[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4506(w_eco4506, !b[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4507(w_eco4507, !a[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4508(w_eco4508, !a[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4509(w_eco4509, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4510(w_eco4510, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4511(w_eco4511, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_4512(w_eco4512, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4513(w_eco4513, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4514(w_eco4514, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4515(w_eco4515, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4516(w_eco4516, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4517(w_eco4517, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4518(w_eco4518, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4519(w_eco4519, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4520(w_eco4520, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4521(w_eco4521, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[1]);
	and _ECO_4522(w_eco4522, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4523(w_eco4523, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4524(w_eco4524, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4525(w_eco4525, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4526(w_eco4526, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4527(w_eco4527, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4528(w_eco4528, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4529(w_eco4529, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4530(w_eco4530, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4531(w_eco4531, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4532(w_eco4532, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4533(w_eco4533, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4534(w_eco4534, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4535(w_eco4535, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4536(w_eco4536, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4537(w_eco4537, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4538(w_eco4538, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4539(w_eco4539, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4540(w_eco4540, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4541(w_eco4541, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4542(w_eco4542, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4543(w_eco4543, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4544(w_eco4544, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4545(w_eco4545, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4546(w_eco4546, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4547(w_eco4547, !a[3], !b[3], a[6], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4548(w_eco4548, !a[3], !b[3], a[6], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4549(w_eco4549, !b[3], a[6], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4550(w_eco4550, !b[3], a[6], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4551(w_eco4551, !a[3], a[6], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4552(w_eco4552, !a[3], a[6], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4553(w_eco4553, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4554(w_eco4554, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4555(w_eco4555, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4556(w_eco4556, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4557(w_eco4557, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4558(w_eco4558, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4559(w_eco4559, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4560(w_eco4560, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4561(w_eco4561, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_4562(w_eco4562, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4563(w_eco4563, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4564(w_eco4564, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4565(w_eco4565, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4566(w_eco4566, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4567(w_eco4567, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4568(w_eco4568, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4569(w_eco4569, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4570(w_eco4570, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[0], op[0], !op[1]);
	and _ECO_4571(w_eco4571, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4572(w_eco4572, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], a[0], op[0], !op[1]);
	and _ECO_4573(w_eco4573, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4574(w_eco4574, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4575(w_eco4575, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4576(w_eco4576, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], !b[0], op[0], !op[1]);
	and _ECO_4577(w_eco4577, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], !a[2], a[0], op[0], !op[1]);
	and _ECO_4578(w_eco4578, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4579(w_eco4579, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !b[1], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4580(w_eco4580, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4581(w_eco4581, a[3], !b[3], !a[6], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4582(w_eco4582, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4583(w_eco4583, b[3], a[4], b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4584(w_eco4584, b[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4585(w_eco4585, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4586(w_eco4586, !a[3], a[4], b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4587(w_eco4587, !a[3], a[4], b[4], a[5], b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4588(w_eco4588, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_4589(w_eco4589, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4590(w_eco4590, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4591(w_eco4591, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4592(w_eco4592, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4593(w_eco4593, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4594(w_eco4594, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4595(w_eco4595, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4596(w_eco4596, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4597(w_eco4597, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4598(w_eco4598, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4599(w_eco4599, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4600(w_eco4600, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4601(w_eco4601, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4602(w_eco4602, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4603(w_eco4603, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4604(w_eco4604, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4605(w_eco4605, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4606(w_eco4606, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4607(w_eco4607, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4608(w_eco4608, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4609(w_eco4609, a[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4610(w_eco4610, !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4611(w_eco4611, a[3], !b[3], !a[4], b[5], b[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4612(w_eco4612, !b[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4613(w_eco4613, !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4614(w_eco4614, !b[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4615(w_eco4615, !b[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4616(w_eco4616, !b[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4617(w_eco4617, !a[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4618(w_eco4618, !a[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4619(w_eco4619, !a[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4620(w_eco4620, !a[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4621(w_eco4621, !a[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4622(w_eco4622, !a[3], !b[3], a[5], b[5], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4623(w_eco4623, !a[3], !b[3], a[5], b[5], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4624(w_eco4624, !a[3], !b[3], a[5], b[5], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4625(w_eco4625, !a[3], !b[3], a[5], b[5], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4626(w_eco4626, !b[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4627(w_eco4627, !b[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4628(w_eco4628, !b[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4629(w_eco4629, !b[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4630(w_eco4630, !a[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4631(w_eco4631, !a[3], a[5], b[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4632(w_eco4632, !a[3], a[5], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4633(w_eco4633, !a[3], a[5], b[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4634(w_eco4634, b[3], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4635(w_eco4635, b[3], a[1], !b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4636(w_eco4636, a[1], !b[1], a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4637(w_eco4637, a[1], !b[1], a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4638(w_eco4638, !a[3], b[3], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4639(w_eco4639, !a[3], b[3], !a[1], b[1], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4640(w_eco4640, b[3], !a[1], b[1], !a[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4641(w_eco4641, b[3], !a[1], b[1], !a[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4642(w_eco4642, !a[3], !a[1], b[1], !a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4643(w_eco4643, !a[3], !a[1], b[1], !a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4644(w_eco4644, !a[3], a[1], b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4645(w_eco4645, !a[3], a[1], b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4646(w_eco4646, !a[3], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4647(w_eco4647, !a[3], a[1], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4648(w_eco4648, !a[3], !a[1], !b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4649(w_eco4649, !a[3], !a[1], !b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4650(w_eco4650, !b[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4651(w_eco4651, !b[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4652(w_eco4652, !a[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4653(w_eco4653, !a[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4654(w_eco4654, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4655(w_eco4655, !a[3], !b[3], a[5], b[5], a[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4656(w_eco4656, !a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4657(w_eco4657, !a[3], !b[3], a[5], b[5], a[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4658(w_eco4658, !a[3], !b[3], a[5], b[5], a[6], !a[1], b[1], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4659(w_eco4659, !a[3], !b[3], a[5], b[5], a[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4660(w_eco4660, !b[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4661(w_eco4661, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4662(w_eco4662, !b[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4663(w_eco4663, !b[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4664(w_eco4664, !b[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4665(w_eco4665, !a[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4666(w_eco4666, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4667(w_eco4667, !a[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4668(w_eco4668, !a[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4669(w_eco4669, !a[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4670(w_eco4670, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4671(w_eco4671, a[4], !b[4], a[5], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4672(w_eco4672, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4673(w_eco4673, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4674(w_eco4674, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4675(w_eco4675, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4676(w_eco4676, !a[3], !a[4], !b[4], a[5], b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4677(w_eco4677, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4678(w_eco4678, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_4679(w_eco4679, a[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4680(w_eco4680, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4681(w_eco4681, a[3], !b[3], b[4], !a[5], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4682(w_eco4682, a[3], !b[3], b[4], !a[5], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4683(w_eco4683, !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4684(w_eco4684, a[3], !b[3], b[4], !a[5], b[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4685(w_eco4685, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4686(w_eco4686, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4687(w_eco4687, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4688(w_eco4688, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4689(w_eco4689, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4690(w_eco4690, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4691(w_eco4691, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4692(w_eco4692, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4693(w_eco4693, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4694(w_eco4694, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4695(w_eco4695, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4696(w_eco4696, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4697(w_eco4697, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4698(w_eco4698, !a[3], !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4699(w_eco4699, !b[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4700(w_eco4700, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4701(w_eco4701, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4702(w_eco4702, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4703(w_eco4703, !a[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4704(w_eco4704, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4705(w_eco4705, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4706(w_eco4706, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4707(w_eco4707, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4708(w_eco4708, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4709(w_eco4709, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4710(w_eco4710, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4711(w_eco4711, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4712(w_eco4712, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4713(w_eco4713, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4714(w_eco4714, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4715(w_eco4715, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4716(w_eco4716, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4717(w_eco4717, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4718(w_eco4718, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4719(w_eco4719, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4720(w_eco4720, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4721(w_eco4721, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4722(w_eco4722, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4723(w_eco4723, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4724(w_eco4724, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4725(w_eco4725, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4726(w_eco4726, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4727(w_eco4727, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4728(w_eco4728, !b[3], a[6], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4729(w_eco4729, !b[3], a[6], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4730(w_eco4730, !a[3], a[6], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4731(w_eco4731, !a[3], a[6], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4732(w_eco4732, !a[3], !b[3], a[6], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4733(w_eco4733, !a[3], !b[3], a[6], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4734(w_eco4734, !a[3], !b[3], a[6], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4735(w_eco4735, !a[3], !b[3], a[6], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4736(w_eco4736, !a[3], !b[3], a[6], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4737(w_eco4737, !a[3], !b[3], a[6], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4738(w_eco4738, !b[3], a[6], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4739(w_eco4739, !b[3], a[6], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4740(w_eco4740, !b[3], a[6], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4741(w_eco4741, !b[3], a[6], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4742(w_eco4742, !b[3], a[6], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4743(w_eco4743, !a[3], a[6], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4744(w_eco4744, !a[3], a[6], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4745(w_eco4745, !a[3], a[6], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4746(w_eco4746, !a[3], a[6], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4747(w_eco4747, !a[3], a[6], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4748(w_eco4748, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4749(w_eco4749, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], !b[0], op[0], !op[1]);
	and _ECO_4750(w_eco4750, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4751(w_eco4751, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4752(w_eco4752, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4753(w_eco4753, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_4754(w_eco4754, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4755(w_eco4755, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4756(w_eco4756, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4757(w_eco4757, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4758(w_eco4758, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4759(w_eco4759, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4760(w_eco4760, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4761(w_eco4761, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4762(w_eco4762, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4763(w_eco4763, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4764(w_eco4764, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4765(w_eco4765, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4766(w_eco4766, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4767(w_eco4767, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4768(w_eco4768, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4769(w_eco4769, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4770(w_eco4770, a[5], !b[5], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4771(w_eco4771, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4772(w_eco4772, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4773(w_eco4773, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4774(w_eco4774, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4775(w_eco4775, !a[3], a[4], b[4], !a[5], !b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4776(w_eco4776, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4777(w_eco4777, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_4778(w_eco4778, a[4], !b[4], !b[5], !a[1], b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4779(w_eco4779, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4780(w_eco4780, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4781(w_eco4781, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4782(w_eco4782, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], b[1], b[2], a[0], op[0], !op[1]);
	and _ECO_4783(w_eco4783, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4784(w_eco4784, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[1], !b[1], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4785(w_eco4785, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], a[0], op[0], !op[1]);
	and _ECO_4786(w_eco4786, a[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4787(w_eco4787, a[3], !b[3], !a[6], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4788(w_eco4788, a[3], !b[3], !a[6], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4789(w_eco4789, a[3], !b[3], !a[6], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4790(w_eco4790, !b[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4791(w_eco4791, a[3], !b[3], !a[6], b[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4792(w_eco4792, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4793(w_eco4793, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4794(w_eco4794, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4795(w_eco4795, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4796(w_eco4796, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4797(w_eco4797, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4798(w_eco4798, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4799(w_eco4799, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4800(w_eco4800, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4801(w_eco4801, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4802(w_eco4802, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4803(w_eco4803, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4804(w_eco4804, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4805(w_eco4805, !a[3], !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4806(w_eco4806, !b[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4807(w_eco4807, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4808(w_eco4808, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4809(w_eco4809, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4810(w_eco4810, !a[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4811(w_eco4811, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4812(w_eco4812, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4813(w_eco4813, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4814(w_eco4814, a[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4815(w_eco4815, a[3], !a[4], b[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4816(w_eco4816, a[3], !a[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4817(w_eco4817, !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4818(w_eco4818, !b[3], !a[4], b[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4819(w_eco4819, !b[3], !a[4], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4820(w_eco4820, a[3], !b[3], !a[4], b[5], b[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4821(w_eco4821, !b[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4822(w_eco4822, !b[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4823(w_eco4823, !b[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4824(w_eco4824, !a[3], a[5], b[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4825(w_eco4825, !a[3], a[5], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4826(w_eco4826, !a[3], a[5], b[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4827(w_eco4827, !b[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4828(w_eco4828, !a[3], a[5], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4829(w_eco4829, b[3], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4830(w_eco4830, b[3], a[1], !b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4831(w_eco4831, b[3], !a[1], b[1], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4832(w_eco4832, b[3], !a[1], b[1], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4833(w_eco4833, a[1], !b[1], a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4834(w_eco4834, a[1], !b[1], a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4835(w_eco4835, !a[3], b[3], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4836(w_eco4836, !a[3], b[3], !a[1], b[1], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4837(w_eco4837, !a[3], b[3], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4838(w_eco4838, !a[3], b[3], a[1], b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4839(w_eco4839, !a[3], b[3], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4840(w_eco4840, !a[3], b[3], !a[1], !b[1], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4841(w_eco4841, !a[3], !a[1], b[1], b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4842(w_eco4842, !a[3], !a[1], b[1], b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4843(w_eco4843, b[3], !a[1], b[1], !a[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4844(w_eco4844, b[3], !a[1], b[1], !a[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4845(w_eco4845, b[3], a[1], b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4846(w_eco4846, b[3], a[1], b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4847(w_eco4847, b[3], !a[1], !b[1], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4848(w_eco4848, b[3], !a[1], !b[1], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4849(w_eco4849, a[1], !b[1], !b[2], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4850(w_eco4850, a[1], !b[1], !b[2], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_4851(w_eco4851, !b[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4852(w_eco4852, !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4853(w_eco4853, !b[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4854(w_eco4854, !b[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4855(w_eco4855, !b[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4856(w_eco4856, !a[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4857(w_eco4857, !a[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4858(w_eco4858, !a[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4859(w_eco4859, !a[3], b[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4860(w_eco4860, !a[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4861(w_eco4861, !a[3], !b[3], a[5], b[5], a[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4862(w_eco4862, !a[3], !b[3], a[5], b[5], a[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4863(w_eco4863, !a[3], !b[3], a[5], b[5], a[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4864(w_eco4864, !a[3], !b[3], a[5], b[5], a[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4865(w_eco4865, !b[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4866(w_eco4866, !b[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4867(w_eco4867, !b[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4868(w_eco4868, !b[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4869(w_eco4869, !a[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4870(w_eco4870, !a[3], a[5], b[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4871(w_eco4871, !a[3], a[5], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4872(w_eco4872, !a[3], a[5], b[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4873(w_eco4873, a[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4874(w_eco4874, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4875(w_eco4875, a[3], !b[3], !a[4], b[5], !a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4876(w_eco4876, a[3], !b[3], !a[4], b[5], !a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4877(w_eco4877, !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4878(w_eco4878, a[3], !b[3], !a[4], b[5], !a[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4879(w_eco4879, a[4], !b[4], a[5], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4880(w_eco4880, a[4], !b[4], a[5], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4881(w_eco4881, a[4], !b[4], a[5], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4882(w_eco4882, a[4], !b[4], a[5], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4883(w_eco4883, a[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4884(w_eco4884, a[3], b[4], !a[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4885(w_eco4885, a[3], b[4], !a[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4886(w_eco4886, !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4887(w_eco4887, !b[3], b[4], !a[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4888(w_eco4888, !b[3], b[4], !a[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4889(w_eco4889, a[3], !b[3], b[4], !a[5], b[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4890(w_eco4890, !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4891(w_eco4891, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4892(w_eco4892, !b[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4893(w_eco4893, !a[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4894(w_eco4894, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4895(w_eco4895, !a[3], a[4], b[4], b[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4896(w_eco4896, !b[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4897(w_eco4897, !a[3], a[4], b[4], b[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4898(w_eco4898, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4899(w_eco4899, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4900(w_eco4900, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4901(w_eco4901, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_4902(w_eco4902, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4903(w_eco4903, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4904(w_eco4904, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4905(w_eco4905, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4906(w_eco4906, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4907(w_eco4907, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4908(w_eco4908, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4909(w_eco4909, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4910(w_eco4910, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4911(w_eco4911, !a[3], !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4912(w_eco4912, !b[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4913(w_eco4913, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4914(w_eco4914, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4915(w_eco4915, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4916(w_eco4916, !a[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4917(w_eco4917, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4918(w_eco4918, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4919(w_eco4919, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4920(w_eco4920, a[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4921(w_eco4921, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4922(w_eco4922, a[3], !b[3], b[4], !a[5], !a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4923(w_eco4923, a[3], !b[3], b[4], !a[5], !a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4924(w_eco4924, !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4925(w_eco4925, a[3], !b[3], b[4], !a[5], !a[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4926(w_eco4926, !b[3], a[6], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4927(w_eco4927, !b[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4928(w_eco4928, !b[3], a[6], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4929(w_eco4929, !b[3], a[6], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4930(w_eco4930, !b[3], a[6], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4931(w_eco4931, !a[3], a[6], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4932(w_eco4932, !a[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4933(w_eco4933, !a[3], a[6], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4934(w_eco4934, !a[3], a[6], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4935(w_eco4935, !a[3], a[6], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4936(w_eco4936, !a[3], !b[3], a[6], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4937(w_eco4937, !a[3], !b[3], a[6], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4938(w_eco4938, !a[3], !b[3], a[6], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4939(w_eco4939, !a[3], !b[3], a[6], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4940(w_eco4940, !b[3], a[6], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4941(w_eco4941, !b[3], a[6], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4942(w_eco4942, !b[3], a[6], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4943(w_eco4943, !b[3], a[6], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4944(w_eco4944, !a[3], a[6], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4945(w_eco4945, !a[3], a[6], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4946(w_eco4946, !a[3], a[6], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4947(w_eco4947, !a[3], a[6], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4948(w_eco4948, a[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4949(w_eco4949, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4950(w_eco4950, a[3], !b[3], !a[5], b[5], b[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4951(w_eco4951, a[3], !b[3], !a[5], b[5], b[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4952(w_eco4952, !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4953(w_eco4953, a[3], !b[3], !a[5], b[5], b[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4954(w_eco4954, a[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4955(w_eco4955, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[0], op[0], !op[1]);
	and _ECO_4956(w_eco4956, a[3], !b[3], !a[5], b[5], !a[6], a[1], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4957(w_eco4957, a[3], !b[3], !a[5], b[5], !a[6], !a[1], !b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_4958(w_eco4958, !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], !b[0], op[0], !op[1]);
	and _ECO_4959(w_eco4959, a[3], !b[3], !a[5], b[5], !a[6], a[1], !b[1], !a[2], b[2], !b[0], op[0], !op[1]);
	and _ECO_4960(w_eco4960, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4961(w_eco4961, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4962(w_eco4962, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4963(w_eco4963, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4964(w_eco4964, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4965(w_eco4965, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4966(w_eco4966, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4967(w_eco4967, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], !a[7], !op[0], !op[1]);
	and _ECO_4968(w_eco4968, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4969(w_eco4969, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !b[0], a[7], !b[7], !op[1]);
	and _ECO_4970(w_eco4970, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4971(w_eco4971, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4972(w_eco4972, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4973(w_eco4973, !a[3], !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4974(w_eco4974, !b[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4975(w_eco4975, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4976(w_eco4976, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4977(w_eco4977, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4978(w_eco4978, !a[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_4979(w_eco4979, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4980(w_eco4980, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !a[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4981(w_eco4981, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !a[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4982(w_eco4982, a[5], !b[5], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4983(w_eco4983, a[5], !b[5], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4984(w_eco4984, a[5], !b[5], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4985(w_eco4985, a[5], !b[5], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4986(w_eco4986, a[4], !b[4], !b[5], !a[1], b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4987(w_eco4987, a[4], !b[4], !b[5], a[1], b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4988(w_eco4988, a[4], !b[4], !b[5], !a[1], !b[1], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4989(w_eco4989, a[4], !b[4], !b[5], a[1], !b[1], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_4990(w_eco4990, a[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4991(w_eco4991, a[3], !a[6], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4992(w_eco4992, a[3], !a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4993(w_eco4993, !b[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_4994(w_eco4994, !b[3], !a[6], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4995(w_eco4995, !b[3], !a[6], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_4996(w_eco4996, a[3], !b[3], !a[6], b[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_4997(w_eco4997, !b[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_4998(w_eco4998, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_4999(w_eco4999, !b[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5000(w_eco5000, !a[3], a[4], b[4], a[5], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5001(w_eco5001, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5002(w_eco5002, !a[3], a[4], b[4], a[5], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5003(w_eco5003, !b[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5004(w_eco5004, !a[3], a[4], b[4], a[5], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5005(w_eco5005, !b[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5006(w_eco5006, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5007(w_eco5007, !b[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5008(w_eco5008, !a[3], a[4], b[4], a[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5009(w_eco5009, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5010(w_eco5010, !a[3], a[4], b[4], a[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5011(w_eco5011, !b[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5012(w_eco5012, !a[3], a[4], b[4], a[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5013(w_eco5013, b[3], !a[1], b[1], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5014(w_eco5014, b[3], !a[1], b[1], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5015(w_eco5015, b[3], a[1], b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5016(w_eco5016, b[3], a[1], b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5017(w_eco5017, b[3], !a[1], !b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5018(w_eco5018, b[3], !a[1], !b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5019(w_eco5019, !a[3], !a[1], b[1], b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5020(w_eco5020, !a[3], !a[1], b[1], b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5021(w_eco5021, !a[3], a[1], b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5022(w_eco5022, !a[3], a[1], b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5023(w_eco5023, !a[3], !a[1], !b[1], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5024(w_eco5024, !a[3], !a[1], !b[1], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5025(w_eco5025, a[1], !b[1], !b[2], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5026(w_eco5026, a[1], !b[1], !b[2], a[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5027(w_eco5027, !b[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5028(w_eco5028, !b[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5029(w_eco5029, !b[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5030(w_eco5030, !a[3], a[5], b[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5031(w_eco5031, !a[3], a[5], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5032(w_eco5032, !a[3], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5033(w_eco5033, !b[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5034(w_eco5034, !a[3], a[5], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5035(w_eco5035, a[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5036(w_eco5036, a[3], !a[4], b[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5037(w_eco5037, a[3], !a[4], b[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5038(w_eco5038, !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5039(w_eco5039, !b[3], !a[4], b[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5040(w_eco5040, !b[3], !a[4], b[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5041(w_eco5041, a[3], !b[3], !a[4], b[5], !a[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_5042(w_eco5042, a[4], !b[4], a[5], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5043(w_eco5043, !b[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5044(w_eco5044, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5045(w_eco5045, !b[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5046(w_eco5046, !a[3], a[4], b[4], b[5], a[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5047(w_eco5047, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5048(w_eco5048, !a[3], a[4], b[4], b[5], a[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5049(w_eco5049, !b[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5050(w_eco5050, !a[3], a[4], b[4], b[5], a[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5051(w_eco5051, a[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5052(w_eco5052, a[3], b[4], !a[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5053(w_eco5053, a[3], b[4], !a[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5054(w_eco5054, !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5055(w_eco5055, !b[3], b[4], !a[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5056(w_eco5056, !b[3], b[4], !a[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5057(w_eco5057, a[3], !b[3], b[4], !a[5], !a[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_5058(w_eco5058, !b[3], a[6], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5059(w_eco5059, !b[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5060(w_eco5060, !b[3], a[6], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5061(w_eco5061, !a[3], a[6], b[6], !a[1], b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5062(w_eco5062, !a[3], a[6], b[6], !a[1], !b[1], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5063(w_eco5063, !a[3], a[6], b[6], a[1], !b[1], !b[2], !a[0], !b[7], !op[0], !op[1]);
	and _ECO_5064(w_eco5064, !b[3], a[6], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5065(w_eco5065, !a[3], a[6], b[6], a[1], b[1], !a[2], !b[2], a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5066(w_eco5066, a[5], !b[5], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5067(w_eco5067, a[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5068(w_eco5068, a[3], !a[5], b[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5069(w_eco5069, a[3], !a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5070(w_eco5070, !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5071(w_eco5071, !b[3], !a[5], b[5], b[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5072(w_eco5072, !b[3], !a[5], b[5], b[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5073(w_eco5073, a[3], !b[3], !a[5], b[5], b[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_5074(w_eco5074, a[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5075(w_eco5075, a[3], !a[5], b[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5076(w_eco5076, a[3], !a[5], b[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5077(w_eco5077, !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], op[0], !op[1]);
	and _ECO_5078(w_eco5078, !b[3], !a[5], b[5], !a[6], a[1], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5079(w_eco5079, !b[3], !a[5], b[5], !a[6], !a[1], !b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5080(w_eco5080, a[3], !b[3], !a[5], b[5], !a[6], a[1], !b[1], !a[2], b[2], a[0], op[0], !op[1]);
	and _ECO_5081(w_eco5081, a[4], !b[4], !b[5], a[1], !b[1], a[0], a[7], !b[7], op[0], !op[1]);
	or _ECO_5082(w_eco5082, w_eco4286, w_eco4287, w_eco4288, w_eco4289, w_eco4290, w_eco4291, w_eco4292, w_eco4293, w_eco4294, w_eco4295, w_eco4296, w_eco4297, w_eco4298, w_eco4299, w_eco4300, w_eco4301, w_eco4302, w_eco4303, w_eco4304, w_eco4305, w_eco4306, w_eco4307, w_eco4308, w_eco4309, w_eco4310, w_eco4311, w_eco4312, w_eco4313, w_eco4314, w_eco4315, w_eco4316, w_eco4317, w_eco4318, w_eco4319, w_eco4320, w_eco4321, w_eco4322, w_eco4323, w_eco4324, w_eco4325, w_eco4326, w_eco4327, w_eco4328, w_eco4329, w_eco4330, w_eco4331, w_eco4332, w_eco4333, w_eco4334, w_eco4335, w_eco4336, w_eco4337, w_eco4338, w_eco4339, w_eco4340, w_eco4341, w_eco4342, w_eco4343, w_eco4344, w_eco4345, w_eco4346, w_eco4347, w_eco4348, w_eco4349, w_eco4350, w_eco4351, w_eco4352, w_eco4353, w_eco4354, w_eco4355, w_eco4356, w_eco4357, w_eco4358, w_eco4359, w_eco4360, w_eco4361, w_eco4362, w_eco4363, w_eco4364, w_eco4365, w_eco4366, w_eco4367, w_eco4368, w_eco4369, w_eco4370, w_eco4371, w_eco4372, w_eco4373, w_eco4374, w_eco4375, w_eco4376, w_eco4377, w_eco4378, w_eco4379, w_eco4380, w_eco4381, w_eco4382, w_eco4383, w_eco4384, w_eco4385, w_eco4386, w_eco4387, w_eco4388, w_eco4389, w_eco4390, w_eco4391, w_eco4392, w_eco4393, w_eco4394, w_eco4395, w_eco4396, w_eco4397, w_eco4398, w_eco4399, w_eco4400, w_eco4401, w_eco4402, w_eco4403, w_eco4404, w_eco4405, w_eco4406, w_eco4407, w_eco4408, w_eco4409, w_eco4410, w_eco4411, w_eco4412, w_eco4413, w_eco4414, w_eco4415, w_eco4416, w_eco4417, w_eco4418, w_eco4419, w_eco4420, w_eco4421, w_eco4422, w_eco4423, w_eco4424, w_eco4425, w_eco4426, w_eco4427, w_eco4428, w_eco4429, w_eco4430, w_eco4431, w_eco4432, w_eco4433, w_eco4434, w_eco4435, w_eco4436, w_eco4437, w_eco4438, w_eco4439, w_eco4440, w_eco4441, w_eco4442, w_eco4443, w_eco4444, w_eco4445, w_eco4446, w_eco4447, w_eco4448, w_eco4449, w_eco4450, w_eco4451, w_eco4452, w_eco4453, w_eco4454, w_eco4455, w_eco4456, w_eco4457, w_eco4458, w_eco4459, w_eco4460, w_eco4461, w_eco4462, w_eco4463, w_eco4464, w_eco4465, w_eco4466, w_eco4467, w_eco4468, w_eco4469, w_eco4470, w_eco4471, w_eco4472, w_eco4473, w_eco4474, w_eco4475, w_eco4476, w_eco4477, w_eco4478, w_eco4479, w_eco4480, w_eco4481, w_eco4482, w_eco4483, w_eco4484, w_eco4485, w_eco4486, w_eco4487, w_eco4488, w_eco4489, w_eco4490, w_eco4491, w_eco4492, w_eco4493, w_eco4494, w_eco4495, w_eco4496, w_eco4497, w_eco4498, w_eco4499, w_eco4500, w_eco4501, w_eco4502, w_eco4503, w_eco4504, w_eco4505, w_eco4506, w_eco4507, w_eco4508, w_eco4509, w_eco4510, w_eco4511, w_eco4512, w_eco4513, w_eco4514, w_eco4515, w_eco4516, w_eco4517, w_eco4518, w_eco4519, w_eco4520, w_eco4521, w_eco4522, w_eco4523, w_eco4524, w_eco4525, w_eco4526, w_eco4527, w_eco4528, w_eco4529, w_eco4530, w_eco4531, w_eco4532, w_eco4533, w_eco4534, w_eco4535, w_eco4536, w_eco4537, w_eco4538, w_eco4539, w_eco4540, w_eco4541, w_eco4542, w_eco4543, w_eco4544, w_eco4545, w_eco4546, w_eco4547, w_eco4548, w_eco4549, w_eco4550, w_eco4551, w_eco4552, w_eco4553, w_eco4554, w_eco4555, w_eco4556, w_eco4557, w_eco4558, w_eco4559, w_eco4560, w_eco4561, w_eco4562, w_eco4563, w_eco4564, w_eco4565, w_eco4566, w_eco4567, w_eco4568, w_eco4569, w_eco4570, w_eco4571, w_eco4572, w_eco4573, w_eco4574, w_eco4575, w_eco4576, w_eco4577, w_eco4578, w_eco4579, w_eco4580, w_eco4581, w_eco4582, w_eco4583, w_eco4584, w_eco4585, w_eco4586, w_eco4587, w_eco4588, w_eco4589, w_eco4590, w_eco4591, w_eco4592, w_eco4593, w_eco4594, w_eco4595, w_eco4596, w_eco4597, w_eco4598, w_eco4599, w_eco4600, w_eco4601, w_eco4602, w_eco4603, w_eco4604, w_eco4605, w_eco4606, w_eco4607, w_eco4608, w_eco4609, w_eco4610, w_eco4611, w_eco4612, w_eco4613, w_eco4614, w_eco4615, w_eco4616, w_eco4617, w_eco4618, w_eco4619, w_eco4620, w_eco4621, w_eco4622, w_eco4623, w_eco4624, w_eco4625, w_eco4626, w_eco4627, w_eco4628, w_eco4629, w_eco4630, w_eco4631, w_eco4632, w_eco4633, w_eco4634, w_eco4635, w_eco4636, w_eco4637, w_eco4638, w_eco4639, w_eco4640, w_eco4641, w_eco4642, w_eco4643, w_eco4644, w_eco4645, w_eco4646, w_eco4647, w_eco4648, w_eco4649, w_eco4650, w_eco4651, w_eco4652, w_eco4653, w_eco4654, w_eco4655, w_eco4656, w_eco4657, w_eco4658, w_eco4659, w_eco4660, w_eco4661, w_eco4662, w_eco4663, w_eco4664, w_eco4665, w_eco4666, w_eco4667, w_eco4668, w_eco4669, w_eco4670, w_eco4671, w_eco4672, w_eco4673, w_eco4674, w_eco4675, w_eco4676, w_eco4677, w_eco4678, w_eco4679, w_eco4680, w_eco4681, w_eco4682, w_eco4683, w_eco4684, w_eco4685, w_eco4686, w_eco4687, w_eco4688, w_eco4689, w_eco4690, w_eco4691, w_eco4692, w_eco4693, w_eco4694, w_eco4695, w_eco4696, w_eco4697, w_eco4698, w_eco4699, w_eco4700, w_eco4701, w_eco4702, w_eco4703, w_eco4704, w_eco4705, w_eco4706, w_eco4707, w_eco4708, w_eco4709, w_eco4710, w_eco4711, w_eco4712, w_eco4713, w_eco4714, w_eco4715, w_eco4716, w_eco4717, w_eco4718, w_eco4719, w_eco4720, w_eco4721, w_eco4722, w_eco4723, w_eco4724, w_eco4725, w_eco4726, w_eco4727, w_eco4728, w_eco4729, w_eco4730, w_eco4731, w_eco4732, w_eco4733, w_eco4734, w_eco4735, w_eco4736, w_eco4737, w_eco4738, w_eco4739, w_eco4740, w_eco4741, w_eco4742, w_eco4743, w_eco4744, w_eco4745, w_eco4746, w_eco4747, w_eco4748, w_eco4749, w_eco4750, w_eco4751, w_eco4752, w_eco4753, w_eco4754, w_eco4755, w_eco4756, w_eco4757, w_eco4758, w_eco4759, w_eco4760, w_eco4761, w_eco4762, w_eco4763, w_eco4764, w_eco4765, w_eco4766, w_eco4767, w_eco4768, w_eco4769, w_eco4770, w_eco4771, w_eco4772, w_eco4773, w_eco4774, w_eco4775, w_eco4776, w_eco4777, w_eco4778, w_eco4779, w_eco4780, w_eco4781, w_eco4782, w_eco4783, w_eco4784, w_eco4785, w_eco4786, w_eco4787, w_eco4788, w_eco4789, w_eco4790, w_eco4791, w_eco4792, w_eco4793, w_eco4794, w_eco4795, w_eco4796, w_eco4797, w_eco4798, w_eco4799, w_eco4800, w_eco4801, w_eco4802, w_eco4803, w_eco4804, w_eco4805, w_eco4806, w_eco4807, w_eco4808, w_eco4809, w_eco4810, w_eco4811, w_eco4812, w_eco4813, w_eco4814, w_eco4815, w_eco4816, w_eco4817, w_eco4818, w_eco4819, w_eco4820, w_eco4821, w_eco4822, w_eco4823, w_eco4824, w_eco4825, w_eco4826, w_eco4827, w_eco4828, w_eco4829, w_eco4830, w_eco4831, w_eco4832, w_eco4833, w_eco4834, w_eco4835, w_eco4836, w_eco4837, w_eco4838, w_eco4839, w_eco4840, w_eco4841, w_eco4842, w_eco4843, w_eco4844, w_eco4845, w_eco4846, w_eco4847, w_eco4848, w_eco4849, w_eco4850, w_eco4851, w_eco4852, w_eco4853, w_eco4854, w_eco4855, w_eco4856, w_eco4857, w_eco4858, w_eco4859, w_eco4860, w_eco4861, w_eco4862, w_eco4863, w_eco4864, w_eco4865, w_eco4866, w_eco4867, w_eco4868, w_eco4869, w_eco4870, w_eco4871, w_eco4872, w_eco4873, w_eco4874, w_eco4875, w_eco4876, w_eco4877, w_eco4878, w_eco4879, w_eco4880, w_eco4881, w_eco4882, w_eco4883, w_eco4884, w_eco4885, w_eco4886, w_eco4887, w_eco4888, w_eco4889, w_eco4890, w_eco4891, w_eco4892, w_eco4893, w_eco4894, w_eco4895, w_eco4896, w_eco4897, w_eco4898, w_eco4899, w_eco4900, w_eco4901, w_eco4902, w_eco4903, w_eco4904, w_eco4905, w_eco4906, w_eco4907, w_eco4908, w_eco4909, w_eco4910, w_eco4911, w_eco4912, w_eco4913, w_eco4914, w_eco4915, w_eco4916, w_eco4917, w_eco4918, w_eco4919, w_eco4920, w_eco4921, w_eco4922, w_eco4923, w_eco4924, w_eco4925, w_eco4926, w_eco4927, w_eco4928, w_eco4929, w_eco4930, w_eco4931, w_eco4932, w_eco4933, w_eco4934, w_eco4935, w_eco4936, w_eco4937, w_eco4938, w_eco4939, w_eco4940, w_eco4941, w_eco4942, w_eco4943, w_eco4944, w_eco4945, w_eco4946, w_eco4947, w_eco4948, w_eco4949, w_eco4950, w_eco4951, w_eco4952, w_eco4953, w_eco4954, w_eco4955, w_eco4956, w_eco4957, w_eco4958, w_eco4959, w_eco4960, w_eco4961, w_eco4962, w_eco4963, w_eco4964, w_eco4965, w_eco4966, w_eco4967, w_eco4968, w_eco4969, w_eco4970, w_eco4971, w_eco4972, w_eco4973, w_eco4974, w_eco4975, w_eco4976, w_eco4977, w_eco4978, w_eco4979, w_eco4980, w_eco4981, w_eco4982, w_eco4983, w_eco4984, w_eco4985, w_eco4986, w_eco4987, w_eco4988, w_eco4989, w_eco4990, w_eco4991, w_eco4992, w_eco4993, w_eco4994, w_eco4995, w_eco4996, w_eco4997, w_eco4998, w_eco4999, w_eco5000, w_eco5001, w_eco5002, w_eco5003, w_eco5004, w_eco5005, w_eco5006, w_eco5007, w_eco5008, w_eco5009, w_eco5010, w_eco5011, w_eco5012, w_eco5013, w_eco5014, w_eco5015, w_eco5016, w_eco5017, w_eco5018, w_eco5019, w_eco5020, w_eco5021, w_eco5022, w_eco5023, w_eco5024, w_eco5025, w_eco5026, w_eco5027, w_eco5028, w_eco5029, w_eco5030, w_eco5031, w_eco5032, w_eco5033, w_eco5034, w_eco5035, w_eco5036, w_eco5037, w_eco5038, w_eco5039, w_eco5040, w_eco5041, w_eco5042, w_eco5043, w_eco5044, w_eco5045, w_eco5046, w_eco5047, w_eco5048, w_eco5049, w_eco5050, w_eco5051, w_eco5052, w_eco5053, w_eco5054, w_eco5055, w_eco5056, w_eco5057, w_eco5058, w_eco5059, w_eco5060, w_eco5061, w_eco5062, w_eco5063, w_eco5064, w_eco5065, w_eco5066, w_eco5067, w_eco5068, w_eco5069, w_eco5070, w_eco5071, w_eco5072, w_eco5073, w_eco5074, w_eco5075, w_eco5076, w_eco5077, w_eco5078, w_eco5079, w_eco5080, w_eco5081);
	xor _ECO_out8(y[1], sub_wire8, w_eco5082);
	and _ECO_5083(w_eco5083, a[4], b[4], a[5], b[5], a[6], b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5084(w_eco5084, a[4], b[4], a[5], b[5], a[6], b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5085(w_eco5085, a[4], b[4], a[5], b[5], !a[6], !b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5086(w_eco5086, a[4], b[4], a[5], b[5], !a[6], !b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5087(w_eco5087, !a[4], !b[4], a[5], b[5], a[6], b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5088(w_eco5088, !a[4], !b[4], a[5], b[5], a[6], b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5089(w_eco5089, !a[4], !b[4], a[5], b[5], !a[6], !b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5090(w_eco5090, !a[4], !b[4], a[5], b[5], !a[6], !b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5091(w_eco5091, a[4], b[4], !a[5], !b[5], a[6], b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5092(w_eco5092, a[4], b[4], !a[5], !b[5], a[6], b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5093(w_eco5093, a[4], b[4], !a[5], !b[5], !a[6], !b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5094(w_eco5094, a[4], b[4], !a[5], !b[5], !a[6], !b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5095(w_eco5095, !a[4], !b[4], !a[5], !b[5], a[6], b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5096(w_eco5096, !a[4], !b[4], !a[5], !b[5], a[6], b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5097(w_eco5097, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5098(w_eco5098, !a[4], !b[4], !a[5], !b[5], !a[6], !b[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5099(w_eco5099, !a[4], !b[4], a[6], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5100(w_eco5100, !a[4], !b[4], a[6], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5101(w_eco5101, !a[4], !b[4], a[5], b[5], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5102(w_eco5102, !a[4], !b[4], a[5], b[5], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5103(w_eco5103, !a[4], !b[4], a[5], b[5], a[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5104(w_eco5104, !a[4], !b[4], a[5], b[5], a[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5105(w_eco5105, !a[5], !b[5], a[6], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5106(w_eco5106, !a[5], !b[5], a[6], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5107(w_eco5107, !a[3], a[4], b[4], a[5], b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5108(w_eco5108, !a[3], a[4], b[4], a[5], b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5109(w_eco5109, b[6], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5110(w_eco5110, b[6], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5111(w_eco5111, b[6], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5112(w_eco5112, b[6], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5113(w_eco5113, !a[6], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5114(w_eco5114, !a[6], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5115(w_eco5115, !a[6], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5116(w_eco5116, !a[6], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5117(w_eco5117, !a[4], !b[4], a[6], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5118(w_eco5118, !a[4], !b[4], a[6], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5119(w_eco5119, !a[4], !b[4], a[5], b[5], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5120(w_eco5120, !a[4], !b[4], a[5], b[5], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5121(w_eco5121, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5122(w_eco5122, !a[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5123(w_eco5123, !a[4], !b[4], a[5], b[5], a[6], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5124(w_eco5124, !a[4], !b[4], a[5], b[5], a[6], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5125(w_eco5125, !a[5], !b[5], a[6], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5126(w_eco5126, !a[5], !b[5], a[6], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5127(w_eco5127, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5128(w_eco5128, !a[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5129(w_eco5129, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5130(w_eco5130, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5131(w_eco5131, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5132(w_eco5132, !a[3], b[3], a[4], b[4], a[5], b[5], a[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5133(w_eco5133, b[3], a[4], b[4], a[5], b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5134(w_eco5134, b[3], a[4], b[4], a[5], b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5135(w_eco5135, !a[3], !b[3], a[5], b[5], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5136(w_eco5136, !a[3], !b[3], a[5], b[5], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5137(w_eco5137, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5138(w_eco5138, !a[3], b[3], !a[4], !b[4], a[5], b[5], a[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5139(w_eco5139, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5140(w_eco5140, b[3], !a[4], !b[4], a[5], b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5141(w_eco5141, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5142(w_eco5142, !a[3], !b[3], a[4], b[4], b[5], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5143(w_eco5143, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5144(w_eco5144, !a[3], b[3], a[4], b[4], !a[5], !b[5], a[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5145(w_eco5145, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5146(w_eco5146, b[3], a[4], b[4], !a[5], !b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5147(w_eco5147, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[0], b[0], op[0], !op[1]);
	and _ECO_5148(w_eco5148, !a[3], b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[0], !b[0], op[0], !op[1]);
	and _ECO_5149(w_eco5149, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5150(w_eco5150, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5151(w_eco5151, b[3], a[4], b[4], a[5], b[5], a[6], !b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5152(w_eco5152, a[4], b[4], a[5], b[5], a[6], !b[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5153(w_eco5153, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5154(w_eco5154, !a[3], !b[3], a[4], b[4], a[5], a[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5155(w_eco5155, !a[3], !b[3], a[5], b[5], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5156(w_eco5156, !a[3], !b[3], a[5], b[5], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5157(w_eco5157, !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5158(w_eco5158, !b[3], a[5], b[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5159(w_eco5159, !a[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5160(w_eco5160, !a[3], a[5], b[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5161(w_eco5161, !a[3], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5162(w_eco5162, !a[3], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5163(w_eco5163, !a[3], !a[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5164(w_eco5164, !a[3], !a[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5165(w_eco5165, !a[3], !b[3], a[5], b[5], a[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5166(w_eco5166, !a[3], !b[3], a[5], b[5], a[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5167(w_eco5167, b[3], !a[4], !b[4], a[5], b[5], a[6], !b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5168(w_eco5168, !a[4], !b[4], a[5], b[5], a[6], !b[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5169(w_eco5169, !a[3], !b[3], a[4], b[4], b[5], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5170(w_eco5170, !a[3], !b[3], a[4], b[4], b[5], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5171(w_eco5171, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5172(w_eco5172, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5173(w_eco5173, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5174(w_eco5174, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5175(w_eco5175, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5176(w_eco5176, !a[3], !b[3], a[4], b[4], b[5], a[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5177(w_eco5177, !a[3], !b[3], a[6], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5178(w_eco5178, !a[3], !b[3], a[6], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5179(w_eco5179, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5180(w_eco5180, !a[3], !b[3], a[4], b[4], a[5], b[6], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5181(w_eco5181, b[3], a[4], b[4], !a[5], !b[5], a[6], !b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5182(w_eco5182, a[4], b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5183(w_eco5183, b[3], !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5184(w_eco5184, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5185(w_eco5185, b[3], a[4], b[4], a[5], b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5186(w_eco5186, b[3], a[4], b[4], a[5], b[5], a[6], a[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5187(w_eco5187, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5188(w_eco5188, a[4], b[4], a[5], b[5], a[6], a[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5189(w_eco5189, !a[3], a[4], b[4], a[5], b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5190(w_eco5190, a[4], b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5191(w_eco5191, !a[3], !b[3], a[4], b[4], a[5], a[6], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5192(w_eco5192, !a[3], !b[3], a[4], b[4], a[5], a[6], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5193(w_eco5193, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5194(w_eco5194, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5195(w_eco5195, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5196(w_eco5196, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5197(w_eco5197, a[3], !b[3], !a[4], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5198(w_eco5198, !b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5199(w_eco5199, !b[3], a[5], b[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5200(w_eco5200, !a[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5201(w_eco5201, !a[3], a[5], b[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5202(w_eco5202, !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5203(w_eco5203, !b[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5204(w_eco5204, !b[3], a[5], b[5], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5205(w_eco5205, !b[3], a[5], b[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5206(w_eco5206, !a[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5207(w_eco5207, !a[3], a[5], b[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5208(w_eco5208, !a[3], a[5], b[5], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5209(w_eco5209, !a[3], a[5], b[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5210(w_eco5210, !a[3], b[3], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5211(w_eco5211, !a[3], b[3], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5212(w_eco5212, !a[3], b[3], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5213(w_eco5213, !a[3], b[3], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5214(w_eco5214, b[3], !a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5215(w_eco5215, b[3], !a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5216(w_eco5216, b[3], !a[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5217(w_eco5217, b[3], !a[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5218(w_eco5218, !a[3], !b[3], a[5], b[5], a[6], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5219(w_eco5219, !a[3], !b[3], a[5], b[5], a[6], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5220(w_eco5220, !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5221(w_eco5221, !b[3], a[5], b[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5222(w_eco5222, !a[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5223(w_eco5223, !a[3], a[5], b[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5224(w_eco5224, b[3], !a[4], !b[4], a[5], b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5225(w_eco5225, b[3], !a[4], !b[4], a[5], b[5], a[6], a[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5226(w_eco5226, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5227(w_eco5227, !a[4], !b[4], a[5], b[5], a[6], a[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5228(w_eco5228, !a[3], !a[4], !b[4], a[5], b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5229(w_eco5229, !a[4], !b[4], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5230(w_eco5230, a[3], !b[3], b[4], !a[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5231(w_eco5231, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5232(w_eco5232, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5233(w_eco5233, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5234(w_eco5234, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5235(w_eco5235, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[1]);
	and _ECO_5236(w_eco5236, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5237(w_eco5237, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !a[2], a[0], !b[0], !a[7], !op[1]);
	and _ECO_5238(w_eco5238, !b[3], a[4], b[4], b[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5239(w_eco5239, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5240(w_eco5240, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5241(w_eco5241, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5242(w_eco5242, !a[3], a[4], b[4], b[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5243(w_eco5243, !a[3], !b[3], a[4], b[4], b[5], a[6], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5244(w_eco5244, !a[3], !b[3], a[4], b[4], b[5], a[6], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5245(w_eco5245, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5246(w_eco5246, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5247(w_eco5247, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5248(w_eco5248, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5249(w_eco5249, !a[3], !b[3], a[6], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5250(w_eco5250, !a[3], !b[3], a[6], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5251(w_eco5251, !b[3], a[6], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5252(w_eco5252, !b[3], a[6], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5253(w_eco5253, !a[3], a[6], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5254(w_eco5254, !a[3], a[6], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5255(w_eco5255, !a[3], !b[3], a[4], b[4], a[5], b[6], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5256(w_eco5256, !a[3], !b[3], a[4], b[4], a[5], b[6], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5257(w_eco5257, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5258(w_eco5258, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5259(w_eco5259, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5260(w_eco5260, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5261(w_eco5261, b[3], a[4], b[4], !a[5], !b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5262(w_eco5262, b[3], a[4], b[4], !a[5], !b[5], a[6], a[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5263(w_eco5263, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5264(w_eco5264, a[4], b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5265(w_eco5265, !a[3], a[4], b[4], !a[5], !b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5266(w_eco5266, a[4], b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5267(w_eco5267, b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5268(w_eco5268, b[3], !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5269(w_eco5269, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], a[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5270(w_eco5270, !a[4], !b[4], !a[5], !b[5], a[6], a[1], a[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5271(w_eco5271, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5272(w_eco5272, !a[4], !b[4], !a[5], !b[5], a[6], !b[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5273(w_eco5273, a[3], !b[3], !a[6], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5274(w_eco5274, b[3], a[4], b[4], a[5], b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5275(w_eco5275, !a[3], a[4], b[4], a[5], b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5276(w_eco5276, a[4], b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5277(w_eco5277, a[4], b[4], a[5], b[5], a[6], a[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5278(w_eco5278, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5279(w_eco5279, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5280(w_eco5280, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5281(w_eco5281, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5282(w_eco5282, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5283(w_eco5283, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5284(w_eco5284, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5285(w_eco5285, !b[3], a[4], b[4], a[5], a[6], !b[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5286(w_eco5286, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5287(w_eco5287, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5288(w_eco5288, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5289(w_eco5289, !a[3], a[4], b[4], a[5], a[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5290(w_eco5290, a[3], !a[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5291(w_eco5291, a[3], !b[3], !a[4], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5292(w_eco5292, a[3], !b[3], !a[4], b[5], b[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5293(w_eco5293, !b[3], !a[4], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5294(w_eco5294, a[3], !b[3], !a[4], b[5], b[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5295(w_eco5295, !b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5296(w_eco5296, !b[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5297(w_eco5297, !b[3], a[5], b[5], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5298(w_eco5298, !b[3], a[5], b[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5299(w_eco5299, !a[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5300(w_eco5300, !a[3], a[5], b[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5301(w_eco5301, !a[3], a[5], b[5], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5302(w_eco5302, !a[3], a[5], b[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5303(w_eco5303, !b[3], a[5], b[5], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5304(w_eco5304, !b[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5305(w_eco5305, !b[3], a[5], b[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5306(w_eco5306, !b[3], a[5], b[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5307(w_eco5307, !a[3], a[5], b[5], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5308(w_eco5308, !a[3], a[5], b[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5309(w_eco5309, !a[3], a[5], b[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5310(w_eco5310, !a[3], a[5], b[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5311(w_eco5311, b[3], !b[1], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5312(w_eco5312, b[3], !b[1], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5313(w_eco5313, !b[1], a[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5314(w_eco5314, !b[1], a[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5315(w_eco5315, !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5316(w_eco5316, !b[3], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5317(w_eco5317, !a[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5318(w_eco5318, !a[3], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5319(w_eco5319, !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5320(w_eco5320, !b[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5321(w_eco5321, !b[3], a[5], b[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5322(w_eco5322, !b[3], a[5], b[5], a[6], !b[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5323(w_eco5323, !a[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5324(w_eco5324, !a[3], a[5], b[5], a[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5325(w_eco5325, !a[3], a[5], b[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5326(w_eco5326, !a[3], a[5], b[5], a[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5327(w_eco5327, a[3], !b[3], !a[4], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5328(w_eco5328, a[4], !b[4], a[5], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5329(w_eco5329, b[3], !a[4], !b[4], a[5], b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5330(w_eco5330, !a[3], !a[4], !b[4], a[5], b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5331(w_eco5331, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[1], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5332(w_eco5332, !a[4], !b[4], a[5], b[5], a[6], a[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5333(w_eco5333, a[3], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5334(w_eco5334, a[3], !b[3], b[4], !a[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5335(w_eco5335, a[3], !b[3], b[4], !a[5], b[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5336(w_eco5336, !b[3], b[4], !a[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5337(w_eco5337, a[3], !b[3], b[4], !a[5], b[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5338(w_eco5338, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[1]);
	and _ECO_5339(w_eco5339, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5340(w_eco5340, a[3], !b[3], a[4], b[4], b[5], b[6], !a[1], b[1], !b[2], a[0], !b[0], !a[7], !op[1]);
	and _ECO_5341(w_eco5341, !b[3], a[4], b[4], b[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5342(w_eco5342, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5343(w_eco5343, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5344(w_eco5344, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5345(w_eco5345, !a[3], a[4], b[4], b[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5346(w_eco5346, a[3], !b[3], a[4], b[4], b[5], b[6], b[1], !a[2], !b[2], !a[0], b[0], !a[7], !op[1]);
	and _ECO_5347(w_eco5347, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5348(w_eco5348, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5349(w_eco5349, !b[3], a[4], b[4], b[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5350(w_eco5350, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5351(w_eco5351, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5352(w_eco5352, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5353(w_eco5353, !a[3], a[4], b[4], b[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5354(w_eco5354, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5355(w_eco5355, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5356(w_eco5356, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5357(w_eco5357, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5358(w_eco5358, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5359(w_eco5359, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5360(w_eco5360, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5361(w_eco5361, !b[3], a[4], b[4], b[5], a[6], !b[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5362(w_eco5362, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5363(w_eco5363, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5364(w_eco5364, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5365(w_eco5365, !a[3], a[4], b[4], b[5], a[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5366(w_eco5366, a[3], !b[3], b[4], !a[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5367(w_eco5367, !b[3], a[6], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5368(w_eco5368, !b[3], a[6], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5369(w_eco5369, !a[3], a[6], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5370(w_eco5370, !a[3], a[6], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5371(w_eco5371, !b[3], a[6], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5372(w_eco5372, !b[3], a[6], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5373(w_eco5373, !b[3], a[6], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5374(w_eco5374, !b[3], a[6], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5375(w_eco5375, !a[3], a[6], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5376(w_eco5376, !a[3], a[6], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5377(w_eco5377, !a[3], a[6], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5378(w_eco5378, !a[3], a[6], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5379(w_eco5379, a[3], !b[3], !a[5], b[5], b[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5380(w_eco5380, a[3], !b[3], !a[5], b[5], !a[6], b[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5381(w_eco5381, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5382(w_eco5382, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5383(w_eco5383, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5384(w_eco5384, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5385(w_eco5385, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5386(w_eco5386, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5387(w_eco5387, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5388(w_eco5388, !b[3], a[4], b[4], a[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5389(w_eco5389, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5390(w_eco5390, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5391(w_eco5391, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5392(w_eco5392, !a[3], a[4], b[4], a[5], b[6], !b[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5393(w_eco5393, a[5], !b[5], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5394(w_eco5394, b[3], a[4], b[4], !a[5], !b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5395(w_eco5395, !a[3], a[4], b[4], !a[5], !b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5396(w_eco5396, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5397(w_eco5397, a[4], b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5398(w_eco5398, a[4], !b[4], !b[5], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5399(w_eco5399, b[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5400(w_eco5400, !a[3], !a[4], !b[4], !a[5], !b[5], a[6], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5401(w_eco5401, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[1], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5402(w_eco5402, !a[4], !b[4], !a[5], !b[5], a[6], a[1], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5403(w_eco5403, a[3], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5404(w_eco5404, !b[3], !a[6], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5405(w_eco5405, a[3], !b[3], !a[6], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5406(w_eco5406, a[3], !b[3], !a[6], b[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5407(w_eco5407, a[3], !b[3], !a[6], b[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5408(w_eco5408, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5409(w_eco5409, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5410(w_eco5410, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5411(w_eco5411, !b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5412(w_eco5412, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5413(w_eco5413, !a[3], b[3], a[4], b[4], a[5], a[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5414(w_eco5414, !a[3], a[4], b[4], a[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5415(w_eco5415, !a[3], a[4], b[4], a[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5416(w_eco5416, !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5417(w_eco5417, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5418(w_eco5418, !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5419(w_eco5419, !b[3], a[4], b[4], a[5], a[6], !a[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5420(w_eco5420, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5421(w_eco5421, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5422(w_eco5422, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5423(w_eco5423, !a[3], a[4], b[4], a[5], a[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5424(w_eco5424, a[3], !a[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5425(w_eco5425, a[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5426(w_eco5426, !b[3], !a[4], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5427(w_eco5427, !b[3], !a[4], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5428(w_eco5428, a[3], !b[3], !a[4], b[5], b[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5429(w_eco5429, !b[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5430(w_eco5430, !b[3], a[5], b[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5431(w_eco5431, !a[3], a[5], b[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5432(w_eco5432, !a[3], a[5], b[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5433(w_eco5433, !b[3], a[5], b[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5434(w_eco5434, !b[3], a[5], b[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5435(w_eco5435, !a[3], a[5], b[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5436(w_eco5436, !a[3], a[5], b[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5437(w_eco5437, b[3], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5438(w_eco5438, b[3], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5439(w_eco5439, b[3], a[1], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5440(w_eco5440, b[3], a[1], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5441(w_eco5441, a[1], !b[1], a[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5442(w_eco5442, a[1], !b[1], a[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5443(w_eco5443, a[1], a[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5444(w_eco5444, a[1], a[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5445(w_eco5445, !a[3], b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5446(w_eco5446, !a[3], b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5447(w_eco5447, !b[1], !b[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5448(w_eco5448, !b[1], !b[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5449(w_eco5449, !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5450(w_eco5450, !b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5451(w_eco5451, !b[3], a[5], b[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5452(w_eco5452, !b[3], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5453(w_eco5453, !a[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5454(w_eco5454, !a[3], b[3], a[5], b[5], a[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5455(w_eco5455, !a[3], a[5], b[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5456(w_eco5456, !a[3], a[5], b[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5457(w_eco5457, !b[3], a[5], b[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5458(w_eco5458, !b[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5459(w_eco5459, !b[3], a[5], b[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5460(w_eco5460, !b[3], a[5], b[5], a[6], !a[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5461(w_eco5461, !a[3], a[5], b[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5462(w_eco5462, !a[3], a[5], b[5], a[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5463(w_eco5463, !a[3], a[5], b[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5464(w_eco5464, !a[3], a[5], b[5], a[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5465(w_eco5465, a[3], !a[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5466(w_eco5466, a[3], !b[3], !a[4], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5467(w_eco5467, a[3], !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5468(w_eco5468, !b[3], !a[4], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5469(w_eco5469, a[3], !b[3], !a[4], b[5], !a[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5470(w_eco5470, a[4], !b[4], a[5], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5471(w_eco5471, a[3], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5472(w_eco5472, a[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5473(w_eco5473, !b[3], b[4], !a[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5474(w_eco5474, !b[3], b[4], !a[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5475(w_eco5475, a[3], !b[3], b[4], !a[5], b[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5476(w_eco5476, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5477(w_eco5477, !b[3], a[4], b[4], b[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5478(w_eco5478, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5479(w_eco5479, !a[3], a[4], b[4], b[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5480(w_eco5480, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5481(w_eco5481, !b[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5482(w_eco5482, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5483(w_eco5483, !a[3], a[4], b[4], b[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5484(w_eco5484, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5485(w_eco5485, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5486(w_eco5486, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5487(w_eco5487, !b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5488(w_eco5488, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5489(w_eco5489, !a[3], b[3], a[4], b[4], b[5], a[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5490(w_eco5490, !a[3], a[4], b[4], b[5], a[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5491(w_eco5491, !a[3], a[4], b[4], b[5], a[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5492(w_eco5492, !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5493(w_eco5493, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5494(w_eco5494, !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5495(w_eco5495, !b[3], a[4], b[4], b[5], a[6], !a[1], !a[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5496(w_eco5496, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5497(w_eco5497, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5498(w_eco5498, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5499(w_eco5499, !a[3], a[4], b[4], b[5], a[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5500(w_eco5500, a[3], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5501(w_eco5501, a[3], !b[3], b[4], !a[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5502(w_eco5502, a[3], !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5503(w_eco5503, !b[3], b[4], !a[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5504(w_eco5504, a[3], !b[3], b[4], !a[5], !a[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5505(w_eco5505, !b[3], a[6], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5506(w_eco5506, !b[3], a[6], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5507(w_eco5507, !b[3], a[6], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5508(w_eco5508, !b[3], a[6], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5509(w_eco5509, !a[3], a[6], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5510(w_eco5510, !a[3], a[6], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5511(w_eco5511, !a[3], a[6], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5512(w_eco5512, !a[3], a[6], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5513(w_eco5513, !b[3], a[6], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5514(w_eco5514, !b[3], a[6], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5515(w_eco5515, !b[3], a[6], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5516(w_eco5516, !b[3], a[6], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5517(w_eco5517, !a[3], a[6], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5518(w_eco5518, !a[3], a[6], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5519(w_eco5519, !a[3], a[6], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5520(w_eco5520, !a[3], a[6], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5521(w_eco5521, a[3], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5522(w_eco5522, a[3], !b[3], !a[5], b[5], b[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5523(w_eco5523, a[3], !b[3], !a[5], b[5], b[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5524(w_eco5524, !b[3], !a[5], b[5], b[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5525(w_eco5525, a[3], !b[3], !a[5], b[5], b[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5526(w_eco5526, a[3], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5527(w_eco5527, a[3], !b[3], !a[5], b[5], !a[6], !a[1], !a[0], b[0], op[0], !op[1]);
	and _ECO_5528(w_eco5528, a[3], !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[0], !b[0], op[0], !op[1]);
	and _ECO_5529(w_eco5529, !b[3], !a[5], b[5], !a[6], b[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5530(w_eco5530, a[3], !b[3], !a[5], b[5], !a[6], !a[2], b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5531(w_eco5531, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5532(w_eco5532, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5533(w_eco5533, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5534(w_eco5534, !b[3], a[4], b[4], a[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5535(w_eco5535, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5536(w_eco5536, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5537(w_eco5537, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5538(w_eco5538, !a[3], a[4], b[4], a[5], b[6], !b[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5539(w_eco5539, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5540(w_eco5540, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5541(w_eco5541, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5542(w_eco5542, !b[3], a[4], b[4], a[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5543(w_eco5543, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[0], b[0], !a[7], !op[0], !op[1]);
	and _ECO_5544(w_eco5544, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5545(w_eco5545, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[0], !b[0], !a[7], !op[0], !op[1]);
	and _ECO_5546(w_eco5546, !a[3], a[4], b[4], a[5], b[6], !a[1], !a[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5547(w_eco5547, a[5], !b[5], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5548(w_eco5548, a[4], !b[4], !b[5], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5549(w_eco5549, a[3], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5550(w_eco5550, a[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5551(w_eco5551, !b[3], !a[6], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5552(w_eco5552, !b[3], !a[6], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5553(w_eco5553, a[3], !b[3], !a[6], b[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5554(w_eco5554, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5555(w_eco5555, !b[3], a[4], b[4], a[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5556(w_eco5556, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5557(w_eco5557, !a[3], a[4], b[4], a[5], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5558(w_eco5558, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5559(w_eco5559, !b[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5560(w_eco5560, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5561(w_eco5561, !a[3], a[4], b[4], a[5], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5562(w_eco5562, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5563(w_eco5563, !b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5564(w_eco5564, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5565(w_eco5565, !a[3], b[3], a[4], b[4], a[5], a[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5566(w_eco5566, !b[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5567(w_eco5567, !b[3], a[4], b[4], a[5], a[6], a[1], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5568(w_eco5568, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5569(w_eco5569, !a[3], a[4], b[4], a[5], a[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5570(w_eco5570, b[3], b[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5571(w_eco5571, b[3], b[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5572(w_eco5572, !a[3], b[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5573(w_eco5573, !a[3], b[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5574(w_eco5574, a[1], !b[1], !b[2], !a[0], b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5575(w_eco5575, a[1], !b[1], !b[2], !a[0], b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5576(w_eco5576, a[1], !b[2], a[0], !b[0], a[7], !b[7], op[0], !op[1]);
	and _ECO_5577(w_eco5577, a[1], !b[2], a[0], !b[0], !a[7], b[7], op[0], !op[1]);
	and _ECO_5578(w_eco5578, !b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5579(w_eco5579, !b[3], a[5], b[5], a[6], !a[1], !b[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5580(w_eco5580, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5581(w_eco5581, !a[3], b[3], a[5], b[5], a[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5582(w_eco5582, !b[3], a[5], b[5], a[6], !a[2], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5583(w_eco5583, !b[3], a[5], b[5], a[6], a[1], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5584(w_eco5584, !a[3], a[5], b[5], a[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5585(w_eco5585, !a[3], a[5], b[5], a[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5586(w_eco5586, a[3], !a[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5587(w_eco5587, a[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5588(w_eco5588, !b[3], !a[4], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5589(w_eco5589, !b[3], !a[4], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5590(w_eco5590, a[3], !b[3], !a[4], b[5], !a[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5591(w_eco5591, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5592(w_eco5592, !b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], a[0], !b[0], !b[7], !op[0], !op[1]);
	and _ECO_5593(w_eco5593, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5594(w_eco5594, !a[3], b[3], a[4], b[4], b[5], a[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5595(w_eco5595, !b[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[0], b[0], !b[7], !op[0], !op[1]);
	and _ECO_5596(w_eco5596, !b[3], a[4], b[4], b[5], a[6], a[1], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5597(w_eco5597, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5598(w_eco5598, !a[3], a[4], b[4], b[5], a[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5599(w_eco5599, a[3], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5600(w_eco5600, a[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5601(w_eco5601, !b[3], b[4], !a[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5602(w_eco5602, !b[3], b[4], !a[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5603(w_eco5603, a[3], !b[3], b[4], !a[5], !a[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5604(w_eco5604, !b[3], a[6], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5605(w_eco5605, !b[3], a[6], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5606(w_eco5606, !a[3], a[6], b[6], !a[1], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5607(w_eco5607, !a[3], a[6], b[6], !a[1], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5608(w_eco5608, !b[3], a[6], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5609(w_eco5609, !b[3], a[6], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5610(w_eco5610, !a[3], a[6], b[6], !a[2], !b[2], !a[0], b[0], a[7], !b[7], !op[1]);
	and _ECO_5611(w_eco5611, !a[3], a[6], b[6], !a[2], !b[2], a[0], !b[0], a[7], !b[7], !op[1]);
	and _ECO_5612(w_eco5612, a[3], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5613(w_eco5613, a[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5614(w_eco5614, !b[3], !a[5], b[5], b[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5615(w_eco5615, !b[3], !a[5], b[5], b[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5616(w_eco5616, a[3], !b[3], !a[5], b[5], b[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5617(w_eco5617, a[3], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5618(w_eco5618, a[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5619(w_eco5619, !b[3], !a[5], b[5], !a[6], !a[1], a[2], !b[2], !a[0], b[0], op[0], !op[1]);
	and _ECO_5620(w_eco5620, !b[3], !a[5], b[5], !a[6], !a[1], b[1], a[2], !b[2], a[0], !b[0], op[0], !op[1]);
	and _ECO_5621(w_eco5621, a[3], !b[3], !a[5], b[5], !a[6], !a[2], b[2], !a[0], b[0], op[0], !op[1]);
	or _ECO_5622(w_eco5622, w_eco5083, w_eco5084, w_eco5085, w_eco5086, w_eco5087, w_eco5088, w_eco5089, w_eco5090, w_eco5091, w_eco5092, w_eco5093, w_eco5094, w_eco5095, w_eco5096, w_eco5097, w_eco5098, w_eco5099, w_eco5100, w_eco5101, w_eco5102, w_eco5103, w_eco5104, w_eco5105, w_eco5106, w_eco5107, w_eco5108, w_eco5109, w_eco5110, w_eco5111, w_eco5112, w_eco5113, w_eco5114, w_eco5115, w_eco5116, w_eco5117, w_eco5118, w_eco5119, w_eco5120, w_eco5121, w_eco5122, w_eco5123, w_eco5124, w_eco5125, w_eco5126, w_eco5127, w_eco5128, w_eco5129, w_eco5130, w_eco5131, w_eco5132, w_eco5133, w_eco5134, w_eco5135, w_eco5136, w_eco5137, w_eco5138, w_eco5139, w_eco5140, w_eco5141, w_eco5142, w_eco5143, w_eco5144, w_eco5145, w_eco5146, w_eco5147, w_eco5148, w_eco5149, w_eco5150, w_eco5151, w_eco5152, w_eco5153, w_eco5154, w_eco5155, w_eco5156, w_eco5157, w_eco5158, w_eco5159, w_eco5160, w_eco5161, w_eco5162, w_eco5163, w_eco5164, w_eco5165, w_eco5166, w_eco5167, w_eco5168, w_eco5169, w_eco5170, w_eco5171, w_eco5172, w_eco5173, w_eco5174, w_eco5175, w_eco5176, w_eco5177, w_eco5178, w_eco5179, w_eco5180, w_eco5181, w_eco5182, w_eco5183, w_eco5184, w_eco5185, w_eco5186, w_eco5187, w_eco5188, w_eco5189, w_eco5190, w_eco5191, w_eco5192, w_eco5193, w_eco5194, w_eco5195, w_eco5196, w_eco5197, w_eco5198, w_eco5199, w_eco5200, w_eco5201, w_eco5202, w_eco5203, w_eco5204, w_eco5205, w_eco5206, w_eco5207, w_eco5208, w_eco5209, w_eco5210, w_eco5211, w_eco5212, w_eco5213, w_eco5214, w_eco5215, w_eco5216, w_eco5217, w_eco5218, w_eco5219, w_eco5220, w_eco5221, w_eco5222, w_eco5223, w_eco5224, w_eco5225, w_eco5226, w_eco5227, w_eco5228, w_eco5229, w_eco5230, w_eco5231, w_eco5232, w_eco5233, w_eco5234, w_eco5235, w_eco5236, w_eco5237, w_eco5238, w_eco5239, w_eco5240, w_eco5241, w_eco5242, w_eco5243, w_eco5244, w_eco5245, w_eco5246, w_eco5247, w_eco5248, w_eco5249, w_eco5250, w_eco5251, w_eco5252, w_eco5253, w_eco5254, w_eco5255, w_eco5256, w_eco5257, w_eco5258, w_eco5259, w_eco5260, w_eco5261, w_eco5262, w_eco5263, w_eco5264, w_eco5265, w_eco5266, w_eco5267, w_eco5268, w_eco5269, w_eco5270, w_eco5271, w_eco5272, w_eco5273, w_eco5274, w_eco5275, w_eco5276, w_eco5277, w_eco5278, w_eco5279, w_eco5280, w_eco5281, w_eco5282, w_eco5283, w_eco5284, w_eco5285, w_eco5286, w_eco5287, w_eco5288, w_eco5289, w_eco5290, w_eco5291, w_eco5292, w_eco5293, w_eco5294, w_eco5295, w_eco5296, w_eco5297, w_eco5298, w_eco5299, w_eco5300, w_eco5301, w_eco5302, w_eco5303, w_eco5304, w_eco5305, w_eco5306, w_eco5307, w_eco5308, w_eco5309, w_eco5310, w_eco5311, w_eco5312, w_eco5313, w_eco5314, w_eco5315, w_eco5316, w_eco5317, w_eco5318, w_eco5319, w_eco5320, w_eco5321, w_eco5322, w_eco5323, w_eco5324, w_eco5325, w_eco5326, w_eco5327, w_eco5328, w_eco5329, w_eco5330, w_eco5331, w_eco5332, w_eco5333, w_eco5334, w_eco5335, w_eco5336, w_eco5337, w_eco5338, w_eco5339, w_eco5340, w_eco5341, w_eco5342, w_eco5343, w_eco5344, w_eco5345, w_eco5346, w_eco5347, w_eco5348, w_eco5349, w_eco5350, w_eco5351, w_eco5352, w_eco5353, w_eco5354, w_eco5355, w_eco5356, w_eco5357, w_eco5358, w_eco5359, w_eco5360, w_eco5361, w_eco5362, w_eco5363, w_eco5364, w_eco5365, w_eco5366, w_eco5367, w_eco5368, w_eco5369, w_eco5370, w_eco5371, w_eco5372, w_eco5373, w_eco5374, w_eco5375, w_eco5376, w_eco5377, w_eco5378, w_eco5379, w_eco5380, w_eco5381, w_eco5382, w_eco5383, w_eco5384, w_eco5385, w_eco5386, w_eco5387, w_eco5388, w_eco5389, w_eco5390, w_eco5391, w_eco5392, w_eco5393, w_eco5394, w_eco5395, w_eco5396, w_eco5397, w_eco5398, w_eco5399, w_eco5400, w_eco5401, w_eco5402, w_eco5403, w_eco5404, w_eco5405, w_eco5406, w_eco5407, w_eco5408, w_eco5409, w_eco5410, w_eco5411, w_eco5412, w_eco5413, w_eco5414, w_eco5415, w_eco5416, w_eco5417, w_eco5418, w_eco5419, w_eco5420, w_eco5421, w_eco5422, w_eco5423, w_eco5424, w_eco5425, w_eco5426, w_eco5427, w_eco5428, w_eco5429, w_eco5430, w_eco5431, w_eco5432, w_eco5433, w_eco5434, w_eco5435, w_eco5436, w_eco5437, w_eco5438, w_eco5439, w_eco5440, w_eco5441, w_eco5442, w_eco5443, w_eco5444, w_eco5445, w_eco5446, w_eco5447, w_eco5448, w_eco5449, w_eco5450, w_eco5451, w_eco5452, w_eco5453, w_eco5454, w_eco5455, w_eco5456, w_eco5457, w_eco5458, w_eco5459, w_eco5460, w_eco5461, w_eco5462, w_eco5463, w_eco5464, w_eco5465, w_eco5466, w_eco5467, w_eco5468, w_eco5469, w_eco5470, w_eco5471, w_eco5472, w_eco5473, w_eco5474, w_eco5475, w_eco5476, w_eco5477, w_eco5478, w_eco5479, w_eco5480, w_eco5481, w_eco5482, w_eco5483, w_eco5484, w_eco5485, w_eco5486, w_eco5487, w_eco5488, w_eco5489, w_eco5490, w_eco5491, w_eco5492, w_eco5493, w_eco5494, w_eco5495, w_eco5496, w_eco5497, w_eco5498, w_eco5499, w_eco5500, w_eco5501, w_eco5502, w_eco5503, w_eco5504, w_eco5505, w_eco5506, w_eco5507, w_eco5508, w_eco5509, w_eco5510, w_eco5511, w_eco5512, w_eco5513, w_eco5514, w_eco5515, w_eco5516, w_eco5517, w_eco5518, w_eco5519, w_eco5520, w_eco5521, w_eco5522, w_eco5523, w_eco5524, w_eco5525, w_eco5526, w_eco5527, w_eco5528, w_eco5529, w_eco5530, w_eco5531, w_eco5532, w_eco5533, w_eco5534, w_eco5535, w_eco5536, w_eco5537, w_eco5538, w_eco5539, w_eco5540, w_eco5541, w_eco5542, w_eco5543, w_eco5544, w_eco5545, w_eco5546, w_eco5547, w_eco5548, w_eco5549, w_eco5550, w_eco5551, w_eco5552, w_eco5553, w_eco5554, w_eco5555, w_eco5556, w_eco5557, w_eco5558, w_eco5559, w_eco5560, w_eco5561, w_eco5562, w_eco5563, w_eco5564, w_eco5565, w_eco5566, w_eco5567, w_eco5568, w_eco5569, w_eco5570, w_eco5571, w_eco5572, w_eco5573, w_eco5574, w_eco5575, w_eco5576, w_eco5577, w_eco5578, w_eco5579, w_eco5580, w_eco5581, w_eco5582, w_eco5583, w_eco5584, w_eco5585, w_eco5586, w_eco5587, w_eco5588, w_eco5589, w_eco5590, w_eco5591, w_eco5592, w_eco5593, w_eco5594, w_eco5595, w_eco5596, w_eco5597, w_eco5598, w_eco5599, w_eco5600, w_eco5601, w_eco5602, w_eco5603, w_eco5604, w_eco5605, w_eco5606, w_eco5607, w_eco5608, w_eco5609, w_eco5610, w_eco5611, w_eco5612, w_eco5613, w_eco5614, w_eco5615, w_eco5616, w_eco5617, w_eco5618, w_eco5619, w_eco5620, w_eco5621);
	xor _ECO_out9(y[0], sub_wire9, w_eco5622);

endmodule