module top(Sync,Gate,Done,clk,ena,rst,Tsync,Tgdel,Tgate,Tlen,prev_cnt,prev_cnt_len,prev_state);
	input clk, ena, rst;
	input [7:0]Tsync, Tgdel;
	input [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	input [4:0]prev_state;
	output Sync, Gate, Done;
	wire clk, ena, rst;
	wire [7:0]Tsync, Tgdel;
	wire [15:0]Tgate, Tlen, prev_cnt, prev_cnt_len;
	wire [4:0]prev_state;
	wire Sync, Gate, Done, n_130, n_142, n_164, n_167, n_290, n_413, n_414, n_415, n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, sub_wire1, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, sub_wire2, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400, w_eco1401;

	nor g63(n_290, Done, n_458);
	not g70(sub_wire1, n_290);
	nor g91(n_130, n_438, prev_cnt_len[5], prev_cnt_len[11], prev_state[1]);
	nor g103(n_142, n_440, prev_cnt_len[15], prev_cnt_len[9], prev_state[3]);
	nor g105(n_167, n_448, prev_cnt[10], prev_cnt[6], prev_cnt[15]);
	nor g111(n_164, n_453, prev_cnt[14], prev_cnt[3], prev_state[3]);
	not g357(n_413, prev_state[1]);
	not g358(n_414, prev_cnt_len[3]);
	not g359(n_415, prev_state[0]);
	not g360(n_416, prev_cnt_len[0]);
	not g361(n_417, prev_cnt_len[7]);
	not g362(n_418, prev_cnt_len[13]);
	not g363(n_419, prev_cnt_len[4]);
	not g364(n_420, prev_cnt_len[10]);
	not g365(n_421, prev_state[2]);
	not g366(n_422, prev_cnt_len[1]);
	not g367(n_423, prev_cnt_len[6]);
	not g368(n_424, prev_cnt_len[12]);
	not g369(n_425, prev_cnt[1]);
	not g370(n_426, prev_state[4]);
	not g371(n_427, rst);
	not g372(n_428, prev_cnt[4]);
	not g373(n_429, prev_cnt[8]);
	not g374(n_430, prev_cnt[12]);
	not g375(n_431, prev_cnt[5]);
	not g376(n_432, prev_cnt[9]);
	not g377(n_433, prev_cnt[13]);
	not g378(n_434, prev_cnt[7]);
	not g379(n_435, prev_cnt[11]);
	not g380(n_436, ena);
	not g381(n_437, prev_cnt[0]);
	nand g382(n_438, n_415, n_414);
	not g383(n_439, n_130);
	nand g384(n_440, n_418, n_417, n_416);
	not g385(n_441, n_142);
	nand g386(n_442, n_421, n_420, n_419);
	nor g387(n_443, n_442, rst, n_426, prev_cnt_len[2]);
	not g388(n_444, n_443);
	nand g389(n_445, n_424, n_423, n_422);
	nor g390(n_446, n_445, n_436, prev_cnt_len[14], prev_cnt_len[8]);
	not g391(n_447, n_446);
	nor g392(sub_wire0, n_439, n_441, n_444, n_447);
	nand g393(n_448, n_427, n_426, n_425);
	not g394(n_449, n_167);
	nand g395(n_450, n_430, n_429, n_428);
	nor g396(n_451, n_450, n_436, n_421, prev_cnt[2]);
	not g397(n_452, n_451);
	nand g398(n_453, n_433, n_432, n_431);
	nand g399(n_454, n_413, n_435, n_434);
	not g400(n_455, n_454);
	nand g401(n_456, n_164, n_455, n_415, n_437);
	nor g402(sub_wire2, n_449, n_452, n_456);
	nand g403(n_457, ena, n_427, n_426, n_421);
	nor g404(n_458, n_457, prev_state[3], prev_state[1], n_415);
	and _ECO_0(w_eco0, prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1(w_eco1, !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_2(w_eco2, !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_3(w_eco3, prev_state[4], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_4(w_eco4, prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_5(w_eco5, !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_6(w_eco6, !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_7(w_eco7, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_8(w_eco8, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_9(w_eco9, !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_10(w_eco10, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_11(w_eco11, prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_12(w_eco12, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_13(w_eco13, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_14(w_eco14, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_15(w_eco15, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_16(w_eco16, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_17(w_eco17, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_18(w_eco18, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_19(w_eco19, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_20(w_eco20, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_21(w_eco21, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_22(w_eco22, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_23(w_eco23, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_24(w_eco24, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_25(w_eco25, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_26(w_eco26, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_27(w_eco27, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_28(w_eco28, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_29(w_eco29, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	or _ECO_30(w_eco30, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29);
	xor _ECO_out0(Done, sub_wire0, w_eco30);
	and _ECO_31(w_eco31, prev_cnt_len[5], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_32(w_eco32, prev_cnt_len[5], prev_state[1], prev_state[0]);
	and _ECO_33(w_eco33, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], prev_cnt_len[8]);
	and _ECO_34(w_eco34, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], !ena, !prev_cnt_len[14]);
	and _ECO_35(w_eco35, prev_cnt_len[5], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_36(w_eco36, prev_cnt_len[5], !prev_state[3], prev_state[0], !prev_state[2], !rst, ena);
	and _ECO_37(w_eco37, prev_cnt_len[5], !prev_state[3], prev_state[0], !prev_state[2], prev_state[4]);
	and _ECO_38(w_eco38, !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_39(w_eco39, prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_40(w_eco40, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_41(w_eco41, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], !ena, !prev_cnt_len[14]);
	and _ECO_42(w_eco42, prev_cnt_len[5], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_43(w_eco43, !prev_state[0], prev_cnt_len[0], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_44(w_eco44, !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_45(w_eco45, prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14]);
	and _ECO_46(w_eco46, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], prev_cnt_len[1], !prev_cnt_len[14]);
	and _ECO_47(w_eco47, !prev_cnt_len[5], !prev_state[1], prev_state[0], !prev_state[4], !ena, !prev_cnt_len[14]);
	and _ECO_48(w_eco48, !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_49(w_eco49, !prev_cnt_len[5], !prev_state[1], prev_state[0], !prev_state[4], rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_50(w_eco50, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], !prev_cnt_len[6], !prev_cnt_len[12], !prev_cnt_len[14]);
	and _ECO_51(w_eco51, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[10], prev_cnt_len[8]);
	and _ECO_52(w_eco52, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_53(w_eco53, prev_cnt_len[5], prev_state[4], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_54(w_eco54, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_55(w_eco55, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_56(w_eco56, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !rst, ena, prev_cnt_len[14]);
	and _ECO_57(w_eco57, prev_state[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_58(w_eco58, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[1], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_59(w_eco59, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_state[4], rst, prev_cnt_len[8]);
	and _ECO_60(w_eco60, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_61(w_eco61, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], prev_cnt_len[8]);
	and _ECO_62(w_eco62, prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_63(w_eco63, prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2]);
	and _ECO_64(w_eco64, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[6], !prev_cnt_len[12], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_65(w_eco65, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], prev_cnt_len[14]);
	and _ECO_66(w_eco66, prev_cnt_len[5], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_67(w_eco67, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_68(w_eco68, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_69(w_eco69, !prev_state[1], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_70(w_eco70, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_71(w_eco71, !prev_state[1], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_72(w_eco72, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_73(w_eco73, !prev_state[0], prev_state[4], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_74(w_eco74, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_75(w_eco75, prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[14]);
	and _ECO_76(w_eco76, !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_77(w_eco77, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_state[4], rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_78(w_eco78, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, prev_cnt_len[8]);
	and _ECO_79(w_eco79, prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_80(w_eco80, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], prev_cnt_len[8]);
	and _ECO_81(w_eco81, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_82(w_eco82, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_cnt_len[14]);
	and _ECO_83(w_eco83, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[1], !prev_cnt_len[6], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_84(w_eco84, !prev_cnt_len[5], !prev_state[1], prev_state[0], !prev_cnt_len[6], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_85(w_eco85, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_state[4], !ena, prev_cnt_len[8]);
	and _ECO_86(w_eco86, prev_cnt_len[5], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_87(w_eco87, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_88(w_eco88, prev_cnt_len[5], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_89(w_eco89, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_90(w_eco90, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_91(w_eco91, !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_92(w_eco92, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_93(w_eco93, !prev_state[1], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_94(w_eco94, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_95(w_eco95, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_96(w_eco96, !prev_state[0], prev_cnt_len[0], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_97(w_eco97, !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_98(w_eco98, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_99(w_eco99, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_100(w_eco100, prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14]);
	and _ECO_101(w_eco101, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], rst, prev_cnt_len[8]);
	and _ECO_102(w_eco102, !prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, ena, !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_103(w_eco103, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_state[2], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_104(w_eco104, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_105(w_eco105, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_106(w_eco106, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2]);
	and _ECO_107(w_eco107, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !ena, prev_cnt_len[8]);
	and _ECO_108(w_eco108, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_109(w_eco109, prev_cnt_len[5], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_110(w_eco110, prev_cnt_len[5], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_111(w_eco111, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_112(w_eco112, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_113(w_eco113, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_114(w_eco114, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_115(w_eco115, !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], rst, ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_116(w_eco116, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_117(w_eco117, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_118(w_eco118, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_119(w_eco119, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_120(w_eco120, !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_121(w_eco121, !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], rst, ena, !prev_cnt_len[8]);
	and _ECO_122(w_eco122, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_123(w_eco123, !prev_state[0], rst, prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_124(w_eco124, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_125(w_eco125, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_126(w_eco126, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_127(w_eco127, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_128(w_eco128, !prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, ena, prev_cnt_len[14]);
	and _ECO_129(w_eco129, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_130(w_eco130, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_131(w_eco131, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_132(w_eco132, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_133(w_eco133, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_134(w_eco134, !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[2]);
	and _ECO_135(w_eco135, prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[2]);
	and _ECO_136(w_eco136, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[6], !prev_state[4], rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_137(w_eco137, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !ena, prev_cnt_len[8]);
	and _ECO_138(w_eco138, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[10], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_139(w_eco139, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_140(w_eco140, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_141(w_eco141, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_142(w_eco142, prev_cnt_len[5], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_143(w_eco143, prev_cnt_len[5], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_144(w_eco144, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14], prev_cnt_len[8]);
	and _ECO_145(w_eco145, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_146(w_eco146, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_147(w_eco147, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_148(w_eco148, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_149(w_eco149, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_150(w_eco150, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_151(w_eco151, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_152(w_eco152, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_153(w_eco153, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], prev_cnt_len[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_154(w_eco154, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_155(w_eco155, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_156(w_eco156, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_157(w_eco157, !prev_state[0], prev_cnt_len[0], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_158(w_eco158, !prev_state[0], prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_159(w_eco159, !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_160(w_eco160, !prev_state[0], prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_161(w_eco161, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_162(w_eco162, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_163(w_eco163, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_164(w_eco164, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_165(w_eco165, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[10], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_166(w_eco166, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_167(w_eco167, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_168(w_eco168, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[14]);
	and _ECO_169(w_eco169, prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], ena, !prev_cnt_len[2]);
	and _ECO_170(w_eco170, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[0], !prev_cnt_len[6], !prev_state[4], rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_171(w_eco171, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[10], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_172(w_eco172, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_173(w_eco173, prev_state[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_174(w_eco174, prev_cnt_len[5], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_175(w_eco175, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_176(w_eco176, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_177(w_eco177, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_178(w_eco178, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_179(w_eco179, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt_len[8]);
	and _ECO_180(w_eco180, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_181(w_eco181, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_182(w_eco182, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_183(w_eco183, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_184(w_eco184, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_state[2], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_185(w_eco185, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_186(w_eco186, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_187(w_eco187, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_188(w_eco188, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_189(w_eco189, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_190(w_eco190, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_191(w_eco191, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_192(w_eco192, !prev_state[0], prev_cnt_len[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_193(w_eco193, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_194(w_eco194, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_195(w_eco195, !prev_state[0], prev_cnt_len[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_196(w_eco196, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_197(w_eco197, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_198(w_eco198, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_199(w_eco199, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_200(w_eco200, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_state[2], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_201(w_eco201, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_202(w_eco202, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_203(w_eco203, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_204(w_eco204, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], prev_cnt_len[10], prev_cnt_len[1], !prev_cnt_len[14]);
	and _ECO_205(w_eco205, !prev_cnt_len[5], !prev_state[1], prev_state[0], prev_cnt_len[10], prev_cnt_len[1], !prev_state[4], rst, !prev_cnt_len[14]);
	and _ECO_206(w_eco206, !prev_cnt_len[5], !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[6], !prev_state[4], !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_207(w_eco207, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[10], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_208(w_eco208, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_209(w_eco209, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_210(w_eco210, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_211(w_eco211, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_212(w_eco212, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt_len[8]);
	and _ECO_213(w_eco213, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_214(w_eco214, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_215(w_eco215, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_216(w_eco216, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_217(w_eco217, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_218(w_eco218, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_219(w_eco219, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_220(w_eco220, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], prev_cnt_len[9], !prev_state[3], !prev_state[0], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_221(w_eco221, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_222(w_eco222, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_223(w_eco223, !prev_state[1], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_224(w_eco224, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_225(w_eco225, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_226(w_eco226, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_227(w_eco227, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_228(w_eco228, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_229(w_eco229, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_230(w_eco230, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], rst, ena, !prev_cnt_len[8]);
	and _ECO_231(w_eco231, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_232(w_eco232, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_233(w_eco233, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_234(w_eco234, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_235(w_eco235, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt_len[8]);
	and _ECO_236(w_eco236, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_237(w_eco237, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_238(w_eco238, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_239(w_eco239, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_cnt_len[12], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_240(w_eco240, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_241(w_eco241, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_state[2], !prev_state[4], !prev_cnt_len[2]);
	and _ECO_242(w_eco242, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_243(w_eco243, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_244(w_eco244, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_245(w_eco245, prev_state[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_246(w_eco246, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_247(w_eco247, !prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, ena, !prev_cnt_len[2]);
	and _ECO_248(w_eco248, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], prev_cnt_len[0], !prev_cnt_len[6], !prev_state[4], rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_249(w_eco249, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_250(w_eco250, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_251(w_eco251, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_252(w_eco252, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_253(w_eco253, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_254(w_eco254, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_255(w_eco255, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_256(w_eco256, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_257(w_eco257, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], prev_cnt_len[4], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_258(w_eco258, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_259(w_eco259, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_260(w_eco260, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_261(w_eco261, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[15], prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_262(w_eco262, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_263(w_eco263, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_264(w_eco264, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_265(w_eco265, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_266(w_eco266, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_267(w_eco267, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_268(w_eco268, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_269(w_eco269, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_270(w_eco270, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_271(w_eco271, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_272(w_eco272, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_273(w_eco273, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_274(w_eco274, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_275(w_eco275, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_276(w_eco276, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_277(w_eco277, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_278(w_eco278, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[0], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_279(w_eco279, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_280(w_eco280, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], prev_cnt_len[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_281(w_eco281, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_282(w_eco282, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_283(w_eco283, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_284(w_eco284, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_285(w_eco285, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_286(w_eco286, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_287(w_eco287, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_288(w_eco288, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_289(w_eco289, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_290(w_eco290, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_291(w_eco291, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_292(w_eco292, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt_len[8]);
	and _ECO_293(w_eco293, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[15], prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_294(w_eco294, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_295(w_eco295, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_296(w_eco296, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2]);
	and _ECO_297(w_eco297, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_298(w_eco298, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_299(w_eco299, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_300(w_eco300, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[13], prev_state[2], !prev_state[4], !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_301(w_eco301, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_302(w_eco302, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_303(w_eco303, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_304(w_eco304, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_305(w_eco305, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_306(w_eco306, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_307(w_eco307, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_308(w_eco308, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_309(w_eco309, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_310(w_eco310, !prev_state[1], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_311(w_eco311, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_312(w_eco312, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_313(w_eco313, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_314(w_eco314, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_315(w_eco315, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_316(w_eco316, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_317(w_eco317, !prev_state[1], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_318(w_eco318, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_319(w_eco319, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_320(w_eco320, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_321(w_eco321, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_322(w_eco322, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_323(w_eco323, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_324(w_eco324, !prev_state[1], !prev_state[0], !prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_325(w_eco325, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_326(w_eco326, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_327(w_eco327, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_328(w_eco328, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_329(w_eco329, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_330(w_eco330, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_331(w_eco331, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_332(w_eco332, prev_cnt_len[5], prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_333(w_eco333, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_334(w_eco334, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_335(w_eco335, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_336(w_eco336, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[6], !prev_state[4], rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_337(w_eco337, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_338(w_eco338, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !ena, !prev_cnt_len[2]);
	and _ECO_339(w_eco339, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_340(w_eco340, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_341(w_eco341, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_342(w_eco342, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !prev_state[4], !rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_343(w_eco343, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_344(w_eco344, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_345(w_eco345, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_346(w_eco346, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], prev_cnt_len[10], !rst, !prev_cnt_len[2]);
	and _ECO_347(w_eco347, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_348(w_eco348, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_349(w_eco349, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_350(w_eco350, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], !prev_cnt_len[10], !prev_state[2], prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_351(w_eco351, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_352(w_eco352, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_353(w_eco353, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_354(w_eco354, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_355(w_eco355, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_356(w_eco356, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_357(w_eco357, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_358(w_eco358, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_359(w_eco359, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_360(w_eco360, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_361(w_eco361, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_362(w_eco362, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt_len[14]);
	and _ECO_363(w_eco363, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_364(w_eco364, prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_365(w_eco365, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_366(w_eco366, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_367(w_eco367, !prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_368(w_eco368, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_369(w_eco369, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_370(w_eco370, !prev_state[1], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_371(w_eco371, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_372(w_eco372, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2]);
	and _ECO_373(w_eco373, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt_len[12], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_374(w_eco374, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_375(w_eco375, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[9], prev_state[0], !prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_376(w_eco376, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt_len[8]);
	and _ECO_377(w_eco377, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_378(w_eco378, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_379(w_eco379, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_380(w_eco380, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], rst, !prev_cnt_len[2], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_381(w_eco381, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_382(w_eco382, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_383(w_eco383, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_384(w_eco384, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], rst, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_385(w_eco385, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_386(w_eco386, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_387(w_eco387, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_388(w_eco388, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_389(w_eco389, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_390(w_eco390, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_391(w_eco391, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_392(w_eco392, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[10], !prev_cnt_len[1], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_393(w_eco393, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_394(w_eco394, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_395(w_eco395, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_396(w_eco396, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_397(w_eco397, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[13], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_398(w_eco398, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[4], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_399(w_eco399, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], prev_cnt_len[10], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_400(w_eco400, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_401(w_eco401, !prev_state[1], !prev_state[0], !prev_cnt_len[13], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_402(w_eco402, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_403(w_eco403, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[12], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_404(w_eco404, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[15], prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_405(w_eco405, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[12], ena, !prev_cnt_len[8]);
	and _ECO_406(w_eco406, prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_407(w_eco407, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, ena, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_408(w_eco408, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_409(w_eco409, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt_len[8]);
	and _ECO_410(w_eco410, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_411(w_eco411, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt_len[2]);
	and _ECO_412(w_eco412, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, ena, prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_413(w_eco413, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], prev_cnt_len[1], !rst, !prev_cnt_len[14]);
	and _ECO_414(w_eco414, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_cnt_len[1], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_415(w_eco415, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_416(w_eco416, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_417(w_eco417, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[8]);
	and _ECO_418(w_eco418, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[1], prev_cnt_len[6], ena, !prev_cnt_len[8]);
	and _ECO_419(w_eco419, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[0], !prev_cnt_len[7], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_state[4], ena, !prev_cnt_len[8]);
	and _ECO_420(w_eco420, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_421(w_eco421, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt_len[8]);
	and _ECO_422(w_eco422, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[1], !prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_423(w_eco423, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_424(w_eco424, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[1], !prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], rst, ena, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_425(w_eco425, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_426(w_eco426, !prev_cnt_len[5], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_427(w_eco427, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt_len[8]);
	or _ECO_428(w_eco428, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427);
	xor _ECO_out1(Sync, sub_wire1, w_eco428);
	and _ECO_429(w_eco429, prev_state[1], prev_state[0], prev_cnt[0]);
	and _ECO_430(w_eco430, !prev_cnt_len[5], prev_state[0], !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_431(w_eco431, prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], !prev_cnt[0], prev_cnt[2]);
	and _ECO_432(w_eco432, prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], !ena, !prev_cnt[0]);
	and _ECO_433(w_eco433, prev_state[3], prev_state[0], !prev_state[2], !rst, prev_cnt[0]);
	and _ECO_434(w_eco434, prev_cnt_len[5], !prev_state[1], prev_state[0], rst, !prev_cnt[0], prev_cnt[2]);
	and _ECO_435(w_eco435, prev_state[0], !prev_state[2], !prev_state[4], !rst, ena, prev_cnt[0]);
	and _ECO_436(w_eco436, !prev_cnt_len[5], prev_state[0], prev_state[2], prev_cnt[0]);
	and _ECO_437(w_eco437, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_state[0], !ena, !prev_cnt[0], prev_cnt[2]);
	and _ECO_438(w_eco438, !prev_cnt_len[5], prev_state[0], prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_439(w_eco439, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_440(w_eco440, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_state[0], prev_state[4], !prev_cnt[0], prev_cnt[2]);
	and _ECO_441(w_eco441, prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[0]);
	and _ECO_442(w_eco442, prev_state[1], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[2]);
	and _ECO_443(w_eco443, prev_cnt_len[5], !prev_state[1], prev_cnt[15], prev_state[0], rst, !prev_cnt[0]);
	and _ECO_444(w_eco444, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_445(w_eco445, !prev_cnt_len[5], prev_state[0], prev_cnt_len[10], prev_cnt[0]);
	and _ECO_446(w_eco446, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_447(w_eco447, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_448(w_eco448, prev_cnt_len[5], !prev_state[1], prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[0]);
	and _ECO_449(w_eco449, prev_cnt_len[5], !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], rst, !prev_cnt[0]);
	and _ECO_450(w_eco450, prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_451(w_eco451, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !ena, !prev_cnt[0]);
	and _ECO_452(w_eco452, prev_cnt_len[5], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_453(w_eco453, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_454(w_eco454, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_455(w_eco455, !prev_cnt_len[5], prev_state[0], prev_cnt_len[1], !prev_cnt_len[12], prev_cnt[0]);
	and _ECO_456(w_eco456, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_457(w_eco457, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_458(w_eco458, prev_state[1], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_459(w_eco459, prev_cnt_len[5], !prev_state[1], prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[0]);
	and _ECO_460(w_eco460, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], rst, !prev_cnt[2]);
	and _ECO_461(w_eco461, prev_cnt_len[5], !prev_state[1], !prev_cnt[6], prev_state[0], prev_cnt[1], rst, !prev_cnt[0]);
	and _ECO_462(w_eco462, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], prev_state[4], !prev_cnt[0]);
	and _ECO_463(w_eco463, prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_state[4], !rst, ena, !prev_cnt[2]);
	and _ECO_464(w_eco464, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_state[4], !rst, !ena, !prev_cnt[0]);
	and _ECO_465(w_eco465, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_466(w_eco466, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[3], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_467(w_eco467, !prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_468(w_eco468, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_469(w_eco469, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_470(w_eco470, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_471(w_eco471, !prev_cnt_len[5], prev_state[0], prev_cnt_len[4], !prev_cnt_len[12], prev_cnt[0]);
	and _ECO_472(w_eco472, !prev_cnt_len[5], !prev_state[3], prev_state[0], !prev_cnt_len[12], prev_state[4], prev_cnt[0]);
	and _ECO_473(w_eco473, !prev_cnt_len[5], prev_state[0], !prev_cnt_len[6], prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_474(w_eco474, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_475(w_eco475, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_476(w_eco476, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_477(w_eco477, prev_state[1], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_478(w_eco478, prev_cnt_len[5], !prev_state[1], !prev_cnt[6], prev_state[0], prev_state[2], !prev_state[4], !rst, !prev_cnt[0]);
	and _ECO_479(w_eco479, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], prev_state[4], !prev_cnt[2]);
	and _ECO_480(w_eco480, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], prev_state[4], !prev_cnt[0]);
	and _ECO_481(w_eco481, prev_cnt_len[5], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_482(w_eco482, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_483(w_eco483, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_484(w_eco484, !prev_state[1], !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !ena, !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_485(w_eco485, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_486(w_eco486, !prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_487(w_eco487, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_488(w_eco488, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_489(w_eco489, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_490(w_eco490, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_491(w_eco491, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_492(w_eco492, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_493(w_eco493, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_494(w_eco494, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_495(w_eco495, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_496(w_eco496, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_497(w_eco497, prev_state[3], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_498(w_eco498, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], prev_cnt[1], prev_state[4], !prev_cnt[0]);
	and _ECO_499(w_eco499, prev_cnt_len[5], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_500(w_eco500, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_501(w_eco501, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_502(w_eco502, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_503(w_eco503, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_504(w_eco504, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_505(w_eco505, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_506(w_eco506, !prev_state[1], !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_507(w_eco507, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], prev_cnt_len[10], !prev_state[2], !prev_cnt[2]);
	and _ECO_508(w_eco508, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_509(w_eco509, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_510(w_eco510, !prev_state[1], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_511(w_eco511, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_512(w_eco512, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_513(w_eco513, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_514(w_eco514, !prev_state[3], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_515(w_eco515, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_516(w_eco516, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_517(w_eco517, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_518(w_eco518, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_519(w_eco519, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_520(w_eco520, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_521(w_eco521, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, prev_cnt[0], !prev_cnt_len[14]);
	and _ECO_522(w_eco522, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_523(w_eco523, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_524(w_eco524, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_525(w_eco525, prev_cnt_len[5], !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], prev_state[2], !prev_cnt[0]);
	and _ECO_526(w_eco526, !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_527(w_eco527, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[3], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_528(w_eco528, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_529(w_eco529, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_530(w_eco530, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_531(w_eco531, prev_cnt_len[5], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_532(w_eco532, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_533(w_eco533, !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_534(w_eco534, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_535(w_eco535, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_536(w_eco536, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !prev_cnt[2]);
	and _ECO_537(w_eco537, !prev_state[1], !prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !ena, !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_538(w_eco538, !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !ena, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_539(w_eco539, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_540(w_eco540, !prev_state[1], !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_541(w_eco541, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_542(w_eco542, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_543(w_eco543, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_544(w_eco544, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_545(w_eco545, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_546(w_eco546, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_547(w_eco547, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_548(w_eco548, !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_549(w_eco549, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_550(w_eco550, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_551(w_eco551, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_552(w_eco552, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[0]);
	and _ECO_553(w_eco553, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_554(w_eco554, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_555(w_eco555, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_556(w_eco556, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_557(w_eco557, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_558(w_eco558, prev_state[1], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_559(w_eco559, prev_cnt_len[5], !prev_state[1], !prev_cnt[6], prev_state[0], prev_state[2], prev_cnt[1], !prev_cnt[0]);
	and _ECO_560(w_eco560, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_561(w_eco561, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_562(w_eco562, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_563(w_eco563, !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_564(w_eco564, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_565(w_eco565, prev_cnt_len[5], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_566(w_eco566, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_567(w_eco567, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_568(w_eco568, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_569(w_eco569, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_570(w_eco570, !prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_571(w_eco571, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_572(w_eco572, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], rst, !prev_cnt[2]);
	and _ECO_573(w_eco573, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_574(w_eco574, !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_575(w_eco575, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !prev_cnt[2]);
	and _ECO_576(w_eco576, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !ena, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_577(w_eco577, !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_578(w_eco578, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_579(w_eco579, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], prev_state[4], !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_580(w_eco580, !prev_state[1], !prev_state[3], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_581(w_eco581, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_582(w_eco582, !prev_cnt_len[5], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt_len[6], !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_583(w_eco583, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_584(w_eco584, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_585(w_eco585, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_586(w_eco586, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_587(w_eco587, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_588(w_eco588, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[7], !ena, !prev_cnt_len[14]);
	and _ECO_589(w_eco589, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_590(w_eco590, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_591(w_eco591, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_592(w_eco592, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[11], !ena, !prev_cnt_len[14]);
	and _ECO_593(w_eco593, !prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_594(w_eco594, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_595(w_eco595, !prev_state[3], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_596(w_eco596, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_597(w_eco597, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_598(w_eco598, !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_599(w_eco599, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[0]);
	and _ECO_600(w_eco600, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_601(w_eco601, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_602(w_eco602, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_603(w_eco603, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_604(w_eco604, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_605(w_eco605, !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_606(w_eco606, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[3], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_607(w_eco607, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_608(w_eco608, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_609(w_eco609, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_610(w_eco610, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_611(w_eco611, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_612(w_eco612, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_613(w_eco613, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_614(w_eco614, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_615(w_eco615, prev_cnt_len[5], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_616(w_eco616, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_617(w_eco617, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_618(w_eco618, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_619(w_eco619, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_620(w_eco620, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_621(w_eco621, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_622(w_eco622, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !prev_cnt[1], rst, !prev_cnt[2]);
	and _ECO_623(w_eco623, !prev_state[1], prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_624(w_eco624, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !ena, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_625(w_eco625, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt[1], prev_state[4], prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_626(w_eco626, !prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_627(w_eco627, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_628(w_eco628, !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_629(w_eco629, !prev_state[1], prev_state[3], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_630(w_eco630, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_631(w_eco631, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[7]);
	and _ECO_632(w_eco632, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_633(w_eco633, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_634(w_eco634, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_635(w_eco635, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_636(w_eco636, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_637(w_eco637, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst);
	and _ECO_638(w_eco638, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[11], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_639(w_eco639, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_640(w_eco640, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_641(w_eco641, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_642(w_eco642, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_643(w_eco643, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_644(w_eco644, !prev_state[3], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_645(w_eco645, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_646(w_eco646, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_647(w_eco647, !prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_648(w_eco648, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_649(w_eco649, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_650(w_eco650, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_651(w_eco651, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_652(w_eco652, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_653(w_eco653, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_654(w_eco654, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_655(w_eco655, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_656(w_eco656, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt[1], prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_657(w_eco657, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_658(w_eco658, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_659(w_eco659, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_660(w_eco660, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_661(w_eco661, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_662(w_eco662, prev_cnt_len[5], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_663(w_eco663, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_664(w_eco664, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_665(w_eco665, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_666(w_eco666, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_667(w_eco667, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_668(w_eco668, prev_cnt_len[5], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_669(w_eco669, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[1], rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_670(w_eco670, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_671(w_eco671, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !prev_cnt[2]);
	and _ECO_672(w_eco672, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_673(w_eco673, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], rst, !prev_cnt[2]);
	and _ECO_674(w_eco674, !prev_state[1], prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_675(w_eco675, !prev_cnt_len[5], !prev_state[3], prev_cnt[6], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt_len[12], prev_state[4], !prev_cnt[2]);
	and _ECO_676(w_eco676, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_677(w_eco677, !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !ena, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_678(w_eco678, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_679(w_eco679, !prev_state[1], prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_680(w_eco680, !prev_state[1], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_681(w_eco681, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_682(w_eco682, !prev_state[1], !prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_683(w_eco683, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_684(w_eco684, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[7]);
	and _ECO_685(w_eco685, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_686(w_eco686, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_687(w_eco687, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_688(w_eco688, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_689(w_eco689, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_690(w_eco690, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[11]);
	and _ECO_691(w_eco691, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst);
	and _ECO_692(w_eco692, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_693(w_eco693, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_694(w_eco694, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_695(w_eco695, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_696(w_eco696, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_697(w_eco697, !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_698(w_eco698, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_699(w_eco699, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_700(w_eco700, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_701(w_eco701, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_702(w_eco702, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_703(w_eco703, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_704(w_eco704, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_705(w_eco705, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_706(w_eco706, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_707(w_eco707, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_708(w_eco708, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_709(w_eco709, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_710(w_eco710, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[0]);
	and _ECO_711(w_eco711, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[0], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_712(w_eco712, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_713(w_eco713, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_714(w_eco714, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_715(w_eco715, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_716(w_eco716, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_717(w_eco717, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_718(w_eco718, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_719(w_eco719, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_720(w_eco720, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_721(w_eco721, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_722(w_eco722, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_723(w_eco723, prev_cnt_len[5], prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_724(w_eco724, prev_cnt_len[5], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_725(w_eco725, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], prev_state[2], !prev_cnt[1], prev_state[4], !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_726(w_eco726, !prev_cnt_len[5], !prev_state[3], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !prev_cnt[2]);
	and _ECO_727(w_eco727, !prev_state[1], prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt[1], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_728(w_eco728, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_729(w_eco729, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt[1], !prev_state[4], rst, !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_730(w_eco730, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_731(w_eco731, !prev_state[1], prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_732(w_eco732, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_733(w_eco733, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_734(w_eco734, !prev_state[1], prev_state[3], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_735(w_eco735, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_736(w_eco736, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_737(w_eco737, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_738(w_eco738, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_739(w_eco739, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_740(w_eco740, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_741(w_eco741, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_742(w_eco742, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[11]);
	and _ECO_743(w_eco743, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_744(w_eco744, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_745(w_eco745, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst);
	and _ECO_746(w_eco746, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_747(w_eco747, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_748(w_eco748, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_749(w_eco749, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_750(w_eco750, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_751(w_eco751, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_752(w_eco752, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_753(w_eco753, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_754(w_eco754, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_755(w_eco755, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !prev_cnt[11], !ena, !prev_cnt_len[14]);
	and _ECO_756(w_eco756, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_757(w_eco757, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_758(w_eco758, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_759(w_eco759, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_760(w_eco760, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_761(w_eco761, !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_762(w_eco762, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_763(w_eco763, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_764(w_eco764, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_765(w_eco765, !prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_766(w_eco766, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_767(w_eco767, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_768(w_eco768, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_769(w_eco769, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_770(w_eco770, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_771(w_eco771, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_772(w_eco772, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[0], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_773(w_eco773, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_774(w_eco774, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_775(w_eco775, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[14], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_776(w_eco776, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_777(w_eco777, prev_cnt_len[5], prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_778(w_eco778, prev_cnt_len[5], !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_779(w_eco779, !prev_state[1], prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_780(w_eco780, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_781(w_eco781, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], prev_state[4], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_782(w_eco782, !prev_state[1], prev_state[3], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_783(w_eco783, !prev_state[1], prev_cnt[15], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_784(w_eco784, !prev_cnt_len[5], !prev_cnt[10], !prev_cnt[15], prev_state[0], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_785(w_eco785, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_786(w_eco786, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[7]);
	and _ECO_787(w_eco787, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[7], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_788(w_eco788, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_789(w_eco789, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_790(w_eco790, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst);
	and _ECO_791(w_eco791, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_792(w_eco792, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_793(w_eco793, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_794(w_eco794, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_795(w_eco795, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_796(w_eco796, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_797(w_eco797, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst);
	and _ECO_798(w_eco798, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_799(w_eco799, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_800(w_eco800, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_801(w_eco801, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_802(w_eco802, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_803(w_eco803, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_804(w_eco804, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !prev_cnt[11], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_805(w_eco805, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_806(w_eco806, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_807(w_eco807, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_808(w_eco808, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[11], !ena, !prev_cnt_len[14]);
	and _ECO_809(w_eco809, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_810(w_eco810, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_811(w_eco811, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_812(w_eco812, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_813(w_eco813, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_814(w_eco814, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_815(w_eco815, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_816(w_eco816, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_817(w_eco817, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_818(w_eco818, !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_819(w_eco819, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_820(w_eco820, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_821(w_eco821, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_822(w_eco822, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_823(w_eco823, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_824(w_eco824, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_825(w_eco825, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_826(w_eco826, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_827(w_eco827, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_828(w_eco828, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_829(w_eco829, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_830(w_eco830, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_831(w_eco831, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[0]);
	and _ECO_832(w_eco832, prev_cnt_len[5], !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_833(w_eco833, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt[1], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_834(w_eco834, !prev_state[1], prev_state[3], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt[1], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_835(w_eco835, !prev_state[1], prev_cnt[10], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_836(w_eco836, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_837(w_eco837, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_838(w_eco838, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[7], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_839(w_eco839, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst);
	and _ECO_840(w_eco840, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[11]);
	and _ECO_841(w_eco841, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst);
	and _ECO_842(w_eco842, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_843(w_eco843, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_844(w_eco844, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_845(w_eco845, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_846(w_eco846, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_847(w_eco847, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_848(w_eco848, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_849(w_eco849, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_850(w_eco850, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_851(w_eco851, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_852(w_eco852, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_853(w_eco853, !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_854(w_eco854, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_855(w_eco855, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_856(w_eco856, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_857(w_eco857, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_858(w_eco858, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_859(w_eco859, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_860(w_eco860, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[11], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_861(w_eco861, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_862(w_eco862, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_863(w_eco863, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_864(w_eco864, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_865(w_eco865, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_866(w_eco866, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_867(w_eco867, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_868(w_eco868, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_869(w_eco869, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_870(w_eco870, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_871(w_eco871, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_872(w_eco872, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_873(w_eco873, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_874(w_eco874, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_875(w_eco875, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_876(w_eco876, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_877(w_eco877, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_878(w_eco878, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_879(w_eco879, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_880(w_eco880, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_881(w_eco881, !prev_cnt_len[15], !prev_state[3], prev_cnt[15], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_882(w_eco882, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_883(w_eco883, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_884(w_eco884, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_885(w_eco885, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_886(w_eco886, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_887(w_eco887, !prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_888(w_eco888, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_889(w_eco889, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_890(w_eco890, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_891(w_eco891, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[11], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_892(w_eco892, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_893(w_eco893, !prev_state[1], !prev_cnt[6], prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], prev_cnt[1], !prev_state[4], rst, ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_894(w_eco894, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[7]);
	and _ECO_895(w_eco895, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_896(w_eco896, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[11]);
	and _ECO_897(w_eco897, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst);
	and _ECO_898(w_eco898, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[11]);
	and _ECO_899(w_eco899, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_900(w_eco900, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_901(w_eco901, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_902(w_eco902, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_903(w_eco903, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_904(w_eco904, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_905(w_eco905, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst);
	and _ECO_906(w_eco906, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_907(w_eco907, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_908(w_eco908, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_909(w_eco909, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_910(w_eco910, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_911(w_eco911, !prev_state[3], prev_cnt[3], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_912(w_eco912, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_913(w_eco913, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_914(w_eco914, !prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_915(w_eco915, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_916(w_eco916, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_917(w_eco917, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_918(w_eco918, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_919(w_eco919, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_920(w_eco920, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_921(w_eco921, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_922(w_eco922, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_923(w_eco923, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_924(w_eco924, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_925(w_eco925, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_926(w_eco926, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_927(w_eco927, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_928(w_eco928, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_929(w_eco929, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_930(w_eco930, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_931(w_eco931, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_932(w_eco932, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[5], !ena, !prev_cnt_len[14]);
	and _ECO_933(w_eco933, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_934(w_eco934, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt[2]);
	and _ECO_935(w_eco935, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_936(w_eco936, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_937(w_eco937, !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], rst, !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_938(w_eco938, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_939(w_eco939, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_940(w_eco940, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_941(w_eco941, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_942(w_eco942, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_943(w_eco943, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_944(w_eco944, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_945(w_eco945, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_946(w_eco946, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_947(w_eco947, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_948(w_eco948, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_949(w_eco949, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_950(w_eco950, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_951(w_eco951, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_952(w_eco952, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_953(w_eco953, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_954(w_eco954, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_955(w_eco955, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_956(w_eco956, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_957(w_eco957, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_958(w_eco958, !prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_959(w_eco959, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_960(w_eco960, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_961(w_eco961, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_962(w_eco962, !prev_cnt_len[5], prev_cnt_len[15], prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_963(w_eco963, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_964(w_eco964, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_965(w_eco965, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_966(w_eco966, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_967(w_eco967, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[11]);
	and _ECO_968(w_eco968, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_969(w_eco969, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_970(w_eco970, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_971(w_eco971, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_972(w_eco972, !prev_cnt_len[5], !prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[11]);
	and _ECO_973(w_eco973, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_974(w_eco974, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_975(w_eco975, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_976(w_eco976, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_977(w_eco977, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst);
	and _ECO_978(w_eco978, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst);
	and _ECO_979(w_eco979, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_980(w_eco980, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_981(w_eco981, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_982(w_eco982, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_983(w_eco983, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_984(w_eco984, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_985(w_eco985, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_986(w_eco986, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_987(w_eco987, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_988(w_eco988, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_989(w_eco989, !prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_990(w_eco990, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_991(w_eco991, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_992(w_eco992, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_993(w_eco993, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_994(w_eco994, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_995(w_eco995, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_996(w_eco996, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_997(w_eco997, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_998(w_eco998, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_999(w_eco999, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1000(w_eco1000, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1001(w_eco1001, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1002(w_eco1002, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt[5], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1003(w_eco1003, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1004(w_eco1004, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1005(w_eco1005, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1006(w_eco1006, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1007(w_eco1007, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1008(w_eco1008, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1009(w_eco1009, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1010(w_eco1010, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1011(w_eco1011, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !ena, !prev_cnt_len[14]);
	and _ECO_1012(w_eco1012, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_1013(w_eco1013, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_1014(w_eco1014, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1015(w_eco1015, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1016(w_eco1016, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1017(w_eco1017, !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1018(w_eco1018, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1019(w_eco1019, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1020(w_eco1020, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1021(w_eco1021, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1022(w_eco1022, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1023(w_eco1023, !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1024(w_eco1024, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1025(w_eco1025, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_1026(w_eco1026, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !ena, !prev_cnt[0]);
	and _ECO_1027(w_eco1027, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_1028(w_eco1028, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1029(w_eco1029, !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1030(w_eco1030, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1031(w_eco1031, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1032(w_eco1032, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1033(w_eco1033, prev_state[1], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1034(w_eco1034, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1035(w_eco1035, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1036(w_eco1036, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1037(w_eco1037, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1038(w_eco1038, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1039(w_eco1039, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_1040(w_eco1040, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1041(w_eco1041, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_1042(w_eco1042, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1043(w_eco1043, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_1044(w_eco1044, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, prev_cnt[5]);
	and _ECO_1045(w_eco1045, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_1046(w_eco1046, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1047(w_eco1047, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1048(w_eco1048, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_1049(w_eco1049, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_1050(w_eco1050, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst);
	and _ECO_1051(w_eco1051, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1052(w_eco1052, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1053(w_eco1053, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_1054(w_eco1054, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1055(w_eco1055, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1056(w_eco1056, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1057(w_eco1057, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1058(w_eco1058, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1059(w_eco1059, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1060(w_eco1060, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1061(w_eco1061, !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1062(w_eco1062, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1063(w_eco1063, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_1064(w_eco1064, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1065(w_eco1065, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1066(w_eco1066, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1067(w_eco1067, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1068(w_eco1068, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1069(w_eco1069, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1070(w_eco1070, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1071(w_eco1071, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1072(w_eco1072, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1073(w_eco1073, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1074(w_eco1074, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1075(w_eco1075, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1076(w_eco1076, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1077(w_eco1077, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1078(w_eco1078, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1079(w_eco1079, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1080(w_eco1080, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1081(w_eco1081, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1082(w_eco1082, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1083(w_eco1083, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1084(w_eco1084, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1085(w_eco1085, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1086(w_eco1086, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1087(w_eco1087, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1088(w_eco1088, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1089(w_eco1089, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1090(w_eco1090, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1091(w_eco1091, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt[2]);
	and _ECO_1092(w_eco1092, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], !ena, !prev_cnt_len[14]);
	and _ECO_1093(w_eco1093, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1094(w_eco1094, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1095(w_eco1095, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1096(w_eco1096, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1097(w_eco1097, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1098(w_eco1098, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1099(w_eco1099, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_1100(w_eco1100, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_1101(w_eco1101, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1102(w_eco1102, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1103(w_eco1103, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1104(w_eco1104, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1105(w_eco1105, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1106(w_eco1106, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1107(w_eco1107, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1108(w_eco1108, prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1109(w_eco1109, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1110(w_eco1110, !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1111(w_eco1111, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1112(w_eco1112, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1113(w_eco1113, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1114(w_eco1114, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1115(w_eco1115, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1116(w_eco1116, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1117(w_eco1117, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1118(w_eco1118, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[11], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1119(w_eco1119, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1120(w_eco1120, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1121(w_eco1121, !prev_cnt_len[5], prev_cnt_len[15], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1122(w_eco1122, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1123(w_eco1123, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1124(w_eco1124, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[11]);
	and _ECO_1125(w_eco1125, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, prev_cnt[5]);
	and _ECO_1126(w_eco1126, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1127(w_eco1127, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_1128(w_eco1128, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1129(w_eco1129, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst);
	and _ECO_1130(w_eco1130, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_1131(w_eco1131, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1132(w_eco1132, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1133(w_eco1133, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_1134(w_eco1134, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_1135(w_eco1135, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1136(w_eco1136, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1137(w_eco1137, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1138(w_eco1138, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1139(w_eco1139, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1140(w_eco1140, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1141(w_eco1141, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1142(w_eco1142, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1143(w_eco1143, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1144(w_eco1144, !prev_cnt_len[15], !prev_state[3], prev_cnt[3], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1145(w_eco1145, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1146(w_eco1146, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_1147(w_eco1147, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1148(w_eco1148, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1149(w_eco1149, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1150(w_eco1150, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1151(w_eco1151, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1152(w_eco1152, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1153(w_eco1153, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1154(w_eco1154, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1155(w_eco1155, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1156(w_eco1156, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_cnt_len[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1157(w_eco1157, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1158(w_eco1158, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1159(w_eco1159, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1160(w_eco1160, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1161(w_eco1161, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1162(w_eco1162, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !rst, !prev_cnt[9], !prev_cnt[13], prev_cnt_len[2], !prev_cnt_len[14]);
	and _ECO_1163(w_eco1163, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1164(w_eco1164, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1165(w_eco1165, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1166(w_eco1166, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1167(w_eco1167, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1168(w_eco1168, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1169(w_eco1169, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1170(w_eco1170, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1171(w_eco1171, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1172(w_eco1172, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1173(w_eco1173, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1174(w_eco1174, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1175(w_eco1175, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1176(w_eco1176, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1177(w_eco1177, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1178(w_eco1178, !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1179(w_eco1179, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1180(w_eco1180, !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_1181(w_eco1181, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !ena, !prev_cnt[0]);
	and _ECO_1182(w_eco1182, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1183(w_eco1183, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1184(w_eco1184, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1185(w_eco1185, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1186(w_eco1186, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1187(w_eco1187, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1188(w_eco1188, !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1189(w_eco1189, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1190(w_eco1190, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1191(w_eco1191, prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1192(w_eco1192, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1193(w_eco1193, prev_state[1], !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1194(w_eco1194, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1195(w_eco1195, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1196(w_eco1196, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1197(w_eco1197, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[11], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1198(w_eco1198, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1199(w_eco1199, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1200(w_eco1200, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1201(w_eco1201, !prev_cnt_len[5], prev_state[1], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1202(w_eco1202, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1203(w_eco1203, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1204(w_eco1204, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[11]);
	and _ECO_1205(w_eco1205, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1206(w_eco1206, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_1207(w_eco1207, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1208(w_eco1208, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst);
	and _ECO_1209(w_eco1209, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1210(w_eco1210, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_1211(w_eco1211, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1212(w_eco1212, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14], prev_cnt[2]);
	and _ECO_1213(w_eco1213, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1214(w_eco1214, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1215(w_eco1215, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1216(w_eco1216, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1217(w_eco1217, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_cnt[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1218(w_eco1218, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1219(w_eco1219, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1220(w_eco1220, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1221(w_eco1221, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1222(w_eco1222, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1223(w_eco1223, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1224(w_eco1224, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !rst, !prev_cnt[2]);
	and _ECO_1225(w_eco1225, !prev_cnt_len[5], prev_cnt_len[15], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1226(w_eco1226, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1227(w_eco1227, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1228(w_eco1228, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1229(w_eco1229, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1230(w_eco1230, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1231(w_eco1231, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1232(w_eco1232, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1233(w_eco1233, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1234(w_eco1234, prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1235(w_eco1235, !prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[13], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1236(w_eco1236, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1237(w_eco1237, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1238(w_eco1238, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1239(w_eco1239, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1240(w_eco1240, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1241(w_eco1241, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1242(w_eco1242, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1243(w_eco1243, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1244(w_eco1244, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1245(w_eco1245, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1246(w_eco1246, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1247(w_eco1247, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1248(w_eco1248, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1249(w_eco1249, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1250(w_eco1250, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1251(w_eco1251, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1252(w_eco1252, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1253(w_eco1253, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1254(w_eco1254, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1255(w_eco1255, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1256(w_eco1256, !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1257(w_eco1257, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1258(w_eco1258, prev_state[1], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1259(w_eco1259, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1260(w_eco1260, !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1261(w_eco1261, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1262(w_eco1262, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1263(w_eco1263, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1264(w_eco1264, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1265(w_eco1265, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1266(w_eco1266, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1267(w_eco1267, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1268(w_eco1268, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1269(w_eco1269, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1270(w_eco1270, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[11]);
	and _ECO_1271(w_eco1271, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_1272(w_eco1272, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, prev_cnt[5]);
	and _ECO_1273(w_eco1273, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst);
	and _ECO_1274(w_eco1274, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_1275(w_eco1275, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1276(w_eco1276, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1277(w_eco1277, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1278(w_eco1278, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1279(w_eco1279, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1280(w_eco1280, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1281(w_eco1281, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1282(w_eco1282, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1283(w_eco1283, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1284(w_eco1284, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1285(w_eco1285, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1286(w_eco1286, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1287(w_eco1287, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1288(w_eco1288, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1289(w_eco1289, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1290(w_eco1290, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1291(w_eco1291, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1292(w_eco1292, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1293(w_eco1293, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1294(w_eco1294, prev_cnt_len[11], prev_state[1], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1295(w_eco1295, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1296(w_eco1296, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1297(w_eco1297, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1298(w_eco1298, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1299(w_eco1299, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8], prev_cnt[2]);
	and _ECO_1300(w_eco1300, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1301(w_eco1301, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1302(w_eco1302, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1303(w_eco1303, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1304(w_eco1304, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1305(w_eco1305, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !ena, !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1306(w_eco1306, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1307(w_eco1307, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1308(w_eco1308, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1309(w_eco1309, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1310(w_eco1310, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1311(w_eco1311, !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1312(w_eco1312, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1313(w_eco1313, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1314(w_eco1314, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1315(w_eco1315, !prev_state[1], !prev_state[3], !prev_cnt[6], prev_cnt[3], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1316(w_eco1316, !prev_state[3], prev_cnt[15], prev_cnt[3], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1317(w_eco1317, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1318(w_eco1318, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1319(w_eco1319, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1320(w_eco1320, prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1321(w_eco1321, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1322(w_eco1322, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1323(w_eco1323, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, prev_cnt[5], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1324(w_eco1324, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1325(w_eco1325, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1326(w_eco1326, !prev_cnt_len[5], prev_cnt_len[15], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1327(w_eco1327, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1328(w_eco1328, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, prev_cnt[5]);
	and _ECO_1329(w_eco1329, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_1330(w_eco1330, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst);
	and _ECO_1331(w_eco1331, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[1], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1332(w_eco1332, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1333(w_eco1333, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1334(w_eco1334, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1335(w_eco1335, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1336(w_eco1336, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1337(w_eco1337, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[3], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1338(w_eco1338, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1339(w_eco1339, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1340(w_eco1340, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1341(w_eco1341, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_state[2], !prev_cnt_len[12], !rst, !prev_cnt[2]);
	and _ECO_1342(w_eco1342, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1343(w_eco1343, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1344(w_eco1344, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1345(w_eco1345, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1346(w_eco1346, !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], prev_cnt_len[3], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1347(w_eco1347, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0], prev_cnt_len[14]);
	and _ECO_1348(w_eco1348, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, prev_cnt_len[2], !prev_cnt_len[14], !prev_cnt[2]);
	and _ECO_1349(w_eco1349, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1350(w_eco1350, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1351(w_eco1351, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1352(w_eco1352, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1353(w_eco1353, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1354(w_eco1354, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1355(w_eco1355, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1356(w_eco1356, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1357(w_eco1357, !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt[2]);
	and _ECO_1358(w_eco1358, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1359(w_eco1359, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1360(w_eco1360, prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1361(w_eco1361, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1362(w_eco1362, prev_state[1], !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1363(w_eco1363, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1364(w_eco1364, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1365(w_eco1365, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1366(w_eco1366, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1367(w_eco1367, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], prev_cnt[14], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst);
	and _ECO_1368(w_eco1368, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1369(w_eco1369, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[4], !prev_cnt_len[12], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1370(w_eco1370, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1371(w_eco1371, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1372(w_eco1372, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_cnt_len[10], !prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1373(w_eco1373, !prev_cnt_len[5], !prev_cnt_len[11], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1374(w_eco1374, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], prev_cnt[6], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1375(w_eco1375, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[12], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[2]);
	and _ECO_1376(w_eco1376, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[8], ena, !prev_cnt[2]);
	and _ECO_1377(w_eco1377, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1378(w_eco1378, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1379(w_eco1379, prev_state[1], !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], !prev_cnt[0]);
	and _ECO_1380(w_eco1380, prev_cnt_len[11], !prev_cnt_len[15], !prev_state[3], !prev_cnt[14], !prev_state[0], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1381(w_eco1381, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1382(w_eco1382, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2], prev_cnt_len[8]);
	and _ECO_1383(w_eco1383, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1384(w_eco1384, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1385(w_eco1385, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1386(w_eco1386, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1387(w_eco1387, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[13], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1388(w_eco1388, !prev_state[1], !prev_state[3], prev_cnt[10], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1389(w_eco1389, !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !rst, !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1390(w_eco1390, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[6], !rst, !prev_cnt[9], !prev_cnt[13], !prev_cnt_len[14], !prev_cnt_len[8]);
	and _ECO_1391(w_eco1391, !prev_cnt_len[5], !prev_cnt_len[11], prev_state[1], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1392(w_eco1392, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_state[3], !prev_cnt[3], !prev_cnt_len[3], !prev_state[0], !prev_cnt_len[0], prev_cnt_len[13], !prev_cnt_len[12], prev_state[4], !rst, !prev_cnt[9], !prev_cnt[13]);
	and _ECO_1393(w_eco1393, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], prev_state[2], !prev_cnt[1], prev_state[4], !rst, !prev_cnt[4], prev_cnt[12], ena, !prev_cnt[2]);
	and _ECO_1394(w_eco1394, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], prev_cnt[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1395(w_eco1395, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_cnt[1], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1396(w_eco1396, !prev_cnt_len[15], !prev_cnt_len[9], !prev_state[3], !prev_cnt[14], !prev_state[0], !prev_cnt_len[7], prev_state[2], !prev_cnt[8], !prev_cnt[12], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], !prev_cnt[0]);
	and _ECO_1397(w_eco1397, !prev_state[1], !prev_state[3], !prev_cnt[6], !prev_cnt[14], !prev_cnt_len[10], !prev_state[2], prev_cnt_len[6], prev_cnt_len[12], prev_cnt[1], prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1398(w_eco1398, !prev_state[3], prev_cnt[15], !prev_cnt[14], !prev_state[0], !prev_cnt_len[4], !prev_cnt_len[10], !prev_state[2], !prev_cnt_len[1], prev_cnt_len[6], !prev_state[4], !prev_cnt[5], prev_cnt[9], !prev_cnt[7], prev_cnt[11], ena, !prev_cnt[0], !prev_cnt_len[2]);
	and _ECO_1399(w_eco1399, !prev_cnt_len[5], !prev_cnt_len[11], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[7], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	and _ECO_1400(w_eco1400, !prev_cnt_len[5], !prev_cnt_len[11], prev_cnt_len[9], !prev_cnt[10], !prev_cnt[15], !prev_cnt_len[3], !prev_cnt_len[0], prev_cnt_len[13], !prev_state[2], !prev_cnt_len[6], !prev_cnt[1], prev_state[4], !rst, !prev_cnt_len[14], !prev_cnt_len[8], !prev_cnt[2]);
	or _ECO_1401(w_eco1401, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462, w_eco463, w_eco464, w_eco465, w_eco466, w_eco467, w_eco468, w_eco469, w_eco470, w_eco471, w_eco472, w_eco473, w_eco474, w_eco475, w_eco476, w_eco477, w_eco478, w_eco479, w_eco480, w_eco481, w_eco482, w_eco483, w_eco484, w_eco485, w_eco486, w_eco487, w_eco488, w_eco489, w_eco490, w_eco491, w_eco492, w_eco493, w_eco494, w_eco495, w_eco496, w_eco497, w_eco498, w_eco499, w_eco500, w_eco501, w_eco502, w_eco503, w_eco504, w_eco505, w_eco506, w_eco507, w_eco508, w_eco509, w_eco510, w_eco511, w_eco512, w_eco513, w_eco514, w_eco515, w_eco516, w_eco517, w_eco518, w_eco519, w_eco520, w_eco521, w_eco522, w_eco523, w_eco524, w_eco525, w_eco526, w_eco527, w_eco528, w_eco529, w_eco530, w_eco531, w_eco532, w_eco533, w_eco534, w_eco535, w_eco536, w_eco537, w_eco538, w_eco539, w_eco540, w_eco541, w_eco542, w_eco543, w_eco544, w_eco545, w_eco546, w_eco547, w_eco548, w_eco549, w_eco550, w_eco551, w_eco552, w_eco553, w_eco554, w_eco555, w_eco556, w_eco557, w_eco558, w_eco559, w_eco560, w_eco561, w_eco562, w_eco563, w_eco564, w_eco565, w_eco566, w_eco567, w_eco568, w_eco569, w_eco570, w_eco571, w_eco572, w_eco573, w_eco574, w_eco575, w_eco576, w_eco577, w_eco578, w_eco579, w_eco580, w_eco581, w_eco582, w_eco583, w_eco584, w_eco585, w_eco586, w_eco587, w_eco588, w_eco589, w_eco590, w_eco591, w_eco592, w_eco593, w_eco594, w_eco595, w_eco596, w_eco597, w_eco598, w_eco599, w_eco600, w_eco601, w_eco602, w_eco603, w_eco604, w_eco605, w_eco606, w_eco607, w_eco608, w_eco609, w_eco610, w_eco611, w_eco612, w_eco613, w_eco614, w_eco615, w_eco616, w_eco617, w_eco618, w_eco619, w_eco620, w_eco621, w_eco622, w_eco623, w_eco624, w_eco625, w_eco626, w_eco627, w_eco628, w_eco629, w_eco630, w_eco631, w_eco632, w_eco633, w_eco634, w_eco635, w_eco636, w_eco637, w_eco638, w_eco639, w_eco640, w_eco641, w_eco642, w_eco643, w_eco644, w_eco645, w_eco646, w_eco647, w_eco648, w_eco649, w_eco650, w_eco651, w_eco652, w_eco653, w_eco654, w_eco655, w_eco656, w_eco657, w_eco658, w_eco659, w_eco660, w_eco661, w_eco662, w_eco663, w_eco664, w_eco665, w_eco666, w_eco667, w_eco668, w_eco669, w_eco670, w_eco671, w_eco672, w_eco673, w_eco674, w_eco675, w_eco676, w_eco677, w_eco678, w_eco679, w_eco680, w_eco681, w_eco682, w_eco683, w_eco684, w_eco685, w_eco686, w_eco687, w_eco688, w_eco689, w_eco690, w_eco691, w_eco692, w_eco693, w_eco694, w_eco695, w_eco696, w_eco697, w_eco698, w_eco699, w_eco700, w_eco701, w_eco702, w_eco703, w_eco704, w_eco705, w_eco706, w_eco707, w_eco708, w_eco709, w_eco710, w_eco711, w_eco712, w_eco713, w_eco714, w_eco715, w_eco716, w_eco717, w_eco718, w_eco719, w_eco720, w_eco721, w_eco722, w_eco723, w_eco724, w_eco725, w_eco726, w_eco727, w_eco728, w_eco729, w_eco730, w_eco731, w_eco732, w_eco733, w_eco734, w_eco735, w_eco736, w_eco737, w_eco738, w_eco739, w_eco740, w_eco741, w_eco742, w_eco743, w_eco744, w_eco745, w_eco746, w_eco747, w_eco748, w_eco749, w_eco750, w_eco751, w_eco752, w_eco753, w_eco754, w_eco755, w_eco756, w_eco757, w_eco758, w_eco759, w_eco760, w_eco761, w_eco762, w_eco763, w_eco764, w_eco765, w_eco766, w_eco767, w_eco768, w_eco769, w_eco770, w_eco771, w_eco772, w_eco773, w_eco774, w_eco775, w_eco776, w_eco777, w_eco778, w_eco779, w_eco780, w_eco781, w_eco782, w_eco783, w_eco784, w_eco785, w_eco786, w_eco787, w_eco788, w_eco789, w_eco790, w_eco791, w_eco792, w_eco793, w_eco794, w_eco795, w_eco796, w_eco797, w_eco798, w_eco799, w_eco800, w_eco801, w_eco802, w_eco803, w_eco804, w_eco805, w_eco806, w_eco807, w_eco808, w_eco809, w_eco810, w_eco811, w_eco812, w_eco813, w_eco814, w_eco815, w_eco816, w_eco817, w_eco818, w_eco819, w_eco820, w_eco821, w_eco822, w_eco823, w_eco824, w_eco825, w_eco826, w_eco827, w_eco828, w_eco829, w_eco830, w_eco831, w_eco832, w_eco833, w_eco834, w_eco835, w_eco836, w_eco837, w_eco838, w_eco839, w_eco840, w_eco841, w_eco842, w_eco843, w_eco844, w_eco845, w_eco846, w_eco847, w_eco848, w_eco849, w_eco850, w_eco851, w_eco852, w_eco853, w_eco854, w_eco855, w_eco856, w_eco857, w_eco858, w_eco859, w_eco860, w_eco861, w_eco862, w_eco863, w_eco864, w_eco865, w_eco866, w_eco867, w_eco868, w_eco869, w_eco870, w_eco871, w_eco872, w_eco873, w_eco874, w_eco875, w_eco876, w_eco877, w_eco878, w_eco879, w_eco880, w_eco881, w_eco882, w_eco883, w_eco884, w_eco885, w_eco886, w_eco887, w_eco888, w_eco889, w_eco890, w_eco891, w_eco892, w_eco893, w_eco894, w_eco895, w_eco896, w_eco897, w_eco898, w_eco899, w_eco900, w_eco901, w_eco902, w_eco903, w_eco904, w_eco905, w_eco906, w_eco907, w_eco908, w_eco909, w_eco910, w_eco911, w_eco912, w_eco913, w_eco914, w_eco915, w_eco916, w_eco917, w_eco918, w_eco919, w_eco920, w_eco921, w_eco922, w_eco923, w_eco924, w_eco925, w_eco926, w_eco927, w_eco928, w_eco929, w_eco930, w_eco931, w_eco932, w_eco933, w_eco934, w_eco935, w_eco936, w_eco937, w_eco938, w_eco939, w_eco940, w_eco941, w_eco942, w_eco943, w_eco944, w_eco945, w_eco946, w_eco947, w_eco948, w_eco949, w_eco950, w_eco951, w_eco952, w_eco953, w_eco954, w_eco955, w_eco956, w_eco957, w_eco958, w_eco959, w_eco960, w_eco961, w_eco962, w_eco963, w_eco964, w_eco965, w_eco966, w_eco967, w_eco968, w_eco969, w_eco970, w_eco971, w_eco972, w_eco973, w_eco974, w_eco975, w_eco976, w_eco977, w_eco978, w_eco979, w_eco980, w_eco981, w_eco982, w_eco983, w_eco984, w_eco985, w_eco986, w_eco987, w_eco988, w_eco989, w_eco990, w_eco991, w_eco992, w_eco993, w_eco994, w_eco995, w_eco996, w_eco997, w_eco998, w_eco999, w_eco1000, w_eco1001, w_eco1002, w_eco1003, w_eco1004, w_eco1005, w_eco1006, w_eco1007, w_eco1008, w_eco1009, w_eco1010, w_eco1011, w_eco1012, w_eco1013, w_eco1014, w_eco1015, w_eco1016, w_eco1017, w_eco1018, w_eco1019, w_eco1020, w_eco1021, w_eco1022, w_eco1023, w_eco1024, w_eco1025, w_eco1026, w_eco1027, w_eco1028, w_eco1029, w_eco1030, w_eco1031, w_eco1032, w_eco1033, w_eco1034, w_eco1035, w_eco1036, w_eco1037, w_eco1038, w_eco1039, w_eco1040, w_eco1041, w_eco1042, w_eco1043, w_eco1044, w_eco1045, w_eco1046, w_eco1047, w_eco1048, w_eco1049, w_eco1050, w_eco1051, w_eco1052, w_eco1053, w_eco1054, w_eco1055, w_eco1056, w_eco1057, w_eco1058, w_eco1059, w_eco1060, w_eco1061, w_eco1062, w_eco1063, w_eco1064, w_eco1065, w_eco1066, w_eco1067, w_eco1068, w_eco1069, w_eco1070, w_eco1071, w_eco1072, w_eco1073, w_eco1074, w_eco1075, w_eco1076, w_eco1077, w_eco1078, w_eco1079, w_eco1080, w_eco1081, w_eco1082, w_eco1083, w_eco1084, w_eco1085, w_eco1086, w_eco1087, w_eco1088, w_eco1089, w_eco1090, w_eco1091, w_eco1092, w_eco1093, w_eco1094, w_eco1095, w_eco1096, w_eco1097, w_eco1098, w_eco1099, w_eco1100, w_eco1101, w_eco1102, w_eco1103, w_eco1104, w_eco1105, w_eco1106, w_eco1107, w_eco1108, w_eco1109, w_eco1110, w_eco1111, w_eco1112, w_eco1113, w_eco1114, w_eco1115, w_eco1116, w_eco1117, w_eco1118, w_eco1119, w_eco1120, w_eco1121, w_eco1122, w_eco1123, w_eco1124, w_eco1125, w_eco1126, w_eco1127, w_eco1128, w_eco1129, w_eco1130, w_eco1131, w_eco1132, w_eco1133, w_eco1134, w_eco1135, w_eco1136, w_eco1137, w_eco1138, w_eco1139, w_eco1140, w_eco1141, w_eco1142, w_eco1143, w_eco1144, w_eco1145, w_eco1146, w_eco1147, w_eco1148, w_eco1149, w_eco1150, w_eco1151, w_eco1152, w_eco1153, w_eco1154, w_eco1155, w_eco1156, w_eco1157, w_eco1158, w_eco1159, w_eco1160, w_eco1161, w_eco1162, w_eco1163, w_eco1164, w_eco1165, w_eco1166, w_eco1167, w_eco1168, w_eco1169, w_eco1170, w_eco1171, w_eco1172, w_eco1173, w_eco1174, w_eco1175, w_eco1176, w_eco1177, w_eco1178, w_eco1179, w_eco1180, w_eco1181, w_eco1182, w_eco1183, w_eco1184, w_eco1185, w_eco1186, w_eco1187, w_eco1188, w_eco1189, w_eco1190, w_eco1191, w_eco1192, w_eco1193, w_eco1194, w_eco1195, w_eco1196, w_eco1197, w_eco1198, w_eco1199, w_eco1200, w_eco1201, w_eco1202, w_eco1203, w_eco1204, w_eco1205, w_eco1206, w_eco1207, w_eco1208, w_eco1209, w_eco1210, w_eco1211, w_eco1212, w_eco1213, w_eco1214, w_eco1215, w_eco1216, w_eco1217, w_eco1218, w_eco1219, w_eco1220, w_eco1221, w_eco1222, w_eco1223, w_eco1224, w_eco1225, w_eco1226, w_eco1227, w_eco1228, w_eco1229, w_eco1230, w_eco1231, w_eco1232, w_eco1233, w_eco1234, w_eco1235, w_eco1236, w_eco1237, w_eco1238, w_eco1239, w_eco1240, w_eco1241, w_eco1242, w_eco1243, w_eco1244, w_eco1245, w_eco1246, w_eco1247, w_eco1248, w_eco1249, w_eco1250, w_eco1251, w_eco1252, w_eco1253, w_eco1254, w_eco1255, w_eco1256, w_eco1257, w_eco1258, w_eco1259, w_eco1260, w_eco1261, w_eco1262, w_eco1263, w_eco1264, w_eco1265, w_eco1266, w_eco1267, w_eco1268, w_eco1269, w_eco1270, w_eco1271, w_eco1272, w_eco1273, w_eco1274, w_eco1275, w_eco1276, w_eco1277, w_eco1278, w_eco1279, w_eco1280, w_eco1281, w_eco1282, w_eco1283, w_eco1284, w_eco1285, w_eco1286, w_eco1287, w_eco1288, w_eco1289, w_eco1290, w_eco1291, w_eco1292, w_eco1293, w_eco1294, w_eco1295, w_eco1296, w_eco1297, w_eco1298, w_eco1299, w_eco1300, w_eco1301, w_eco1302, w_eco1303, w_eco1304, w_eco1305, w_eco1306, w_eco1307, w_eco1308, w_eco1309, w_eco1310, w_eco1311, w_eco1312, w_eco1313, w_eco1314, w_eco1315, w_eco1316, w_eco1317, w_eco1318, w_eco1319, w_eco1320, w_eco1321, w_eco1322, w_eco1323, w_eco1324, w_eco1325, w_eco1326, w_eco1327, w_eco1328, w_eco1329, w_eco1330, w_eco1331, w_eco1332, w_eco1333, w_eco1334, w_eco1335, w_eco1336, w_eco1337, w_eco1338, w_eco1339, w_eco1340, w_eco1341, w_eco1342, w_eco1343, w_eco1344, w_eco1345, w_eco1346, w_eco1347, w_eco1348, w_eco1349, w_eco1350, w_eco1351, w_eco1352, w_eco1353, w_eco1354, w_eco1355, w_eco1356, w_eco1357, w_eco1358, w_eco1359, w_eco1360, w_eco1361, w_eco1362, w_eco1363, w_eco1364, w_eco1365, w_eco1366, w_eco1367, w_eco1368, w_eco1369, w_eco1370, w_eco1371, w_eco1372, w_eco1373, w_eco1374, w_eco1375, w_eco1376, w_eco1377, w_eco1378, w_eco1379, w_eco1380, w_eco1381, w_eco1382, w_eco1383, w_eco1384, w_eco1385, w_eco1386, w_eco1387, w_eco1388, w_eco1389, w_eco1390, w_eco1391, w_eco1392, w_eco1393, w_eco1394, w_eco1395, w_eco1396, w_eco1397, w_eco1398, w_eco1399, w_eco1400);
	xor _ECO_out2(Gate, sub_wire2, w_eco1401);

endmodule