module ex_or(yor, a, b);
  input a, b;
  output yor;
  wire a, b;
  wire yor;
  or g1 (yor, a, b);
endmodule

