module top(a_gtet_b,a,b);
	input [7:0]a, b;
	output a_gtet_b;
	wire [7:0]a, b;
	wire a_gtet_b, n_8, n_13, n_43, n_52, n_59, n_64, n_67, n_149, n_156, n_158, n_171, n_403, n_407, n_410, n_415, n_425, n_432, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517, n_518, n_519, n_520, n_521, n_522, n_523, n_524;
	wire sub_wire0, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461, w_eco462;

	nand g47(n_52, n_8, a[2]);
	nand g58(n_149, n_485, n_496);
	nor g133(n_158, n_43, a[1]);
	not g468(n_442, a[2]);
	not g469(n_443, a[1]);
	not g470(n_444, b[2]);
	not g471(n_445, b[5]);
	not g472(n_446, a[5]);
	not g473(n_447, b[7]);
	not g474(n_448, a[7]);
	not g475(n_449, a[3]);
	not g476(n_450, b[4]);
	not g477(n_451, a[4]);
	not g478(n_452, b[6]);
	not g479(n_453, a[6]);
	not g480(n_454, b[1]);
	not g481(n_455, a[0]);
	nand g482(n_8, n_449, b[3]);
	not g483(n_456, n_8);
	nand g484(n_13, a[7], n_447);
	not g485(n_457, n_13);
	nor g486(n_458, a[6], n_452);
	not g487(n_459, n_458);
	nor g488(n_407, n_442, b[2]);
	not g489(n_460, n_407);
	nor g490(n_43, n_449, b[3]);
	not g491(n_461, n_43);
	not g492(n_462, n_158);
	nor g493(n_463, n_43, n_454);
	not g494(n_464, n_463);
	nand g495(n_465, n_462, n_464);
	nand g496(n_466, n_460, n_465, b[0]);
	nor g497(n_403, a[2], n_444);
	not g498(n_467, n_403);
	nand g499(n_410, n_467, n_8, n_454);
	not g500(n_468, n_410);
	nand g501(n_469, n_460, n_461, n_443);
	nor g502(n_470, n_468, n_469);
	not g503(n_471, n_470);
	nor g504(n_472, n_456, n_461);
	not g505(n_473, n_472);
	nor g506(n_474, n_456, b[2]);
	not g507(n_475, n_474);
	nand g508(n_476, n_52, n_473, n_475);
	nor g509(n_477, n_468, n_476);
	not g510(n_478, n_477);
	nand g511(n_59, n_466, n_471, n_478);
	not g512(n_479, n_59);
	nor g513(n_480, n_59, n_451);
	not g514(n_481, n_480);
	nor g515(n_482, n_479, a[4]);
	not g516(n_483, n_482);
	nand g517(n_484, n_483, n_450);
	nand g518(n_64, n_481, n_484);
	nand g519(n_485, n_13, n_459, n_64);
	nand g520(n_67, n_448, b[7]);
	not g521(n_486, n_67);
	nor g522(n_487, n_453, b[6]);
	not g523(n_488, n_487);
	nand g524(n_489, n_67, n_488, n_446);
	nor g525(n_415, n_486, a[6]);
	not g526(n_490, n_415);
	nand g527(n_425, n_13, n_490);
	not g528(n_491, n_425);
	nor g529(n_492, n_13, n_491);
	not g530(n_493, n_492);
	nor g531(n_494, n_491, n_452);
	not g532(n_495, n_494);
	nand g533(n_496, n_489, n_493, n_495);
	nor g534(n_497, a[5], n_445);
	not g535(n_498, n_497);
	nand g536(n_156, n_467, n_498);
	nor g537(n_499, n_156, n_453, n_455);
	not g538(n_500, n_499);
	nor g539(n_501, n_156, n_455, b[6]);
	not g540(n_502, n_501);
	nand g541(n_503, n_500, n_502);
	not g542(n_504, n_503);
	nor g543(n_505, a[4], n_450);
	not g544(n_506, n_505);
	nand g545(n_171, n_8, n_506);
	nor g546(n_507, n_457, n_171, n_443);
	not g547(n_508, n_507);
	nor g548(n_509, n_457, n_171, b[1]);
	not g549(n_510, n_509);
	nand g550(n_511, n_508, n_510);
	not g551(n_512, n_511);
	nor g552(n_513, n_504, n_512);
	not g553(n_514, n_513);
	nor g554(n_515, n_486, n_452, n_445);
	not g555(n_516, n_515);
	nor g556(n_517, n_490, n_445);
	not g557(n_518, n_517);
	nand g558(n_432, n_516, n_518);
	not g559(n_519, n_432);
	nor g560(n_520, n_519, a[5]);
	not g561(n_521, n_520);
	nor g562(n_522, n_519, n_64);
	not g563(n_523, n_522);
	nand g564(n_524, n_149, n_521, n_523);
	nand g565(sub_wire0, n_514, n_524);
	and _ECO_0(w_eco0, a[2], !a[1], b[2], !b[5], a[5], b[7], b[4]);
	and _ECO_1(w_eco1, !a[1], b[2], !b[5], a[5], b[7], !a[3], b[4]);
	and _ECO_2(w_eco2, !a[2], !a[1], !b[5], a[5], b[7], !a[3], b[4]);
	and _ECO_3(w_eco3, a[2], b[2], !b[5], a[5], b[7], a[3], b[4], !b[1]);
	and _ECO_4(w_eco4, a[2], !a[1], b[2], !b[5], a[5], b[7], !a[4]);
	and _ECO_5(w_eco5, a[2], !a[1], b[2], !b[5], a[7], b[4], b[6]);
	and _ECO_6(w_eco6, a[2], !a[1], b[2], !b[5], a[5], !a[7], b[4]);
	and _ECO_7(w_eco7, a[2], !a[1], !b[2], b[5], !a[5], b[7], a[3], !b[4]);
	and _ECO_8(w_eco8, a[2], !a[1], !b[2], b[5], !a[5], !a[7], a[3], !b[4]);
	and _ECO_9(w_eco9, !a[1], !b[5], a[5], b[7], b[4], !a[4]);
	and _ECO_10(w_eco10, !a[1], !b[5], a[5], b[7], !b[6]);
	and _ECO_11(w_eco11, !a[1], b[2], !b[5], a[5], !a[7], !a[3], b[4]);
	and _ECO_12(w_eco12, !a[2], !a[1], !b[5], a[5], !a[7], !a[3], b[4]);
	and _ECO_13(w_eco13, b[2], !b[5], a[5], b[7], b[4], b[1], !a[0]);
	and _ECO_14(w_eco14, a[2], b[2], !b[5], a[5], b[7], a[3], !a[4], !b[1]);
	and _ECO_15(w_eco15, !b[5], a[5], b[7], b[4], !a[4], !b[1]);
	and _ECO_16(w_eco16, a[2], b[2], !b[5], a[5], !a[7], a[3], b[4], !b[1]);
	and _ECO_17(w_eco17, a[2], !a[1], b[2], a[7], b[4], b[6], a[6]);
	and _ECO_18(w_eco18, !a[1], b[5], !a[5], b[7], !b[4], a[4]);
	and _ECO_19(w_eco19, b[5], !a[5], !b[7], a[7], !b[6], !b[1]);
	and _ECO_20(w_eco20, !a[1], b[5], !a[5], !a[7], !b[4], a[4]);
	and _ECO_21(w_eco21, a[2], !a[1], b[2], !b[5], a[7], !a[4], b[6]);
	and _ECO_22(w_eco22, a[2], !a[1], b[2], !b[5], a[5], !a[7], !a[4]);
	and _ECO_23(w_eco23, a[2], !a[1], !b[2], a[5], b[7], a[3], !b[4], !b[6]);
	and _ECO_24(w_eco24, a[2], !a[1], !b[2], a[5], !a[7], a[3], !b[4], !b[6]);
	and _ECO_25(w_eco25, a[2], !a[1], !b[2], b[5], !a[5], b[7], a[3], a[4]);
	and _ECO_26(w_eco26, a[2], !a[1], !b[2], b[5], !a[5], !a[7], a[3], a[4]);
	and _ECO_27(w_eco27, !a[1], !b[5], a[5], b[7], a[6]);
	and _ECO_28(w_eco28, !a[1], !b[5], a[5], !a[7], b[4], !a[4]);
	and _ECO_29(w_eco29, !a[2], b[2], !b[5], a[7], b[4], !a[4], !b[1]);
	and _ECO_30(w_eco30, !a[1], b[2], !b[5], a[5], !a[7], !a[3], !a[4]);
	and _ECO_31(w_eco31, !a[2], !a[1], !b[5], a[7], !a[3], b[4], b[6]);
	and _ECO_32(w_eco32, !a[2], !a[1], !b[5], a[5], !a[7], !a[3], !a[4]);
	and _ECO_33(w_eco33, b[5], !a[5], b[7], !b[4], a[4], !b[1]);
	and _ECO_34(w_eco34, b[5], !a[5], !a[7], !b[4], a[4], !b[1]);
	and _ECO_35(w_eco35, b[2], !b[5], a[5], b[7], b[4], !b[0]);
	and _ECO_36(w_eco36, a[5], b[7], !b[4], a[4], !b[6], !b[1]);
	and _ECO_37(w_eco37, b[2], !b[5], a[5], b[7], !a[4], b[1], !a[0]);
	and _ECO_38(w_eco38, !b[5], a[5], b[7], !b[6], !b[1]);
	and _ECO_39(w_eco39, a[2], b[2], !b[5], a[7], a[3], b[4], b[6], !b[1]);
	and _ECO_40(w_eco40, b[2], !b[5], a[5], !a[7], b[4], b[1], !a[0]);
	and _ECO_41(w_eco41, a[2], b[2], !b[5], a[5], !a[7], a[3], !a[4], !b[1]);
	and _ECO_42(w_eco42, !b[5], a[5], !a[7], b[4], !a[4], !b[1]);
	and _ECO_43(w_eco43, !b[5], a[5], b[7], b[4], !a[4], !a[0]);
	and _ECO_44(w_eco44, !b[5], a[7], b[4], !a[4], b[6], !b[1]);
	and _ECO_45(w_eco45, !b[7], a[7], !b[6], !a[6], !b[1]);
	and _ECO_46(w_eco46, a[2], !a[1], b[2], a[7], !a[4], b[6], a[6]);
	and _ECO_47(w_eco47, !a[1], a[5], b[7], !b[4], a[4], a[6]);
	and _ECO_48(w_eco48, !b[7], a[7], !a[6], !b[1], a[0]);
	and _ECO_49(w_eco49, !b[7], a[7], !b[6], !b[1], !a[0]);
	and _ECO_50(w_eco50, !a[1], a[5], !a[7], !b[4], a[4], !b[6]);
	and _ECO_51(w_eco51, !a[1], !b[7], !a[7], b[6], a[6]);
	and _ECO_52(w_eco52, !a[1], b[5], !a[5], !b[4], a[4], !b[6]);
	and _ECO_53(w_eco53, a[2], !a[1], b[2], !b[5], !b[7], !a[7], b[4], !a[6]);
	and _ECO_54(w_eco54, a[2], !a[1], b[2], !b[5], !b[7], !a[7], !a[4], !a[6]);
	and _ECO_55(w_eco55, a[2], !a[1], !b[2], a[5], b[7], a[3], a[4], !b[6]);
	and _ECO_56(w_eco56, a[2], !a[1], !b[2], a[5], !a[7], a[3], a[4], !b[6]);
	and _ECO_57(w_eco57, a[2], !a[1], !b[2], b[5], !a[5], a[4], !b[6]);
	and _ECO_58(w_eco58, a[2], !a[1], !b[2], b[5], !a[5], !b[4], !b[6]);
	and _ECO_59(w_eco59, !a[1], !b[5], a[5], !a[7], !b[6]);
	and _ECO_60(w_eco60, !a[1], b[7], a[7], b[6], a[6]);
	and _ECO_61(w_eco61, !a[1], !b[5], b[7], a[7], !b[6], !a[6]);
	and _ECO_62(w_eco62, !a[1], !b[5], !b[7], !a[7], !b[6], !a[6]);
	and _ECO_63(w_eco63, a[1], !b[5], a[7], b[4], !a[4], !a[0]);
	and _ECO_64(w_eco64, !a[2], b[2], !b[5], !b[7], b[4], !a[4], !b[1]);
	and _ECO_65(w_eco65, !a[1], b[2], a[7], !a[3], b[4], b[6], a[6]);
	and _ECO_66(w_eco66, !a[2], !a[1], a[7], !a[3], b[4], b[6], a[6]);
	and _ECO_67(w_eco67, !a[1], !b[2], b[5], !a[5], !a[7], a[3], a[4], !b[3]);
	and _ECO_68(w_eco68, !a[1], !b[2], b[5], !a[5], !a[7], a[3], !b[4], !b[3]);
	and _ECO_69(w_eco69, a[2], b[2], a[7], a[3], b[4], b[6], a[6], !b[1]);
	and _ECO_70(w_eco70, a[5], !a[7], !b[4], a[4], !b[6], !b[1]);
	and _ECO_71(w_eco71, b[5], !a[5], b[4], !a[4], !b[6], !b[1]);
	and _ECO_72(w_eco72, b[5], !a[5], b[7], !b[4], a[4], !a[0]);
	and _ECO_73(w_eco73, a[1], !b[7], a[7], !b[6], !a[0]);
	and _ECO_74(w_eco74, b[5], !a[5], !a[7], !b[4], a[4], !a[0]);
	and _ECO_75(w_eco75, a[5], b[7], !b[4], a[4], a[6], !b[1]);
	and _ECO_76(w_eco76, a[5], b[7], !b[4], a[4], !b[6], !a[0]);
	and _ECO_77(w_eco77, b[2], !b[5], a[5], b[7], !a[4], !b[0]);
	and _ECO_78(w_eco78, b[2], !b[5], a[5], !a[7], b[4], !b[0]);
	and _ECO_79(w_eco79, b[2], !b[5], a[5], !a[7], !a[4], b[1], !a[0]);
	and _ECO_80(w_eco80, !b[5], a[5], !a[7], !b[6], !b[1]);
	and _ECO_81(w_eco81, a[2], b[2], !b[5], a[7], a[3], !a[4], b[6], !b[1]);
	and _ECO_82(w_eco82, a[1], !b[5], !a[5], b[7], !a[7], a[3], !b[4], b[1], a[0], b[0]);
	and _ECO_83(w_eco83, a[2], b[2], !b[5], !b[7], a[3], b[4], b[6], !b[1]);
	and _ECO_84(w_eco84, a[2], b[2], !b[5], !b[7], a[3], !a[4], b[6], !b[1]);
	and _ECO_85(w_eco85, !b[5], !b[7], b[4], !a[4], b[6], !b[1]);
	and _ECO_86(w_eco86, a[7], b[4], !a[4], b[6], a[6], !b[1]);
	and _ECO_87(w_eco87, a[1], !b[2], b[5], !a[5], !a[7], a[4], !b[1], b[0]);
	and _ECO_88(w_eco88, a[1], !b[2], b[5], !a[5], !a[7], !b[4], !b[1], b[0]);
	and _ECO_89(w_eco89, !b[5], a[5], b[7], a[6], !b[1]);
	and _ECO_90(w_eco90, !b[5], a[5], b[7], !b[6], !a[0]);
	and _ECO_91(w_eco91, !b[5], a[5], b[7], b[4], !a[4], !b[0]);
	and _ECO_92(w_eco92, !b[5], a[5], !a[7], b[4], !a[4], !a[0]);
	and _ECO_93(w_eco93, !a[1], b[5], !a[5], !b[4], a[4], !a[6]);
	and _ECO_94(w_eco94, a[2], !a[1], !b[2], b[7], a[7], a[4], !b[6], !a[6]);
	and _ECO_95(w_eco95, a[2], !a[1], !b[2], b[7], a[7], !b[4], !b[6], !a[6]);
	and _ECO_96(w_eco96, a[2], !a[1], !b[2], a[5], !a[7], a[3], a[4], a[6]);
	and _ECO_97(w_eco97, a[2], !a[1], !b[2], a[5], !a[7], a[3], !b[4], a[6]);
	and _ECO_98(w_eco98, a[2], !a[1], !b[2], a[5], !a[7], a[4], !b[6], !a[6]);
	and _ECO_99(w_eco99, a[2], !a[1], !b[2], a[5], !a[7], !b[4], !b[6], !a[6]);
	and _ECO_100(w_eco100, a[2], !a[1], !b[2], b[5], !a[5], !a[7], a[4], b[1]);
	and _ECO_101(w_eco101, a[2], !a[1], !b[2], b[5], !a[5], !a[7], !b[4], b[1]);
	and _ECO_102(w_eco102, !a[1], !b[5], a[7], b[4], !a[4], b[6]);
	and _ECO_103(w_eco103, !a[2], b[2], b[4], !a[4], !b[6], !b[1]);
	and _ECO_104(w_eco104, !a[2], b[2], !b[7], a[7], !b[1], a[0]);
	and _ECO_105(w_eco105, !a[2], a[1], b[2], !b[7], a[7], a[0], !b[0]);
	and _ECO_106(w_eco106, !a[2], a[1], b[5], !a[5], !a[7], a[4], !b[1], b[0]);
	and _ECO_107(w_eco107, !a[2], a[1], b[5], !a[5], !a[7], !b[4], !b[1], b[0]);
	and _ECO_108(w_eco108, b[5], !a[5], !b[4], a[4], !a[6], !a[0]);
	and _ECO_109(w_eco109, b[2], !b[5], a[7], b[4], b[6], b[1], !a[0]);
	and _ECO_110(w_eco110, b[2], !b[5], a[7], !a[4], b[6], b[1], !a[0]);
	and _ECO_111(w_eco111, !a[2], b[2], !a[3], !b[6], !b[1], b[3]);
	and _ECO_112(w_eco112, a[1], !b[5], !b[7], b[4], !a[4], !a[0]);
	and _ECO_113(w_eco113, !a[1], b[2], !b[5], !b[7], !a[3], b[4], b[6]);
	and _ECO_114(w_eco114, !a[1], b[2], !b[5], !b[7], !a[3], !a[4], b[6]);
	and _ECO_115(w_eco115, !a[1], !b[2], a[5], b[7], a[3], a[4], !b[6], !b[3]);
	and _ECO_116(w_eco116, !a[1], !b[2], a[5], b[7], a[3], !b[4], !b[6], !b[3]);
	and _ECO_117(w_eco117, !a[2], !a[1], a[7], !a[3], !a[4], b[6], a[6]);
	and _ECO_118(w_eco118, !a[1], !b[2], a[5], !a[7], a[3], a[4], !b[6], !b[3]);
	and _ECO_119(w_eco119, !a[1], !b[2], a[5], !a[7], a[3], !b[4], !b[6], !b[3]);
	and _ECO_120(w_eco120, !a[1], !b[2], b[5], b[7], a[3], a[4], !b[6], !b[3]);
	and _ECO_121(w_eco121, !a[1], !b[2], b[5], b[7], a[3], !b[4], !b[6], !b[3]);
	and _ECO_122(w_eco122, !a[2], !a[1], !b[5], a[7], !a[3], !a[4], b[6]);
	and _ECO_123(w_eco123, !a[2], !a[1], !b[5], a[5], b[4], b[6], b[3]);
	and _ECO_124(w_eco124, !a[2], !a[1], !b[5], a[5], !a[4], b[6], b[3]);
	and _ECO_125(w_eco125, !a[2], !a[1], !b[5], !b[7], !a[3], b[4], b[6]);
	and _ECO_126(w_eco126, !a[2], !a[1], !b[5], !b[7], !a[3], !a[4], b[6]);
	and _ECO_127(w_eco127, b[4], !a[4], !b[6], !a[6], !b[1]);
	and _ECO_128(w_eco128, b[7], a[7], b[6], a[6], !b[1]);
	and _ECO_129(w_eco129, a[1], b[2], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], a[0], b[0]);
	and _ECO_130(w_eco130, a[1], b[2], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], a[0], b[0]);
	and _ECO_131(w_eco131, b[2], a[7], b[4], b[6], a[6], b[1], !a[0]);
	and _ECO_132(w_eco132, a[1], b[5], !a[5], !b[7], a[7], a[0], !b[0]);
	and _ECO_133(w_eco133, a[1], !b[7], a[7], b[4], b[6], a[0], !b[0]);
	and _ECO_134(w_eco134, a[2], b[2], a[7], a[3], !a[4], b[6], a[6], !b[1]);
	and _ECO_135(w_eco135, !b[7], !a[7], b[6], a[6], !b[1]);
	and _ECO_136(w_eco136, a[5], !a[7], !b[4], a[4], !b[6], !a[0]);
	and _ECO_137(w_eco137, a[1], b[4], !a[4], !b[6], !a[0]);
	and _ECO_138(w_eco138, b[5], !a[5], b[7], !b[4], a[4], !b[0]);
	and _ECO_139(w_eco139, b[5], !a[5], !a[3], !b[6], !b[1], b[3]);
	and _ECO_140(w_eco140, b[5], !a[5], b[4], !a[4], !b[1], a[0]);
	and _ECO_141(w_eco141, a[1], b[5], !a[5], b[4], !a[4], a[0], !b[0]);
	and _ECO_142(w_eco142, b[5], !a[5], !a[7], !b[4], a[4], !b[0]);
	and _ECO_143(w_eco143, a[5], b[7], !b[4], a[4], a[6], !a[0]);
	and _ECO_144(w_eco144, a[5], b[7], !b[4], a[4], !b[6], !b[0]);
	and _ECO_145(w_eco145, b[2], !b[5], a[5], !a[7], !a[4], !b[0]);
	and _ECO_146(w_eco146, !b[5], a[7], !b[6], !a[6], !b[1]);
	and _ECO_147(w_eco147, a[1], !b[5], !a[5], b[7], !a[7], a[3], a[4], b[1], a[0], b[0]);
	and _ECO_148(w_eco148, !a[3], !b[6], !a[6], !b[1], b[3]);
	and _ECO_149(w_eco149, b[2], !b[5], !b[7], b[4], b[6], b[1], !a[0]);
	and _ECO_150(w_eco150, !b[5], !b[7], !b[6], !a[6], !b[1]);
	and _ECO_151(w_eco151, b[2], !b[5], !b[7], !a[4], b[6], b[1], !a[0]);
	and _ECO_152(w_eco152, a[1], !b[2], a[5], b[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_153(w_eco153, a[1], !b[2], a[5], b[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_154(w_eco154, a[7], b[4], !a[4], b[6], a[6], !a[0]);
	and _ECO_155(w_eco155, a[1], !b[2], a[5], !b[7], a[7], !b[4], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_156(w_eco156, a[1], !b[7], a[7], !a[6], a[0], !b[0]);
	and _ECO_157(w_eco157, a[2], a[1], !b[2], a[5], !b[7], a[7], !b[4], !a[4], b[6], a[6], b[1], a[0]);
	and _ECO_158(w_eco158, a[1], a[7], !a[4], b[6], a[6], !b[0]);
	and _ECO_159(w_eco159, a[1], !b[2], a[5], !a[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_160(w_eco160, a[1], !b[2], a[5], !a[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_161(w_eco161, a[1], !b[2], b[5], b[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_162(w_eco162, a[1], !b[2], b[5], b[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_163(w_eco163, a[2], !b[2], b[5], !a[5], !a[7], a[4], !a[0], b[0]);
	and _ECO_164(w_eco164, a[2], !b[2], b[5], !a[5], !a[7], !b[4], !a[0], b[0]);
	and _ECO_165(w_eco165, a[2], !b[2], b[5], !a[5], a[4], !a[6], !a[0], b[0]);
	and _ECO_166(w_eco166, a[2], !b[2], b[5], !a[5], !b[4], !a[6], !a[0], b[0]);
	and _ECO_167(w_eco167, b[5], !a[5], a[7], b[6], a[6], !b[1], a[0]);
	and _ECO_168(w_eco168, a[1], a[7], b[4], b[6], a[6], !b[0]);
	and _ECO_169(w_eco169, a[2], a[1], !b[2], a[5], !b[7], a[7], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_170(w_eco170, a[1], !b[2], a[5], !b[7], a[7], !b[6], a[6], b[1], b[0]);
	and _ECO_171(w_eco171, a[1], !b[5], a[7], b[4], !a[6], !b[0]);
	and _ECO_172(w_eco172, a[1], !b[5], a[7], !a[4], !a[6], !b[0]);
	and _ECO_173(w_eco173, a[2], a[1], !b[2], !b[5], !b[7], a[7], !b[4], a[6], b[1], a[0], b[0]);
	and _ECO_174(w_eco174, !b[5], a[5], !a[7], !b[6], !a[0]);
	and _ECO_175(w_eco175, !b[5], a[5], !a[7], b[4], !a[4], !b[0]);
	and _ECO_176(w_eco176, a[2], a[1], !b[2], !b[5], !b[7], a[7], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_177(w_eco177, a[2], !a[1], !b[2], a[5], b[7], a[4], a[6], b[1]);
	and _ECO_178(w_eco178, a[2], !a[1], !b[2], a[5], b[7], !b[4], a[6], b[1]);
	and _ECO_179(w_eco179, a[2], !a[1], !b[2], a[5], !a[7], a[4], a[6], b[1]);
	and _ECO_180(w_eco180, a[2], !a[1], !b[2], a[5], !a[7], !b[4], a[6], b[1]);
	and _ECO_181(w_eco181, a[2], !a[1], !b[2], b[5], !a[5], !b[1], a[0]);
	and _ECO_182(w_eco182, !a[1], !b[5], !b[7], b[4], !a[4], b[6]);
	and _ECO_183(w_eco183, !a[2], a[1], a[5], b[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_184(w_eco184, !a[2], a[1], a[5], b[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_185(w_eco185, !a[2], b[2], b[4], !a[4], !b[1], a[0]);
	and _ECO_186(w_eco186, !a[2], a[1], b[2], b[4], !a[4], a[0], !b[0]);
	and _ECO_187(w_eco187, !a[2], a[1], a[5], !a[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_188(w_eco188, !a[2], a[1], a[5], !a[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_189(w_eco189, !a[2], a[1], b[5], b[7], a[4], !b[6], !b[1], b[0]);
	and _ECO_190(w_eco190, !a[2], a[1], b[5], b[7], !b[4], !b[6], !b[1], b[0]);
	and _ECO_191(w_eco191, !a[2], b[2], !a[3], !b[1], a[0], b[3]);
	and _ECO_192(w_eco192, a[1], !a[3], !b[6], !a[0], b[3]);
	and _ECO_193(w_eco193, !a[2], a[1], b[2], !a[3], a[0], b[3], !b[0]);
	and _ECO_194(w_eco194, a[1], !b[5], !a[5], b[7], !a[7], !b[4], b[1], a[0], !b[3], b[0]);
	and _ECO_195(w_eco195, !a[1], b[2], a[7], !a[4], b[6], a[6], b[1]);
	and _ECO_196(w_eco196, !a[2], b[5], !a[5], !a[7], a[3], a[4], !b[1], !b[3], b[0]);
	and _ECO_197(w_eco197, !a[2], b[5], !a[5], !a[7], a[3], !b[4], !b[1], !b[3], b[0]);
	and _ECO_198(w_eco198, !a[1], b[2], !b[5], a[7], b[4], b[6], b[1]);
	and _ECO_199(w_eco199, !a[1], !b[2], a[5], !a[7], a[3], a[4], a[6], !b[3]);
	and _ECO_200(w_eco200, !a[1], !b[2], a[5], !a[7], a[3], !b[4], a[6], !b[3]);
	and _ECO_201(w_eco201, !a[2], !a[1], a[7], b[4], b[6], a[6], b[3]);
	and _ECO_202(w_eco202, !a[2], !a[1], a[7], !a[4], b[6], a[6], b[3]);
	and _ECO_203(w_eco203, !a[1], !b[2], b[5], !a[5], a[3], a[4], !a[6], !b[3]);
	and _ECO_204(w_eco204, !a[1], !b[2], b[5], !a[5], a[3], !b[4], !a[6], !b[3]);
	and _ECO_205(w_eco205, !a[2], !a[1], !b[5], a[7], b[4], b[6], b[3]);
	and _ECO_206(w_eco206, !a[2], !a[1], !b[5], a[7], !a[4], b[6], b[3]);
	and _ECO_207(w_eco207, !a[2], !a[1], !b[5], !b[7], b[4], b[6], b[3]);
	and _ECO_208(w_eco208, !a[2], !a[1], !b[5], !b[7], !a[4], b[6], b[3]);
	and _ECO_209(w_eco209, a[1], b[2], b[5], b[7], a[3], b[4], a[4], !b[6], b[1], a[0], b[0]);
	and _ECO_210(w_eco210, b[4], !a[4], !a[6], !b[1], a[0]);
	and _ECO_211(w_eco211, a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !b[6], b[1], a[0], b[0]);
	and _ECO_212(w_eco212, a[2], a[1], b[5], a[5], b[7], !a[7], b[4], !a[4], a[6], b[1], a[0], b[0]);
	and _ECO_213(w_eco213, a[1], b[4], !a[4], !a[6], a[0], !b[0]);
	and _ECO_214(w_eco214, a[2], a[1], a[5], !b[7], a[7], !b[6], a[6], b[1], b[0]);
	and _ECO_215(w_eco215, !b[7], !a[7], b[6], a[6], !a[0]);
	and _ECO_216(w_eco216, a[1], b[2], b[5], !a[7], a[3], b[4], a[4], !b[6], b[1], a[0], b[0]);
	and _ECO_217(w_eco217, a[5], !a[7], !b[4], a[4], !b[6], !b[0]);
	and _ECO_218(w_eco218, a[1], b[2], b[5], !a[7], a[3], !b[4], !a[4], !b[6], b[1], a[0], b[0]);
	and _ECO_219(w_eco219, !b[7], !a[7], b[6], a[6], !b[0]);
	and _ECO_220(w_eco220, a[1], b[5], a[5], !a[7], a[3], !b[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_221(w_eco221, b[5], !a[5], !a[3], !b[1], a[0], b[3]);
	and _ECO_222(w_eco222, a[5], b[7], !b[4], a[4], a[6], !b[0]);
	and _ECO_223(w_eco223, a[1], a[5], b[7], a[3], !b[4], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_224(w_eco224, a[2], b[2], !b[5], a[5], b[4], !a[6], !b[1], a[0]);
	and _ECO_225(w_eco225, !a[3], !a[6], !b[1], a[0], b[3]);
	and _ECO_226(w_eco226, b[4], !a[4], !b[6], !b[1], !a[0]);
	and _ECO_227(w_eco227, !a[3], !b[6], !b[1], !a[0], b[3]);
	and _ECO_228(w_eco228, a[2], b[2], !b[5], a[5], !a[4], !a[6], !b[1], !b[3]);
	and _ECO_229(w_eco229, b[7], a[7], b[6], a[6], !a[0]);
	and _ECO_230(w_eco230, b[7], a[7], !b[4], a[4], !b[6], !a[6], !a[0]);
	and _ECO_231(w_eco231, a[2], a[1], !b[5], !a[5], b[7], !a[7], a[6], b[1], a[0], b[0]);
	and _ECO_232(w_eco232, a[1], !a[3], !a[6], a[0], b[3], !b[0]);
	and _ECO_233(w_eco233, a[2], a[1], !b[5], !b[7], a[7], !b[6], a[6], b[1], b[0]);
	and _ECO_234(w_eco234, !b[5], !b[7], !a[7], !b[6], !a[6], !a[0]);
	and _ECO_235(w_eco235, a[2], !b[2], a[5], b[7], a[4], !b[6], !a[0], b[0]);
	and _ECO_236(w_eco236, a[2], !b[2], a[5], b[7], !b[4], !b[6], !a[0], b[0]);
	and _ECO_237(w_eco237, a[1], !b[2], a[5], !a[7], a[4], a[6], !b[1], b[0]);
	and _ECO_238(w_eco238, a[1], !b[2], a[5], !a[7], !b[4], a[6], !b[1], b[0]);
	and _ECO_239(w_eco239, a[2], !b[2], a[5], !a[7], a[4], !b[6], !a[0], b[0]);
	and _ECO_240(w_eco240, a[2], !b[2], a[5], !a[7], !b[4], !b[6], !a[0], b[0]);
	and _ECO_241(w_eco241, !b[5], a[5], !a[7], a[6], !a[0]);
	and _ECO_242(w_eco242, a[2], a[1], !b[2], !b[5], a[5], !a[7], a[3], b[4], a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_243(w_eco243, a[1], !b[5], a[5], b[4], !a[6], !b[0]);
	and _ECO_244(w_eco244, !b[5], a[5], !a[7], a[6], !b[0]);
	and _ECO_245(w_eco245, a[2], a[1], !b[2], !b[5], a[5], !a[7], a[3], !b[4], !a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_246(w_eco246, a[1], !b[5], a[5], !a[4], !a[6], !b[0]);
	and _ECO_247(w_eco247, a[2], a[1], !b[2], !b[5], !b[7], !a[7], a[3], b[4], a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_248(w_eco248, a[1], !b[5], !b[7], b[4], !a[6], !b[0]);
	and _ECO_249(w_eco249, a[2], a[1], !b[5], !a[5], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_250(w_eco250, b[2], !b[5], !b[7], !a[7], !a[4], !a[6], !b[0]);
	and _ECO_251(w_eco251, a[2], a[1], !b[2], !b[5], !b[7], !a[7], a[3], !b[4], !a[4], b[6], !a[6], b[1], a[0]);
	and _ECO_252(w_eco252, a[1], !b[5], !b[7], !a[4], !a[6], !b[0]);
	and _ECO_253(w_eco253, !a[1], b[7], a[7], !b[4], a[4], !b[6], !a[6]);
	and _ECO_254(w_eco254, a[2], !a[1], !b[2], a[5], !a[7], a[4], a[6], !b[3]);
	and _ECO_255(w_eco255, a[2], !a[1], !b[2], a[5], !a[7], !b[4], a[6], !b[3]);
	and _ECO_256(w_eco256, !a[1], a[7], b[4], !a[4], b[6], a[6]);
	and _ECO_257(w_eco257, a[2], !a[1], !b[2], b[5], !a[5], a[4], !a[6], a[0]);
	and _ECO_258(w_eco258, a[2], !a[1], !b[2], b[5], !a[5], !b[4], !a[6], a[0]);
	and _ECO_259(w_eco259, !a[2], a[1], a[5], !a[7], a[4], a[6], !b[1], b[0]);
	and _ECO_260(w_eco260, !a[2], a[1], a[5], !a[7], !b[4], a[6], !b[1], b[0]);
	and _ECO_261(w_eco261, a[1], b[2], b[5], b[7], !a[7], b[4], a[4], b[1], a[0], !b[3], b[0]);
	and _ECO_262(w_eco262, a[1], b[2], b[5], b[7], !a[7], !b[4], !a[4], b[1], a[0], !b[3], b[0]);
	and _ECO_263(w_eco263, b[2], a[7], !a[4], b[6], a[6], b[1], !a[0]);
	and _ECO_264(w_eco264, !a[2], a[1], b[5], !a[5], a[4], !a[6], !b[1], b[0]);
	and _ECO_265(w_eco265, !a[2], a[1], b[5], !a[5], !b[4], !a[6], !b[1], b[0]);
	and _ECO_266(w_eco266, a[1], !b[5], !a[5], b[7], !a[7], a[4], b[1], a[0], !b[3], b[0]);
	and _ECO_267(w_eco267, a[1], !b[2], b[5], a[5], b[7], !a[7], b[4], !a[4], a[6], b[1], a[0], b[0]);
	and _ECO_268(w_eco268, !a[2], a[1], !b[2], b[5], a[5], b[7], !a[7], !a[3], b[4], a[6], b[1], a[0], b[0]);
	and _ECO_269(w_eco269, !a[2], a[1], !b[2], b[5], a[5], b[7], !a[7], !a[3], !a[4], a[6], b[1], a[0], b[0]);
	and _ECO_270(w_eco270, !a[2], a[1], !a[5], b[7], !a[7], a[3], b[4], a[4], b[1], a[0], b[3], b[0]);
	and _ECO_271(w_eco271, !b[2], b[5], !a[5], !a[7], a[3], a[4], !a[0], !b[3], b[0]);
	and _ECO_272(w_eco272, !a[2], a[1], !a[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], a[0], b[3], b[0]);
	and _ECO_273(w_eco273, !b[2], b[5], !a[5], !a[7], a[3], !b[4], !a[0], !b[3], b[0]);
	and _ECO_274(w_eco274, !a[2], !b[5], a[7], !a[3], b[4], b[6], b[1], !a[0]);
	and _ECO_275(w_eco275, !a[2], !b[5], a[7], !a[3], !a[4], b[6], b[1], !a[0]);
	and _ECO_276(w_eco276, a[1], !b[2], !b[5], !a[5], b[7], !a[7], a[6], b[1], a[0], b[0]);
	and _ECO_277(w_eco277, a[1], !b[2], !b[5], !b[7], a[7], !b[4], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_278(w_eco278, a[1], !b[2], !b[5], !b[7], a[7], !b[6], a[6], b[1], b[0]);
	and _ECO_279(w_eco279, !a[2], a[5], b[7], a[3], a[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_280(w_eco280, !a[2], a[5], b[7], a[3], !b[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_281(w_eco281, !a[2], a[5], !a[7], a[3], a[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_282(w_eco282, !a[2], a[5], !a[7], a[3], !b[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_283(w_eco283, !a[2], b[5], b[7], a[3], a[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_284(w_eco284, !a[2], b[5], b[7], a[3], !b[4], !b[6], !b[1], !b[3], b[0]);
	and _ECO_285(w_eco285, !a[1], !b[2], b[5], !a[5], a[3], a[4], !b[6], !b[3]);
	and _ECO_286(w_eco286, !a[1], !b[2], b[5], !a[5], a[3], !b[4], !b[6], !b[3]);
	and _ECO_287(w_eco287, a[1], b[5], a[5], b[7], a[3], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_288(w_eco288, a[2], a[1], b[5], a[5], b[4], !a[4], !b[6], a[6], b[1], b[0]);
	and _ECO_289(w_eco289, a[1], b[5], a[5], b[7], a[3], !b[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_290(w_eco290, a[2], a[1], b[2], b[5], a[5], b[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_291(w_eco291, a[2], a[1], b[2], b[5], a[5], !a[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_292(w_eco292, a[1], a[5], !a[7], !a[3], a[4], a[6], !b[1], b[3], b[0]);
	and _ECO_293(w_eco293, a[1], a[5], !a[7], !a[3], !b[4], a[6], !b[1], b[3], b[0]);
	and _ECO_294(w_eco294, a[2], a[1], a[5], !b[7], a[7], !b[4], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_295(w_eco295, a[2], b[2], a[7], b[4], b[6], a[6], !b[1], !b[3]);
	and _ECO_296(w_eco296, a[2], b[2], a[7], !a[4], b[6], a[6], !b[1], !b[3]);
	and _ECO_297(w_eco297, a[1], b[5], a[5], !a[7], a[3], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_298(w_eco298, a[1], b[2], b[5], !a[7], b[4], a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_299(w_eco299, a[1], b[2], b[5], !a[7], !b[4], !a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_300(w_eco300, a[1], b[2], b[5], b[7], a[3], b[4], a[4], !a[6], b[1], a[0], b[0]);
	and _ECO_301(w_eco301, a[1], b[2], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], a[0], b[0]);
	and _ECO_302(w_eco302, a[2], b[2], !b[5], a[5], b[4], !b[1], !a[0], !b[3]);
	and _ECO_303(w_eco303, a[1], a[5], b[7], !b[4], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_304(w_eco304, a[1], a[5], !a[7], a[3], !b[4], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_305(w_eco305, !b[5], b[7], a[7], !b[6], !a[6], !a[0]);
	and _ECO_306(w_eco306, a[1], !b[2], !b[5], !a[5], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_307(w_eco307, b[7], a[7], b[6], a[6], !b[0]);
	and _ECO_308(w_eco308, a[1], !b[5], b[7], a[3], !b[4], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_309(w_eco309, b[7], a[7], !b[4], a[4], !b[6], !a[6], !b[0]);
	and _ECO_310(w_eco310, a[1], !b[5], !a[5], b[7], a[3], !b[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_311(w_eco311, a[2], b[2], !b[5], a[7], b[4], !a[6], !b[1], !b[3]);
	and _ECO_312(w_eco312, a[2], b[2], !b[5], a[7], !a[4], !a[6], !b[1], !b[3]);
	and _ECO_313(w_eco313, a[2], a[1], !b[5], !b[7], a[7], !b[4], a[4], a[6], b[1], a[0], b[0]);
	and _ECO_314(w_eco314, a[1], !b[5], !a[7], a[3], !b[4], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_315(w_eco315, !b[7], !a[7], !b[4], a[4], !b[6], !a[6], !b[0]);
	and _ECO_316(w_eco316, a[1], !b[5], !a[5], !a[7], a[3], !b[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_317(w_eco317, a[2], b[2], !b[5], !b[7], b[4], !a[6], !b[1], !b[3]);
	and _ECO_318(w_eco318, a[2], b[2], !b[5], !b[7], !a[4], !a[6], !b[1], !b[3]);
	and _ECO_319(w_eco319, a[2], !b[2], a[5], !a[7], a[4], a[6], !a[0], b[0]);
	and _ECO_320(w_eco320, a[2], !b[2], a[5], !a[7], !b[4], a[6], !a[0], b[0]);
	and _ECO_321(w_eco321, a[1], b[5], a[5], b[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_322(w_eco322, a[1], b[5], a[5], b[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_323(w_eco323, a[1], b[5], a[5], !a[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_324(w_eco324, a[1], !b[2], b[5], !a[5], !b[1], a[0], b[0]);
	and _ECO_325(w_eco325, a[2], !b[2], b[5], b[7], a[4], a[6], !a[0], b[0]);
	and _ECO_326(w_eco326, a[2], !b[2], b[5], b[7], !b[4], a[6], !a[0], b[0]);
	and _ECO_327(w_eco327, a[1], b[5], !a[5], !a[3], a[0], b[3], !b[0]);
	and _ECO_328(w_eco328, !a[2], a[1], !a[5], b[7], !a[7], !a[3], b[4], a[4], b[1], a[0], !b[3], b[0]);
	and _ECO_329(w_eco329, !a[2], a[1], !a[5], b[7], !a[7], !a[3], !b[4], !a[4], b[1], a[0], !b[3], b[0]);
	and _ECO_330(w_eco330, a[1], b[2], b[5], b[7], b[4], a[4], !b[6], b[1], a[0], !b[3], b[0]);
	and _ECO_331(w_eco331, a[1], b[2], b[5], b[7], !b[4], !a[4], !b[6], b[1], a[0], !b[3], b[0]);
	and _ECO_332(w_eco332, a[1], b[5], !a[5], !a[7], !a[3], a[4], !b[1], b[3], b[0]);
	and _ECO_333(w_eco333, a[1], b[5], !a[5], !a[7], !a[3], !b[4], !b[1], b[3], b[0]);
	and _ECO_334(w_eco334, a[2], a[1], !b[2], a[5], b[7], a[3], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_335(w_eco335, !b[5], a[5], b[7], a[6], !b[0]);
	and _ECO_336(w_eco336, a[2], a[1], !b[2], a[5], b[7], a[3], !b[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_337(w_eco337, a[2], a[1], !b[2], a[5], b[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_338(w_eco338, a[2], a[1], !b[2], a[5], b[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_339(w_eco339, a[2], a[1], !b[2], a[5], !a[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_340(w_eco340, a[2], a[1], !b[2], !b[5], b[7], a[3], a[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_341(w_eco341, a[2], a[1], !b[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], b[1], a[0], b[0]);
	and _ECO_342(w_eco342, a[2], a[1], !b[2], !b[5], b[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_343(w_eco343, a[2], a[1], !b[2], !b[5], !a[7], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_344(w_eco344, a[2], !a[1], !b[2], a[5], b[7], a[4], a[6], !b[3]);
	and _ECO_345(w_eco345, a[2], !a[1], !b[2], a[5], b[7], !b[4], a[6], !b[3]);
	and _ECO_346(w_eco346, a[2], !b[2], a[5], !a[7], a[4], a[6], !b[1], b[0]);
	and _ECO_347(w_eco347, a[2], !b[2], a[5], !a[7], !b[4], a[6], !b[1], b[0]);
	and _ECO_348(w_eco348, a[7], !a[3], b[4], b[6], a[6], !b[1], b[3], !b[0]);
	and _ECO_349(w_eco349, a[7], !a[3], !a[4], b[6], a[6], !b[1], b[3], !b[0]);
	and _ECO_350(w_eco350, !b[5], a[5], !a[3], b[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_351(w_eco351, !b[5], a[5], !a[3], !a[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_352(w_eco352, a[2], !a[1], !b[2], b[5], !a[5], a[4], !a[6], b[1]);
	and _ECO_353(w_eco353, a[2], !a[1], !b[2], b[5], !a[5], !b[4], !a[6], b[1]);
	and _ECO_354(w_eco354, a[2], !a[1], !b[2], b[5], !a[5], !a[7], a[4], !b[3]);
	and _ECO_355(w_eco355, a[2], !a[1], !b[2], b[5], !a[5], !a[7], !b[4], !b[3]);
	and _ECO_356(w_eco356, !b[5], !b[7], !a[3], b[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_357(w_eco357, !b[5], !b[7], !a[3], !a[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_358(w_eco358, a[1], !b[5], !a[5], b[7], a[3], a[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_359(w_eco359, a[1], !b[5], !a[5], !a[7], a[3], a[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_360(w_eco360, !a[2], a[1], b[5], b[7], a[3], b[4], a[4], !b[6], a[0], b[3], b[0]);
	and _ECO_361(w_eco361, !b[2], a[5], b[7], a[3], a[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_362(w_eco362, a[1], !b[2], b[5], a[5], b[4], !a[4], !b[6], a[6], b[1], b[0]);
	and _ECO_363(w_eco363, !a[2], a[1], b[5], b[7], a[3], !b[4], !a[4], !b[6], a[0], b[3], b[0]);
	and _ECO_364(w_eco364, !b[2], a[5], b[7], a[3], !b[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_365(w_eco365, !a[2], a[1], !b[2], b[5], a[5], !a[3], b[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_366(w_eco366, !a[2], a[1], !b[2], b[5], a[5], !a[3], !a[4], !b[6], a[6], b[1], a[0], b[0]);
	and _ECO_367(w_eco367, !a[2], a[7], !a[3], b[4], b[6], a[6], b[1], !a[0]);
	and _ECO_368(w_eco368, !a[2], a[7], !a[3], !a[4], b[6], a[6], b[1], !a[0]);
	and _ECO_369(w_eco369, !a[2], a[1], b[5], !a[7], a[3], b[4], a[4], !b[6], a[0], b[3], b[0]);
	and _ECO_370(w_eco370, !b[2], a[5], !a[7], a[3], a[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_371(w_eco371, !a[2], a[1], b[5], !a[7], a[3], !b[4], !a[4], !b[6], a[0], b[3], b[0]);
	and _ECO_372(w_eco372, !b[2], a[5], !a[7], a[3], !b[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_373(w_eco373, !a[2], a[1], b[5], !a[7], !a[3], b[4], a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_374(w_eco374, !b[2], b[5], b[7], a[3], a[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_375(w_eco375, !b[2], b[5], b[7], a[3], !b[4], !b[6], !a[0], !b[3], b[0]);
	and _ECO_376(w_eco376, !a[2], a[1], b[5], b[7], !a[3], b[4], a[4], !b[6], a[0], !b[3], b[0]);
	and _ECO_377(w_eco377, !a[2], a[1], b[5], b[7], !a[3], !b[4], !a[4], !b[6], a[0], !b[3], b[0]);
	and _ECO_378(w_eco378, !a[2], a[1], b[5], !a[7], !a[3], !b[4], !a[4], !b[6], a[0], !b[3], b[0]);
	and _ECO_379(w_eco379, !a[2], !b[5], a[5], !a[3], b[4], b[6], b[1], !a[0]);
	and _ECO_380(w_eco380, !a[2], !b[5], a[5], !a[3], !a[4], b[6], b[1], !a[0]);
	and _ECO_381(w_eco381, a[1], !b[2], a[5], b[7], a[3], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_382(w_eco382, !a[2], !b[5], a[5], b[4], b[6], b[1], !a[0], b[3]);
	and _ECO_383(w_eco383, a[1], !b[2], a[5], b[7], a[3], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_384(w_eco384, !a[2], !b[5], a[5], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_385(w_eco385, !a[2], !b[5], !b[7], !a[3], b[4], b[6], b[1], !a[0]);
	and _ECO_386(w_eco386, !a[2], !b[5], !b[7], !a[3], !a[4], b[6], b[1], !a[0]);
	and _ECO_387(w_eco387, !a[2], a[5], !a[7], a[3], a[4], a[6], !b[1], !b[3], b[0]);
	and _ECO_388(w_eco388, !a[2], a[5], !a[7], a[3], !b[4], a[6], !b[1], !b[3], b[0]);
	and _ECO_389(w_eco389, !a[1], b[2], a[7], b[4], b[6], a[6], a[0]);
	and _ECO_390(w_eco390, !a[2], b[5], !a[5], a[3], a[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_391(w_eco391, !a[2], b[5], !a[5], a[3], !b[4], !a[6], !b[1], !b[3], b[0]);
	and _ECO_392(w_eco392, b[2], a[7], b[4], b[6], a[6], !b[0]);
	and _ECO_393(w_eco393, b[2], a[7], !a[4], b[6], a[6], !b[0]);
	and _ECO_394(w_eco394, !a[1], b[2], !b[5], a[7], !a[4], b[6], b[1]);
	and _ECO_395(w_eco395, b[2], !b[5], a[7], b[4], !a[6], !b[1], !b[0]);
	and _ECO_396(w_eco396, b[2], !b[5], a[7], !a[4], !a[6], !b[1], !b[0]);
	and _ECO_397(w_eco397, !a[1], b[2], !b[5], a[5], b[4], b[6], b[1]);
	and _ECO_398(w_eco398, !a[1], b[2], !b[5], a[5], !a[4], b[6], b[1]);
	and _ECO_399(w_eco399, !a[1], b[2], !b[5], !b[7], b[4], b[6], b[1]);
	and _ECO_400(w_eco400, b[2], !b[5], !b[7], b[4], !a[6], !b[1], !b[0]);
	and _ECO_401(w_eco401, a[1], a[5], b[7], !a[3], a[4], !b[1], a[0], b[3], b[0]);
	and _ECO_402(w_eco402, a[1], a[5], b[7], !a[3], !b[4], !b[1], a[0], b[3], b[0]);
	and _ECO_403(w_eco403, a[2], a[1], b[2], b[5], a[5], b[7], !a[7], b[4], a[6], b[1], a[0], b[0]);
	and _ECO_404(w_eco404, a[2], a[1], b[2], b[5], a[5], b[7], !a[7], !a[4], a[6], b[1], a[0], b[0]);
	and _ECO_405(w_eco405, a[1], b[2], b[5], b[7], b[4], a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_406(w_eco406, a[1], b[5], !a[5], !a[3], a[4], !a[6], !b[1], b[3], b[0]);
	and _ECO_407(w_eco407, a[1], b[2], b[5], b[7], !b[4], !a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_408(w_eco408, a[1], b[5], !a[5], !a[3], !b[4], !a[6], !b[1], b[3], b[0]);
	and _ECO_409(w_eco409, a[1], b[2], b[5], !a[7], a[3], b[4], a[4], !a[6], b[1], a[0], b[0]);
	and _ECO_410(w_eco410, a[1], b[2], b[5], !a[7], a[3], !b[4], !a[4], !a[6], b[1], a[0], b[0]);
	and _ECO_411(w_eco411, a[1], b[2], b[5], !a[7], b[4], a[4], !b[6], b[1], a[0], !b[3], b[0]);
	and _ECO_412(w_eco412, a[1], b[2], !a[5], !a[7], !b[4], !a[4], !b[6], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_413(w_eco413, a[1], a[5], !a[7], !b[4], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_414(w_eco414, a[1], !b[5], b[7], !b[4], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_415(w_eco415, a[1], !b[5], !a[5], b[7], !b[4], !b[6], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_416(w_eco416, a[1], !b[5], !a[7], !b[4], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_417(w_eco417, a[1], !b[5], !a[5], !a[7], a[4], !b[6], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_418(w_eco418, a[1], b[5], a[5], !a[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_419(w_eco419, a[2], a[1], !b[2], a[5], !a[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_420(w_eco420, a[2], a[1], !b[2], !b[5], b[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_421(w_eco421, a[2], a[1], !b[2], !b[5], !a[7], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_422(w_eco422, a[2], !b[2], a[5], b[7], a[4], a[6], !b[1], b[0]);
	and _ECO_423(w_eco423, a[2], !b[2], a[5], b[7], !b[4], a[6], !b[1], b[0]);
	and _ECO_424(w_eco424, a[2], !a[1], !b[2], b[5], !a[5], a[4], !a[6], !b[3]);
	and _ECO_425(w_eco425, a[2], !a[1], !b[2], b[5], !a[5], !b[4], !a[6], !b[3]);
	and _ECO_426(w_eco426, a[2], !a[1], !b[2], b[5], !a[5], a[3], a[4], !a[6]);
	and _ECO_427(w_eco427, a[2], !a[1], !b[2], b[5], !a[5], a[3], !b[4], !a[6]);
	and _ECO_428(w_eco428, !b[5], a[7], !a[3], b[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_429(w_eco429, !b[5], a[7], !a[3], !a[4], !b[1], !a[0], b[3], !b[0]);
	and _ECO_430(w_eco430, a[1], !b[5], !a[5], b[7], a[4], !b[6], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_431(w_eco431, !a[2], a[1], b[5], b[7], !a[7], a[3], b[4], a[4], b[1], a[0], b[3], b[0]);
	and _ECO_432(w_eco432, !b[2], a[5], !a[7], a[3], a[4], a[6], !a[0], !b[3], b[0]);
	and _ECO_433(w_eco433, !a[2], a[1], b[5], b[7], !a[7], a[3], !b[4], !a[4], b[1], a[0], b[3], b[0]);
	and _ECO_434(w_eco434, !b[2], a[5], !a[7], a[3], !b[4], a[6], !a[0], !b[3], b[0]);
	and _ECO_435(w_eco435, a[1], !b[2], a[5], !b[7], a[7], a[3], a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_436(w_eco436, !a[2], a[7], b[4], b[6], a[6], b[1], !a[0], b[3]);
	and _ECO_437(w_eco437, a[1], !b[2], a[5], !b[7], a[7], a[3], !b[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_438(w_eco438, !a[2], a[7], !a[4], b[6], a[6], b[1], !a[0], b[3]);
	and _ECO_439(w_eco439, !a[2], a[1], b[5], b[7], a[3], b[4], a[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_440(w_eco440, !b[2], b[5], !a[5], a[3], a[4], !a[6], !a[0], !b[3], b[0]);
	and _ECO_441(w_eco441, !a[2], a[1], b[5], b[7], a[3], !b[4], !a[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_442(w_eco442, !b[2], b[5], !a[5], a[3], !b[4], !a[6], !a[0], !b[3], b[0]);
	and _ECO_443(w_eco443, !a[2], a[1], b[5], b[7], !a[3], b[4], a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_444(w_eco444, !a[2], a[1], b[5], b[7], !a[3], !b[4], !a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_445(w_eco445, !a[2], a[1], b[5], !a[7], a[3], b[4], a[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_446(w_eco446, !a[2], a[1], b[5], !a[7], a[3], !b[4], !a[4], !a[6], b[1], a[0], b[3], b[0]);
	and _ECO_447(w_eco447, !a[2], a[1], !a[5], !a[7], !a[3], b[4], a[4], !b[6], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_448(w_eco448, !a[2], a[1], b[5], !a[7], !a[3], !b[4], !a[4], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_449(w_eco449, a[1], !b[2], a[5], !a[7], a[3], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_450(w_eco450, a[1], !b[2], a[5], !a[7], a[3], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_451(w_eco451, a[1], !b[2], !b[5], b[7], a[3], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_452(w_eco452, !a[2], !b[5], a[7], b[4], b[6], b[1], !a[0], b[3]);
	and _ECO_453(w_eco453, a[1], !b[2], !b[5], b[7], a[3], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_454(w_eco454, !a[2], !b[5], a[7], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_455(w_eco455, a[1], !b[2], !b[5], !b[7], a[7], a[3], a[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_456(w_eco456, a[1], !b[2], !b[5], !b[7], a[7], a[3], !b[4], a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_457(w_eco457, a[1], !b[2], !b[5], !a[7], a[3], a[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_458(w_eco458, !a[2], !b[5], !b[7], b[4], b[6], b[1], !a[0], b[3]);
	and _ECO_459(w_eco459, a[1], !b[2], !b[5], !a[7], a[3], !b[4], b[6], !a[6], b[1], a[0], !b[3], b[0]);
	and _ECO_460(w_eco460, !a[2], !b[5], !b[7], !a[4], b[6], b[1], !a[0], b[3]);
	and _ECO_461(w_eco461, !a[1], b[2], !b[5], !b[7], !a[4], b[6], b[1]);
	or _ECO_462(w_eco462, w_eco0, w_eco1, w_eco2, w_eco3, w_eco4, w_eco5, w_eco6, w_eco7, w_eco8, w_eco9, w_eco10, w_eco11, w_eco12, w_eco13, w_eco14, w_eco15, w_eco16, w_eco17, w_eco18, w_eco19, w_eco20, w_eco21, w_eco22, w_eco23, w_eco24, w_eco25, w_eco26, w_eco27, w_eco28, w_eco29, w_eco30, w_eco31, w_eco32, w_eco33, w_eco34, w_eco35, w_eco36, w_eco37, w_eco38, w_eco39, w_eco40, w_eco41, w_eco42, w_eco43, w_eco44, w_eco45, w_eco46, w_eco47, w_eco48, w_eco49, w_eco50, w_eco51, w_eco52, w_eco53, w_eco54, w_eco55, w_eco56, w_eco57, w_eco58, w_eco59, w_eco60, w_eco61, w_eco62, w_eco63, w_eco64, w_eco65, w_eco66, w_eco67, w_eco68, w_eco69, w_eco70, w_eco71, w_eco72, w_eco73, w_eco74, w_eco75, w_eco76, w_eco77, w_eco78, w_eco79, w_eco80, w_eco81, w_eco82, w_eco83, w_eco84, w_eco85, w_eco86, w_eco87, w_eco88, w_eco89, w_eco90, w_eco91, w_eco92, w_eco93, w_eco94, w_eco95, w_eco96, w_eco97, w_eco98, w_eco99, w_eco100, w_eco101, w_eco102, w_eco103, w_eco104, w_eco105, w_eco106, w_eco107, w_eco108, w_eco109, w_eco110, w_eco111, w_eco112, w_eco113, w_eco114, w_eco115, w_eco116, w_eco117, w_eco118, w_eco119, w_eco120, w_eco121, w_eco122, w_eco123, w_eco124, w_eco125, w_eco126, w_eco127, w_eco128, w_eco129, w_eco130, w_eco131, w_eco132, w_eco133, w_eco134, w_eco135, w_eco136, w_eco137, w_eco138, w_eco139, w_eco140, w_eco141, w_eco142, w_eco143, w_eco144, w_eco145, w_eco146, w_eco147, w_eco148, w_eco149, w_eco150, w_eco151, w_eco152, w_eco153, w_eco154, w_eco155, w_eco156, w_eco157, w_eco158, w_eco159, w_eco160, w_eco161, w_eco162, w_eco163, w_eco164, w_eco165, w_eco166, w_eco167, w_eco168, w_eco169, w_eco170, w_eco171, w_eco172, w_eco173, w_eco174, w_eco175, w_eco176, w_eco177, w_eco178, w_eco179, w_eco180, w_eco181, w_eco182, w_eco183, w_eco184, w_eco185, w_eco186, w_eco187, w_eco188, w_eco189, w_eco190, w_eco191, w_eco192, w_eco193, w_eco194, w_eco195, w_eco196, w_eco197, w_eco198, w_eco199, w_eco200, w_eco201, w_eco202, w_eco203, w_eco204, w_eco205, w_eco206, w_eco207, w_eco208, w_eco209, w_eco210, w_eco211, w_eco212, w_eco213, w_eco214, w_eco215, w_eco216, w_eco217, w_eco218, w_eco219, w_eco220, w_eco221, w_eco222, w_eco223, w_eco224, w_eco225, w_eco226, w_eco227, w_eco228, w_eco229, w_eco230, w_eco231, w_eco232, w_eco233, w_eco234, w_eco235, w_eco236, w_eco237, w_eco238, w_eco239, w_eco240, w_eco241, w_eco242, w_eco243, w_eco244, w_eco245, w_eco246, w_eco247, w_eco248, w_eco249, w_eco250, w_eco251, w_eco252, w_eco253, w_eco254, w_eco255, w_eco256, w_eco257, w_eco258, w_eco259, w_eco260, w_eco261, w_eco262, w_eco263, w_eco264, w_eco265, w_eco266, w_eco267, w_eco268, w_eco269, w_eco270, w_eco271, w_eco272, w_eco273, w_eco274, w_eco275, w_eco276, w_eco277, w_eco278, w_eco279, w_eco280, w_eco281, w_eco282, w_eco283, w_eco284, w_eco285, w_eco286, w_eco287, w_eco288, w_eco289, w_eco290, w_eco291, w_eco292, w_eco293, w_eco294, w_eco295, w_eco296, w_eco297, w_eco298, w_eco299, w_eco300, w_eco301, w_eco302, w_eco303, w_eco304, w_eco305, w_eco306, w_eco307, w_eco308, w_eco309, w_eco310, w_eco311, w_eco312, w_eco313, w_eco314, w_eco315, w_eco316, w_eco317, w_eco318, w_eco319, w_eco320, w_eco321, w_eco322, w_eco323, w_eco324, w_eco325, w_eco326, w_eco327, w_eco328, w_eco329, w_eco330, w_eco331, w_eco332, w_eco333, w_eco334, w_eco335, w_eco336, w_eco337, w_eco338, w_eco339, w_eco340, w_eco341, w_eco342, w_eco343, w_eco344, w_eco345, w_eco346, w_eco347, w_eco348, w_eco349, w_eco350, w_eco351, w_eco352, w_eco353, w_eco354, w_eco355, w_eco356, w_eco357, w_eco358, w_eco359, w_eco360, w_eco361, w_eco362, w_eco363, w_eco364, w_eco365, w_eco366, w_eco367, w_eco368, w_eco369, w_eco370, w_eco371, w_eco372, w_eco373, w_eco374, w_eco375, w_eco376, w_eco377, w_eco378, w_eco379, w_eco380, w_eco381, w_eco382, w_eco383, w_eco384, w_eco385, w_eco386, w_eco387, w_eco388, w_eco389, w_eco390, w_eco391, w_eco392, w_eco393, w_eco394, w_eco395, w_eco396, w_eco397, w_eco398, w_eco399, w_eco400, w_eco401, w_eco402, w_eco403, w_eco404, w_eco405, w_eco406, w_eco407, w_eco408, w_eco409, w_eco410, w_eco411, w_eco412, w_eco413, w_eco414, w_eco415, w_eco416, w_eco417, w_eco418, w_eco419, w_eco420, w_eco421, w_eco422, w_eco423, w_eco424, w_eco425, w_eco426, w_eco427, w_eco428, w_eco429, w_eco430, w_eco431, w_eco432, w_eco433, w_eco434, w_eco435, w_eco436, w_eco437, w_eco438, w_eco439, w_eco440, w_eco441, w_eco442, w_eco443, w_eco444, w_eco445, w_eco446, w_eco447, w_eco448, w_eco449, w_eco450, w_eco451, w_eco452, w_eco453, w_eco454, w_eco455, w_eco456, w_eco457, w_eco458, w_eco459, w_eco460, w_eco461);
	xor _ECO_out0(a_gtet_b, sub_wire0, w_eco462);

endmodule